`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
bo49trehcslJg4im271Q32rlKfgWB3uwD/eNJhEuEToQZgacWRy2tbSPUU/O75ei
iNgfLX9Xv28pMqt4S7MJuJWBmGSmJiq8V6zd+RWJDGpmzq3C/uCz96ZJR2CvuMzz
8Zfw7KZ5csUXnr0u/BSxlozX23wgS42PkFWIvotXBV9Ve47pgGAsE2dgnk+ynj+U
jw220cdPSfxe9gBZk4RAue5SqqQtu5MHMvqdVBrVfuIy9ArUeA5tl7T3r1XIePNH
ykUi+3jTeglWhYLpXH2RCx4lxVsvThpKVwc+6+2f2c7Oc6ULpavnaXa1ZyU1VUtA
8nUMgpNsaNthmFAyEbC0e4Tey2u6zxbXVlylVmfMpk8DNrIDKLgT03n/qn4K8SuJ
q6PZkIG6f/9uL9GbQrrK0UJpugVOGWO3MH6GmQlo3rsbZEohahr8B9Lidq8nEwqp
mQ70g64i0wQFXcSDOCyhnvG183tlo6/IUR/3pOksIi4dV9AvwgTunUXLa7H7jLiQ
S/PSVr9qDSTlPCFR+LKIucksE/Oz0VdzluJDup4daJgtwn+QPUiT46+E8BRmww8J
ZJxrhQRMAe7I1YVPEiopUWc1je0aVTgowGHHSaX/po60BzZqbbQyS/YGm7RVzJ+e
EQvfoUh/JzQ9/RTcUxD3FyGuSamUfyglTkmFhScQxf7k94lE7h0UNWNBzLMgioBt
ySmokTZ1MY8KUNHMISdBELoQeKwAuhYUpWyNoQq3+TBWb3/7BJMxBr+pW47wi+3G
qoSfhPguB+quWlV1I9/ewQ/o1uvQ/uPTQoHO8iV6iB485imgil+XRLzJCfitF3rJ
XJ7xi2pfqv4Apm3bgKVutrnG66uodErFBa2zWWX3Gg6IzgYRfGAEVrNhiCDRcYLu
532vTfA4RTQJQ+5l6IOyB41Tk+udWqXOaVh52Gh3FX/A3zFAzkC8QkqZC1EICeTF
UIVx9/1d2MVBUJcWeHQ7QmYo5wGKGMUshDOzFZJpYfHhrfPGHHwf23jaVpIXd18J
j4jmkfjDc3h/9CRoonrhdeyUYi8F9Qy96mE+fL66fmPQMaBKYHajlVdPjsTTHWFA
P73s+kAqT/PoMDteME/dRpzDPW7PbBmztfrRbpQoaBXby5iWpgaiVcUF3c5sUzNY
5L1s8UAu5Thgt+1+cuzowPw66UFa+hZZfe0t0FvFapeIIaM3NL9KwP2QeAmVclHf
HfvaW77Om3NkIHAVBWLNHIscdzdMSeajXli6idu2tcTBzonPfrl5bjOMlu8f29S3
kOMlb0C2GfChy6F4g9PjcLI6fcTbPylCJuq2eOGEuujZI3lvlhJKjJ7UX0z1cGgh
W/467yPq/2ojo3Qey3QCBgrfBZOJIi3ewJHjiz+qYQVNO/DrryZBJ3dVeKpaQ3e+
CT2d+MPtM0mr4GVnAYAW6tT6+1rojRRsq8vwk7+NS6TK5pWyUrDhx404OBivjg9C
B7/FuMSmivmLgpuaXgb6+vMvm93HU/Th0MU06qp/Nw80j4riNR8oebqEAJ0BVnsR
qHlud8pUVsgEeQBdlXnunaDuDolsDGQybInY0vvdv1JMnPpT3JTAI6SZ5ViV3cpn
moizSLhrgqgd9oBZXRbYdPTxmNCwTnEhb09mNQxPq6cWMymJAllTV33/Jo7aek6i
lWI6yQCnTPhvIVGoVGDsp9RUFHs3qvnB1tHe+yWh/PtveWujM2Z0SVlX6NG7pGUc
826UUWdKbTlkPDL1+AbU4heO18tO5Yo4Ole79PbZL9o9N5GrpIYmMHW9wbB7pN6i
1hwZ8gNTttWPItTImNvv3Co7x6zH8++Zf3nnYeD8IBW73QDAEyWetuVAYu5/Toni
WHihVEUEQJNLB38DHzaxJndJPZnoPahqdF1Cq71Lyc9D+if+yW6RcBkhKoHGgPp3
nYS+fzMoCI7D1yATlQW2mnOK5PAXIuhfdV9XYfREfQlT7BuxXmM/oJxzlrhIiHdK
3eE5Q9GDZLif2jRrwCbJmg/YhgbWYjouoSM8T7p0u/NO9/6pe7+JnRPmjC3VaDuN
ERKm7JTwVhLjXGLjsp5lVNt8bDdjyHH9NG6O8obLw7jISpwke2XBVKYntDNcIFeL
DR7vAm1c+KLfc/+G/0zDQw7sHMCDzkVvIMvGOQnQd9Bx9AFO9/vvjnCAA04/6DxZ
JZV6xzzHkn7Tld1efYUeea27s/EppwuPnB5ZcA2tuslv70D//T5wmjjPrusXWjzb
etn9l1X8tmtXrj2qhhjyXU7Fux1if60NFCKgJZu2i8uG9AFIJCojJHtGEZKpaxCv
C9K3sZRJBUf9xJubf8GzpkyuTnMUnzUiYiMuFMDSe7O0uJc6UlwgmK1NbfXH6gHa
1O0EIYF+fauYzoqcAL3fsQGPnPRzNIEUroF2cthB21BwrYCz6klS54LDj2bSS17M
/cnnciXzGAgl32V1Q0Ps7khvUbXvG9V4JY+rqk7woZv6reaXEfdq2tJj2D7P2Ujs
4sjBBiAnAn26byKkvsxFm3dFAaSkCMdn0EeS3jtwqV8g3dlJZt9CeUnzKwvxLgAu
BP12qjQJoJR5OpNkwN7QbuP3m0532XTVtNE5lYe2sDJi1qdGWCaznonTtnG+6sOA
kQtCcDCZE1ivsEUgTm2TVI+TFN+D099eFGdyD3SW5crGZyUrM/6SA6y0zIdGz13A
FMZeH7586Zzpl1hqoF6y+sWOlOHRuGnkJv6iCZLkEd895OTCCzZ4/W1C+eMx6ITK
4ubo/ZrhjsVtajQfqxh39hKdia5K1lHIvZRMX52CgZYk7q9KR5WIcDD58f4kLpVx
oW/BqHTirzw6gVGRizUxRpgU9CdqUa8/+0G6NnJrjfR7oJeGrnspKJxVZVcpfBt4
NywGXeU1pNlR6/Q3l1QwDLMm7pk+bA3zumMPLDVnkhDNyk4GiUWZHf2ZF6lqxlde
CwFajwUzdozgIvkRiLKe9GvZsNa680WnsugKdhM0sfq7FaiRqXOxOOnrphtkEF8b
T7PkNzfAYEhv5k59TvU1DUJubcOV4MbpLDix+ltRFpvWiHy0BrxGMrJ+UZUwGhNl
kEOsMDB2OawUk0C4XCkwgLx744Jsx2H4kkr4kPUn7pY2R6OO82LJMNzEtmiHP85H
VTmfC2Qmh/giVyO50lFNYeSV4s9bQrSCPnshnxcWCOZiyx2W440N9td7AIVEUzu4
PhnnxEiRukObVgQ1QpCz9ddp7l88k1EpDpCoCsCi1qMynZ4yenl5QgpqMF/b13v9
gri5dTT2EBF2MhM/uq5IqY1qSz+sZHtX5Ax0HqlHSu3ihnCZRMOBOViachY7X86f
QFpg1XjrtdH2FWM5RgTBSJWUy4q0vUz3MVlyWhee9/wim+Aiz1jYJUc39DKQB3oe
mkQgNyqGIChskC/vDFpgj2jVFKZNOzOA1R7ZsFU322uBbYjy/fOi/j3D79AJFcBF
NLMzhK9OwZy88Hf1pDHY/BjLVHYWqPmGYdek91OMdUZtffsSmIFuofilt86K5N5x
cF5eUkmkOS69EXT5wqbp7lS4daq043HTg/KrINXw1LcHBJt4kwMCT0UrMZjxHHY6
zj+tVp4D0xZcIeycRCJeeSTbW0uPFpSapuNv5mRfNHJhLxWPvZyNyxmhGCfL9kwo
0OKQjlP4T3vv3QpFhgnKHhMvACIU9k9ima5qyonf0EMtTdmPyIieOaVSrJEu3MXv
BrGXnv0YyUxFqrfod4IsnU6lttXb/rNihUqLVJzy94tRjcCSgc1snhXacXp5mXlI
MxTFzEsltLUajC6vsA9CKj4SrwX96sWrijln5Mf8jymOGR5QFRw8FZ4QN/ldOTmg
iH+sPG9qB42c657DvRMeat0YHSkr+TvrrCPTjRA2ZAyJyraea9YguRKAfSV/9Igm
zkzx7zqea1pCKpmV8pUAzuu5qf1/HA+rcNKQfuUMaPVa7TmFVw5/BAilAMeWTL4R
HhuiB+SpbK3FLklg4xQYQno0PWu3T6ct3Vew21LwOzFDN+0Xoxqntc8u2jYvzeGp
m9Cly5rPXK54z3HECzhHw4OvpB9xedyyhSY/5Ckbbce8b7vQg18eryzCWj0Oegog
b8RiY9X1B2+FKCi12xY6ocSEW4sQUed/bm9hm+30xNw+UfPVRZ0Bt1bUkV9RygMj
5IuVpS38TPsmXRCEUg4XZQtJCL2Zo3p2SJ6IkBde5N4r0XTXk3huD9nvgamX/0z/
pB/SWudCtU03KsFZORxzTs7LuwcPJrREwqoiW9qAbCtPygw0LjxUtcfIG83vSyXk
+5n5LV1dlr2K23V0wyYfN68F8R8UqkkPlA6KHByrSYAFmWuOcgjcxgVFP4DXVFM7
lm30DQeaA5/vIbnhL5A0QPApQnAgG3pTmMYEA8knxos1ns0CwejFuMd1j0/LDEML
Brll93C+N0gQaMnAUHjjdyyWtyJlFBtfNX1LHHlon4KKNAB2DDyE8jDLmxffZj07
yP3bB0yZkOKjGxfQ/oofFCIwSKlt5p/VvNPN60ZM9c5zIkcY44MEFdk/sH+tBnuP
5t2eJ6feC3mrEUYrzA/tkftG1TOOM2yK3RfWRgVfds+GgdvuI7cCqLYa3P+pn+IZ
ATFGUQMbl2CWX+24kvZsB2+pzK0JyS/H0x68pjtLlYC83DyBv/oX4PT4bd6loqHs
sTILaQp9euL9F8bbrz90JuwaGsrOf9bbeBLAEiATyHOwNDkTcozTbJHUX+lNBfEn
yvFFa3/4Wxo0W+55swDSbXZ6+YG9oaspMXPPvphuoFHBD94dHLQ7ccmgolcVIUYz
jtd7Cd0kZIoA85H+1DZJCpUyCICSkl/qwpimSMf5xqAjieuaH3OpWxxRIGSHJtid
IbreyUuofYljdWoGGYxRpNAr+TL5v1JBwdFxFVwSA3gkJtlBWOxJR5YfgEIFCKvc
ZqGMRsNsogu4mBr80LM1ZHrVRjTrr1iqahu52L97xGID+Knktv8KH447DFAvnFfQ
PII6Au0tlw5cXi/0uaAcK+tMtLOsQfOwEXxA+z+We/TjE/+AiI/3SKvgNy2+/aAl
44NoG5qr2h75CCBa+AuilHsm6dDYnM+BcW7ZNfygLarGoIUw7bFl+HilSrdb6v4y
JlJCfNvBEFCP0GKSrwewNlnyqQXbhfAsTdw37cloNGOGWj0YWjATSyMxPFji7CUj
zIHYfhnv/hBNi1A7kb2vJPHJ0hI1dR3Vh21LKO1hmLf4zDD8z+2QjvVq49GwCYAE
1Lw2AOzLCQg37PvlMRNGIhb1KjuWhlpDoN57qHR86/F3XYvHHVKeaZaU8rcpxcQp
au0y/TPaXt/ZKdNK5ku4eoxhMGMrxpw/wmm9xvluToQpP50x0Y6/KUwVVGM9AjDJ
W1rvrpTF5vtnWy8Rl0LHrWOwQoqyLT0iHj4FGD5yUPQMhoArQbCF9f9Z3fMGBmu7
JapnfKocZKUERy366UMXvJC+lRH3aW7XjLnPgFgxIMTSakHLDqKszDMDJ0iMvEgh
HeSJZXf+sXdVStGM42h4WtUHaYsX/2zFLR2wenG47ErbmQhx2cgMSycRtC3ernbG
CIkaTHKcjcUp24he1mERjA75KMdeXf5zM8677y/v39apW8yt5/nnnpHjGkYnSQAI
uqcFnNmBbvkJfw3nWCpCpi6P1z5s5HOLmFNOH5LnN/GBhbVCboXVfKIRp2eLqQZV
plZwaHQtLVCPnpZyrXRXW5dFufgAMZv6rd9xXbMZ1NkQSuGigDfmOPTAhTaAl6uA
lJiD39N9EfAkhIdwuhkKFIOUV/1qz6+7vYzhXC1RKGHPtAltN5yWvWfXoWCYPaAH
h4K7qSBmiv6/oOe9BvFH60ZxKdiijq2CqNq+rPFBFx8zOpMiMJ29xUNMNsbmllqc
6TTIO8bLbE52LzSXMGtyP1fa6uSJIYRoXTro3BjR0vi2TYc/lxeC6lk22MEu8pZf
l/eeHi7gG/oaaZm5T88DUJKUBqcC5Jp+uMOy5ZPGO8V1R8ejDAaEvjaEporbs3vA
p9CzryouU9wren079nu1Fk0mKwsRFLKdVl/A62GFhYf4l/3PLTRteqM2vg4X2ys4
DV2BMwlIHotlyPsustx0rew8rANSqBXz32Qt+KviITcULuOf6isjyIGsS9Nu2ScD
qCn7kO3BGKtoSrh2JR5tRhsp7G8+Yy5cnujL5q3wY45fUzfC9SNcUQTjJtK/pQto
CGBtEwpXR/fZsiANvCXj9S/m3l1kkgzkncR6Vz2PZGJjTUugdhbtIrukpEORYqFD
Df1L5zW2M1TbvBJbTCUacYrVXykWaRG3eh7TNFi2c6fIi0C68VilRAL/lw2aQKXt
0hG+lEVZYNPqXi3JoFtizla29nZqYXF7kyzQKRuVqtntyyeVRLOgBzEzxH/qCNe0
gBO2jLEt1O8Z27hGN0UekA65+P1sElnnE1RVhJBXEonMn11opj9sQ2Bph52E/435
qLDSJ/ZesUeob9B5hUHPonwULseEMQ8wIom/MwV7AH/XzyQWNTSTPSUGIzktvC4t
r6onuMQiOwSAylU+NPg9YpTtaBNq/jL3z8Q1nR8sEE8zJ7ohJwRL1JYk49t/W2DA
d+4AC67WHvVoxxjuUP7U7iRkCDIpE4bpS8tWGozecsIuHF5+C1URU0Re1MY+BZwX
eUPZO6081fg/CTzwTWO9yMCUmHIykl8WG3E75Dajb9SehQsCmP6nLbMc9GJFwev0
WDiA4Hu4/laqjy+/dDkVKZ627UUYxlLMbelXC3KuQVFRJATZ565R6lOmYHqDdHa9
brabrP9MqdGcls+C04OxKGzn3VYZjyDlzw/JVdVUoNxedLUDnizG5zWB+DC8lqnw
8ZIR3QD0f4fa/f6+qZxCTLUmPCU73MxMW73D35DwmylG/XAvQ7NIRUSubXu/a5cm
fzLVS9kaHcH2u57M7ceK6Nu4OqMs7QzovToB95J7gcSsX0HxXIUkUJ2C2nQvyzbe
Z4xfOJ3L7m94vPH8jAjaqC1zR/Bz6cHD7PxbrYzctOpbtOrMCoXoV2OIHvYeo3zG
9Ac5vKx/Eev1N/t8mjnjFCc8ex6swuPJQAxtEB9clHOSXy5DFx+Y/hKSvgx1eXvO
tf2E8hbyEjFZWdvIH8PDjE4wEn0fp3mZhPtOkNZLOCanAgZwPzgSyeQA8Gx5dUIU
S1CIu3KKMfL0FOj98IHok1dLIjoaApqKQbQxaCG369hz3YYmfAc2TchP89S+mmZd
Z0aF5RBMT/1ZD6EI2B/Yfs268ilwwo3iFqrIwY9cQvkJ0PNw1jI40k03qiAhwDQr
NuE4YS95wCQUIUXcbC0yN3YT3cVuTD6nRmeyqWCnRsr8Mi3hKUn9EugAKSPpVHPK
BB0+twIwoeYj4Ee8Bfl8gRLR8a86PNpg6NQ0Iq+1SN3LrxoaCpDmyWlKslFozrCO
h3PPW7OfKXevvi4FzKDYuHqwqROL/DY34S9Ju8pRoDkEl8DQnMBkgM+xMcXoMMoW
YcSHxFo3UkVhQCa4qIeuMF/DHbuCw8dhcEF2rkPS0faNM/g8JmdhWCU5DQJtaU6C
8NqoLDKQRJdmv2sKOsUk2B+SJBP7muui6it4xwzDqJEflIxN535rFW3ZZsz+dqlZ
+miS4Csj4rm9JXcEDf/39Bq+LKqd8s+IraWyyuQiGSmqXZE/AznU2pDAUIVrofjA
suPnXVfnl73BXg0KQv07kv63bLEUaaHD380CXrIUcOylC+i6DCxc5rWBkxFW7Aaz
3DYTye+c4/KPAbb468oRzdDDMpTQcShBCzAvypiRYrZgQHJBEYaixZqscWP+4qVW
Ohvhwis5nLJxyGHSHv1DIJOKy4ND+rpviPSLXYO+ozzweJoulhNi5FnBPMtUUfH9
KpOU9B7NyrRe/Wx87sreklJUvA+RczC5U+Ct/8xl85DXmZkVX+qeD0ciG0YtEJbr
QOU9FHghsb43QtzyfR7VS5G0cXbA4rw2WuNdva1fxwy48tUnXoxY8zrzuGEFNvPR
WVT2FD9BMsq4wzVBAraKp8ltboSK9Xl3f0CCVzPQtfZp/Kz7sZ5K+VjSDcbxQepc
qU4ihr60eCDCK/hRCQ02ilRfn2sSKwBowEurP1T+I/eFqJkK/++fOLEVkGZ2AJNA
7UjcVeCidoK9EONyqupiG+TwUnK8oeZg4T5FeYwVpwxnL2wTgQFbZqeNqW3YcgV5
MrJkbLW+9izEbS+5zxkeZKLV5zV/IvKG80NxKgB5SZDfSURev0yq3YhNVRyMKvOo
K9qqkAyXtEuT/OpzZvEC2zTuNVAUKiCx/9dHQAs2ojMAxmWcKsb0Ca9DZ6S9/ek/
kygVMBB9V/6OBU/Wmb82WBbmXZyHG8T6H5IEadfoy70FQw/x/DwblXA9LsnPALIE
kRigiV8DV96dsgzoAqc29wg2ojUAAkq8NJaXxA/lLkikqzLb7l1GX2swCtKlvtwY
BWvdoCHM5x+F6Q5WOTnX5vjXW+WRCU/vZGj3aOIoLIFQbGSqCJALN60CuuCQyxos
0dN0pYZuJgbK26kjxX13Dt8Hz4OBFX5TeD1tlpj5M/lqi3tZEcTzbRroJXCUkLO9
j+l5nBLX/+eii9QnRiyS5VPwDVXiwSm7oYi1KfuuLK6VTqL/R2yEQEUb9zA5DGpV
gWXX5z7S+ue+OIgfVITltndZTUQ+dEmAWwaLBrqmqGneIU1u76Sv+/2oIapGuPtf
xvAH0CHcQKy/AtSZLJ7ssqTZ+3s6cJ1demTJa7TxZ46hx6Z0dkCBJEXO5GnbX8Oc
Du9qvZctK8XETHSy7hZwvr1B9YC68Wl4HXrpaBg7UcAfILPasHgNJWzMkQem+4Fa
T/bjsJK+KxrdGod5vrJQvihy+395wT7+QD0j9wBwIIfTV74kmIgbw4aCDAImL72H
KUDXvxpXp1A8eU059H9A0R4nnNaEKbLXXMELDpwc24jUoFhXPA33AFYw/GRbTnU9
qvuA/Aw9iyZ/H/ETsXilOEhvv3gRNVBO5pXzTaRGmRce96ldZ2zEB8OWiaULgNYv
FZ2kO8+bfXAGIhEcYuF/voSEcXZECnMjtX5R//+UawmLplGmLC+FAy+gJVK13ksG
Sj/IfnAG/e3//sck/6lV3Az5EZ2ZfRFxoJj8m10x7eIuTTyPOs8h2ap9XrYN86MC
I3jsY/FxD4mT3oEBY6TpjbgitXTCe4p8zmvLRzlGSI5RcsE+XLQEzq1TivPIeCX0
yw4JkdSQs/rXAuWGnofRBpPvzCNQlcNRzsSz2kOrzgCoBpPKBDVArlTfHDQI9esi
ubVUvW/wcbz/3gEblKeizt2V9rqRCnu7lDylZzX7AlXUBp62dHjfYVHr+svDe5Cx
grDUwLe2qQhqaDL8oQFs3J99Go+EGUwprCgfzJkoJ7P3iwWGaWcgXj11n9U5mTQO
64qZxcKY5g58UCNWgJLoX4EFcXhEnXWATp0eSeMD4LhaODexXOYVh4DgzdilUii6
GjK6PKDQzx1Z48WRuZxpZtKXv0CrphSEC8KigNCepMLbl7j5gHkUhlR2hTagzYnt
zHXSaggAJ+lhzSlefAKEhYOk3OBlvE7+vAMETCCjUAvV9hbDVksfsEYzLM0SOECv
Cp2tZ5O/ePt/E+FZdAvSlIBhsouydWWCm3aMmTewxMx6kv1bJ+de/nFSb6C5YLTq
XBgD/IYZDjuD/7/MLtL1G6uwcyKvJPfqryWF6cMe0Em0BlVXz9ly+YFZE0FbwJ3L
ySrrRwds0TPaY3g3NYvQYOF21YDmLC/9sypLxLVo+3MS2+R5Dqz6p7f6kAe4lX7w
x9Temum/8n86ZDWgfVkyH0nk816zQJJ1UbQ/Nz6rlaXsnfUrxCeoRw6yX7ayNrtI
g1EZGjFZ0u2WYFMkqQ/d1LX2M1KPcrF4X3wKfno6408y/MuHV+FRWt5+UG3VS6Od
OkTI2oBHuhLoghbN1C1OTXg5TruntHCzkmgJgfbiXRlRkCLNWdVKyFHiv1e529LL
7af0o3zh5FTvrm8Sn1iw7qz1N47qCW1si5CpJjYAMuVljawRDdsxliROKWTAC2vK
vRMUwwd1GmebfCVXnI7LZ85Pgb/58iC6xQumNkgNZBxoFV4Sf9RPHDYfyHIPEHgO
fnTwYkpOBVFwqyDPR212BdyCL6VIFR108HhXPzsvheSJAt7crFN0djBhcD2J5AS0
DWsHSiGqGBdpw4jJqHE45Gj03i/wzIxKUdeP42JLAfGZpyE4KY9k9Zt18FjYsqQm
HXQcCrY4nGP2RGSN6t+/n6MS/RG25T8HO6i3JD35yG4/zRs7IEZFgh6XTNHrJr2R
j45JHu+NxNd3mkZ227buQoQLO9e2b0xianuUoJ2SCb24tKI3yRIsz1lsB8wYCrSa
gZykphlJzch/q6O0ob2n0kQaa76q2iRMxro6Q1evt9vP/R8Gr2cwG5tsE158ikBL
txgHgq0CRtCibQAscd/QnW5sMdsCobYLmyM8JR+uBHMXKztP901vo6LdmcuRa3bk
ska3JgSL7kL6zX0CzkfzOXN1VbCWqr6GPzRqY4XgVdvf+ad1s3bBa/NFJe9m+veg
srsRlA5/fuyei+2yMQa5tFE1ObPhNVM3c7DiT0zSanOnsURIzGtAD+25Dz5UUPN/
b6AETQVLdzq+s+v5lYPWHdABL9ESZn2PHOpb4ZXQtIr7Phh16K1S6itddJAIBE81
mbxbdUqlf/vP5Xgea3F0fhiDk6v0A/K8/lrR6/hPjCsczWwdcuDbTotHqufhVfEe
KggTn0PRJsrtbtBrLimqVCVvC/1zGAC/jAGps+tvLepsN1gS6byePd8kpes5zO5E
7wkvmJg/tJlsbQc5+GngkrGhtC4U1p8rC91QByd+bpftKDgyXqyQVlb24tlWLy+6
HFb6AKPmKFa3AeUxYf9B+RRVwx9VL1xN+n1PGPp5pntqwYF7/Lk9H+dSxcQUHX0+
Y7bfGi6EZuECjOckGv3rAfOv9Sjz+h15988trR+KuVBeV411rc/nK62y6hhe/jfX
XlLce499vyqKYIZ1KO/5S22XZG1IZs6i2uRTlJEj5ieooZC0WG2LNmBFJUVVxrgv
xEC+dmhRI46q3qrdonzB6L7k1e+kAL68TMzQZ2ecRY9/IxPgENxDtT6kkuSiM5RM
qcD8HbYZn36T6tB1VykoVz+tYhmEjwbqLuEGbRFnQyZPwUhqJYHAPkncXrtUR7Ds
Pv/bFTHON45UeC4ULlrp3QXgTGSd8ElZamEi+2EcYMJ5/9KjRVdc2KMkAtuRYKMN
konCfYGScqh5gbaAlj6gcSWwnwx6md//CM3LGJDyg6N1oqOs50Xj0Ii4+SbQ20su
6VS4RC7yt+hFYd4io/BCZW4eoutDbX69TcdUhS2m3k+8Mwxnvc27JrLshQdbDd0q
BQQ+rIrvZOX1BrVzP62cmUMLjYsdRRRFTEbUqEOVHO3xWwDAtDcDj3rhHO3Co/uw
a3j4xzhAeUwBjy2Y2thbS4wpWTOJNoSuw91zx8qhKT3uH7sUxCTFB+C9n3wcZlky
1UwOBf6iKJEMaivrrVbquZqxPQ/AkpJapppivDbGnJ3zWUXfNbOte0Mtl3LWv2Qw
4sCf7lPEioKSDNOUKGGe8MZqCGSMGQ1rv54Ve4ukiLZWMhhg3MqXqfhYa4mZ6UMl
Wp+FWx/1Z4wM4IuCDu0mRYGKiTBdj8FXykPN0URVLucX1nLo0NIolj/V0kcbM7o1
qcRAG2EJUVGwbDG+E2ExNa8e0hV+AQeTsYvpaGRSsTrF1iQAkrb0OoAR1bBUn9qP
4Blc+qLmIQlIfnI+qqrV/bC8yXylhaxIFBoCKn3BXl/ldgwDkzoJBFYr9A67uNyd
sWhy3lyBog/fucFQs3hAyotBzof5HRr4206Vb8YTjsScPjUMZNUdBYV32v09ntBJ
lXBUJ99dJoxL5m3eIVsshHwcVjkGHlJdZ/EXL+EPjoyyOraYvnWCz9AIrJ5XO8rT
hypeYt7Tqz/s/6pq4mcock+GYjZ6HrqxmnaH6tj+vFwJhlvsK3dr5BjvhyGFbD9A
1B7A0Mwz76ui2EcavHKzFbEXN6qAX98VoMvicKzIiRp5Wi42D5Tgv4Y0/uL1HRj8
yiDlYHA1gC0wfAKyViTun/bk3/HLq4+MwL3kk8F40jg7J7HsVy+TH6X8BQGwnxc7
VxxzIK8e9CdHZn6H7Usya0fyTrcZRgkXdV5Nqe4Zb0PobyXbQ2RQmVyUYthGPfZC
goeULOiXYLbaQe74FZu/ISrd4m2cNuMTh+c/i1rKWgqWIYOwLF8jjh/MpW8LR31B
ZkfBU3GIGAJeGUj2ds5cps2UthmqxBrHtFsVZH5dlgWdh5C9Zx8TS1+RjIhPhvje
b+3Yom8bViIAxTdY+imXRex0fyF2p+h+Ge8liy+yCsGL6Wv3Wa+ZWIy8lkcKzfjI
SF/KfgLJu9ooZLj0VTWIX58AtZY76SF/rI0WBd7VH7b80DYBHVf7BW4PTn37bm60
5IsT2f3fph303F91yk5CixzeUagaYq+kEyo+hlnX4vE3kdVroQtTwcfLtJUiJVnz
xaUK1vfCdtHVEmw3Glvl2Xi3soqLKInZpqK2p+fvTqsJbCv5VYMZV1WsU2g7xVOe
2+JERYRgLfU0zs9ShvqUvj6PwN+V2BVVhEN1ZMB8rcDC4wdk6d984zKXbfIB31tu
k6CNkGgiv4nGorrizjeAv+Cm6ecJjIC/z0wCqIi1PX6PGvowtRd5BT6OAjmuLw8I
GQY1wWNx5aylKAqSjuML7iNpTtDzGnRH+ytijHONL13NC3ATuwNkXrY1JfVVu1G3
bbtH3VVAn9V5zE5oCH/iJBVfZF6zmwL6suyt9/chwwUqnpcAviqjCxRvxutRR+VM
PQ4J+Y7hkGq16AumYqGtYhJ7Pu9j6DGpxIza66TQ15s3d1yAIK8FlOUAKBGzoPX0
UadJ0Uqm4V7u+nE/8t7hZSIewPtd/DQ6Pg69aOXK+n5t8nCh2ehso6oT9WDgvZWU
0o6O1lRMtKfd/w/LbHcjNSE1BehblQgtoJ3q/cwcpyQ7PjYxZ55Lo/O+eXooVm1n
qMDjfgt/gsX3Zsnk7zltAqZ3X2bMtomeDcHfthMI85fbS6+4ZF0PSxTLhpEcibwr
1UXyQC/KHJTM8IXwAziMTPWktMqCRBRUPu+l3WiAIsCi2xQAB1PFTa3eK4lB1LSM
KkemLrSxvBumrhCAWPE3jSU4g/kQX9an6Y/wx/F506vG/pP10+w3mNCt5YEnvT0u
yQGiJs+OYxbio63SywbxO9X2/yP0DjuVe3qSVyQmIwdODTp6Vrf9/jWIeuylVbip
+NY+xTmOq6LAVPr4mHXYrqxqRaIrYwfe5awIpELjJ3+bDHU+hlBjNZ55zKTj7Xr8
zhwTXlRbtkdB2cHqZdCqHHgfZY7U7N+9tVCW+QpfGgrishwkmJjg2nxxcltX53jm
Auj83CIUzPvPj1PTIl2FKzcs069hQ5WtvD8M5sZLGFUAQBmvdR/1R5/xPMozxP1d
reXRZXIV6U/ShUxPOmA/GnDijxJAcJ2EYhkk4bq0vFW1kFy+Ys66PZyrau7yxq0Y
/vGbK+iR1GXRd26xssQikLEuh8AgRZioolGkBcslmDA9FkX9AULJKn5Sru4W0KTQ
r76tbsalUZcZhcnvKUiiNkImfShsAo417gXlK9dPofsTgZf+wG2MXztRGjtHkncQ
4lYmoSdCtqL64X7q7DODjz6z+66gZsK0+2zi99mCYEmjju1gS8ei916NyMg1R4Bd
OojjZczP24nIJ2MkPRu8W4WSSSb0l1cbk/EL8f/7kEaAyGDzv7VZXY7nO14Ux5lE
rT//hN/5EDgeyW5vKNSr4z9shPqGlj26kC7ASkKEJinyopB7HlMmmmVukyiTKSFO
4xDNoYD3EP6C+uS1mGlJdxh0lRkgqmGKOckGM4c03y1emRQ9+R58scRL7TnLR03D
wO9b8EfqfleGa8TTuqT7d2NJHc1rSlT8znzl6ZhVu5JypPo7hwJ9uMMbmCTbirc/
8C1enAWJ6SRzuYBVQj+o19fju+fglSOLJk6J93PeyqxfRDHo2hu+zX2A95Dyqnhf
lTulo6iafWG2O/rXd5RNxYF8kT5+EDytohMjs7YyneDKE78vRQY0e5zxVw4AaKcV
RPbzacFzIXEg7SoBDH7SxIqj9bf19vtF2kG6KJPQ5eGUdTEH3RRlAxAzToRHRQ8b
L7cOWWXFxKHx4TsBKvKCZy9Z/aLUJr9avQtWYNSmNZIk35MpUzblPwtWGZel/02n
gq2uQLotLeleAVAeaN2VZ1wOjYpnd34yCVJSpVf0lsxA1Xk6kK9v+XcAmLbIV7df
EpD6V8V3iyXn6zjUju7xGdrEuvs4O1XRiRHFJEgpBt5iCQmk7icl6uLr7ygy07FQ
ZIulIe9vwhUV1KhtPPedxnipO/+FJbjSvDv1xTk1i2tL8TEQnkXMOHRAPEagsrCw
UAYYp0v0QHDWMXz7CTPLtUlVRWdrpeILaHKbXY1RGHQ9pNvokiXv0XBV/EVyslj/
AtH5/e7U5cR8yRa8lFa51tRRIFJ+dCrc+gsJve6eETFsm0NF99/8DmFjWcSg1mZI
qa5IE4UP9I/uH5Ms91TgWv0dBFjs6NgiQrTtkfyz44HIbghERXZfKbJ3pS4ChNNX
0/f/iErjaxEfQd4VT4yVwo+tdrb6oUcOfOld548KmPZgiAQn3zxVycPAfJ3lTTxB
gF5CucF50CMsr76WzyMttJ+yHAf4o4NuhGUOiJbfWaT1yZyfyceGG4P6MUWRU5nO
RP7vvNWnEIzGUb6O5ZXKK+G7diI615NOe5sqvWohvsWoxHcagQnJYlo5w3aSVI3d
xHslyM3MUa8kATz9WXCOLB3w/gXhMNjH/lN//hDj+cnlWhgVKri9qAHMzLeaMbaw
qys17AvEJdcDLSm50nhHYsp0popHNv8BIe76naUpjDg4ezLt9PzZlfTBFupmXxgc
q+mP2+47ojVs6M4C6cL86O03BH+cXb2tLOlIv2MKH8j5fcsgaBnhaLk5yWPdp8+A
JgD1ej7WPVYkFcvlIYa/6QR7YW0YU+77IB1WSfblVUv/L/SQVU893GrQtomjPgKo
0RWGI5jw9egv9wWqPB7x5g4wx5a8tukOTU5M9KAsLZHdZOfy95CZ1qZPVtq+Ih5a
sVpcML99qnjCjqfSrV4UY9zHkUYm2qQ+yhVYgLsGqd2gIhuWizAP1jkPqnvR6sGu
PFSkmB7wdCNheJf8Rj3roZY2UbUgHgtWUZLC9bGDU3ksgKh+6Kxu4rxnd96WJjhP
W4rE9/KeGxwkrkLEeJSCPrG94Pu6kEh7KVTJA34TEMGqqNk2LTmlZYmAT6Kx3eeM
X7kNZw0XAi6qj8HB3mAAE+BpgPgkZn1pyZX5SCbzwKMStt8GvFs1haj3Jyn0qpE4
yVsCNoySS5ho0rCckBH1bVabcsNDbsXkR4aTXx2xCZ0c8F8UQJ8mD/UplNkqSs/b
Jar2d++gruv62Y7pO4rQB0N+R9qR07UYKFqWvKcWSkYkG0sq9o16C5+5BEzcQkUk
7j8i49tRr4SWSyQEQc5KZVmJQwkqT8clEDXBrnBGKnwoTWGw2XPRqAI5MNPQtN5w
cv4TJ1ofZsJXwebfs5B6NfS8dTXPKZY+DMqEnli77VddSfx8OoiPTnczkmGnT0St
dMQ5wkTH0OT9Yq1Uu9GS3pINtlZdAHcXxFGKu6bEBFozZZYzBNiv9XMuWoeG3YG5
4wZUhIaD1XIGKNh8/c6mVTdGexOvLCUe7BWpB0gg/EPJdmD8pHFMWFuKoyAWgTw6
Oh6lYd9lACDEbuc+dihzoHFR6HOOPsKmADH/AQxTTnhOkkfrUgeKnQ7TGyfbQBua
tuQelk+ydGPQ4EDwxLZ8rrxdBaV3Sm0yutxAW+MCr7ZJHnN484QW7fjRQrnApZJs
KlW2AVlnEjTHqt95bPPaF1GCewFUPUhZnbKOp7CM+y0gstYZIhzXw2Tapcz7WSOR
5y1Xb8VrZn96mrFSWoCbhT2QTZaqR5wGe0PkCQEtzedKRXU9eur6YXAmhSAHU5vB
Tqs36jtqP6jewltAa3biImAk32nwd8885WUcuIFhrECualfcv/U18y8uCCAJYmKd
z+fIPJDK40+TOlIdinABISRwLQ5jVrD28bVP8Y5tDwJoN3c+oQFac0CvDokg6Cu/
5Zdztx5DQW4UPYmI3Fem0fNqW2Mnfd/yA4YcHBEzCYGC5BKQKdUrPU2JKCiCxD4x
BmkPR4yHK5a5ycig0xsm7Alu2fSDgquOCZCGzbPjcnIaxBkWgPtUMKcRLvjlV352
tAOX7ZbplJla51WdU2nCMajRQohPM6uZ+10uCZu0MLg0C9MaSs0txphUTs5WZTuM
iarmmA/bSE5ukp4v5h/b7jfFCJTmnvSiL6NLwACg/IYGtFvLV/5eC5y6mZ+b00co
5kTPRyw6znP+ricoaDJr3CaLkIy+IVFN8aNlYlZMxUHwqi5f/dBmj1k41dAQJZYz
WnYyWVvlWK9JQDzMqvJs8lek5yxEJapD1RqC+kBC30EESdKRehfLwqHMkXYvUWy0
ANNTngbx2r3NJBpN1+KXxQAidzC6iocsF7HG+dk+6e4xzpQecH8NXk+A+M36j7bk
l3b5B+P9gFhPH37Usolqm+WsiFx0b4WZ/uCUx9EtuZvlAVUK8apvWCUabE2n7noi
xqT3JQ8LQjZaML4iZ71jS3YU1rzrJ36CTZXwCWt2CBXSvKdisvBAGvIo/B9H1z9z
Pa3TeS+43AKtQBX/cj4Bgwf5Kmrh1a10QDBM80z2DvQUp10kWMiB5IcMNZZh06pq
POrWLrYQsC/pKYBlqTO6FPrjgQsn59jsCUOn5gNvjwNAQfws7L8eIMx4YArj3vcD
5JRukJVp5SOgsNxZ19nhaosxWh5Lh2vqOipMKDIBIzCiIQ3qZkzfXTyn7n77yE5k
U9HwA4orQOdBPIkAd1W9Rn/OKk51HSIcCRuoDXZRPnseM3VbIAta3qdlfjwmK3Du
TD/N6FJwM/EX27HOUZIq8uGTB0JWwgh9cKa+1UENN4V3A4cZliMrVBjOp2bnZ9EG
IACTjrYwDoMpEPBktav1MHed2JJDfm44frs1AYqFgq/SOhdEIjMWjPJCxgwOPuyj
l2M89rVjO3u8iFpGpx6VJ1TlNapT/azb1TbnJ6QzRVQdItFEDRRMCKHTwRC/Zgzp
HqKKtddjcHkgurYkvbdJ7gizFtZwvo1Y6+kZksKNrsPP+8keD9+0K5FgoJe4z/QA
DKGdBmM0Su2G4sTpgpntKuyzPd65LQ3O3QaAUzQ7eNy+LioWP2yRC4+f7sZj8FL3
0pyTcnlXmKNvEo3lT6Ql1EI1yAiDkzKHSbUfcdTpartjjLMDjlUSqw2XmAqsUR4N
pxduaU3I8qPbjrhpGdPpNhGCZQ66+SsfGPdnOZ8dnCy9ejr0pwcoiT+8ocjFM3Tr
iSoSsOeKZKHF7wq+q4k883fEZl/s7UbY3RPgts6OmRMqES5TW0ugium0gkpT5wme
1wA6cJ79jBa00etTSAj+S7WnpHph+VlExnmYQgnQCUuvpBnhLk0rz8mLCeOhpIUp
T510n91gnTXS7yT4ZxjK5g==
`protect end_protected