`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
K1W7uuA+c2p+j1DoODqY++P+/YtfLyhXpeXPJVL9NCocmHmzHSnOMvJ8d39fD+OM
2Nop4nv0zMn/K+550rtBQggVvD2bdtClfOFrBb6fX1lwV96pH3hcZ8sgvuTgWOwp
L7MRxFi+hOHdR3tKQW5vOqQxKHvKAHDQQuglgOOo7nifO/oJeJ+ZpTVchuZ6laPK
aQMMC8cR8wCOoRBfws0sSv53+5JvEgZyWmFzXQhne9oeVzBnZOf3+S2gQPy4FWc6
yaGsYeNao7Z9VPqq0ynSA8bpGVvJ0X6mR4IHOYy40qkwiliw2HY0ETmN+NiuZAks
cQtYCC8yoRxDD0LJRHj/JPPCdeauD6wUaAf9bwUDr3JkdysWkL6M/2jchYK2txqy
2gOq94MLljsmJDwKzOkUvcxTRGnHE497yAa9rEq7wgLKIDfyKnnFYIee1acLxoZi
C6RFjNbYWbtgFjQ/HgXNAIX0DUDn8hZO5c2FqFQhdqM6lUPZ5J1eYxkFfA/lExcx
rneW3XlBf8y2JXb62p+1I2f1JrYFbHvGC5Bpy40YYan81P7kJGqMkTKmB//g2BMa
4OdmEY4DdRKlJ8TrtRZBZYSoQk+r0AwBFkGyvLjiMdqSOFFxhqkVG17DOKQR9mtH
V/yvXb0Y7Jd8flh68vV9NqEwbrkTuSpvPLDhxPNFerEgIIO6dE3YFlPQKVPyYGmf
HUtm8yZeQ/0A5VRlCdjttg9r5eVma0dcK2VSlY/aRhJR7974IfY1WADKlKBnaBD1
EBPCB+WBeo2nvA3vq7rgkc5CF+PNAqALfnTmZ8q2d/ctyaTBhhRWrmBlTkFldiwY
S5/slsKumkVx+gWPHiRPuuuPKisxb6kLLZHOIQlCtNe5ARnfpuRTqkxYbFWnqYm3
OJbViKjheOWZInkNqxUc3AG6qrgMADBfNAzvnBN8AUe0OcPcfwCS9BYZw3sMJreo
hPf36WzkNGaFc2psQcVveaSLOGHGn7IBL1jOdf2BOGQyXmk7BE6HtuFoDQIRkt73
Hz4pvkrt0cTUys3fPKLm31Vi83+LUMG9ZKJGuTP6vPEzlN4Wf9JsAXlC9H12/Geq
drB+VBbb8yrL5vGRgWWWD5/ltiH0JDGaVugLulKAbqSLQKHwIZGku1aixO5GCI2b
NcLH2sMa8Xm04of75tgqXSk1y6OgulCDoUW9LPK49uvZbIPaESzowWxI6bTcJHHw
XV31rhHE1kZh23qBgeJQ9GExV8AH7og5hw22XkH5w/IqgAeaXOAFwi700QNDKOfX
heklzNbDCqKMP7IOtZwgUPEOmJDuEDczw66teJfMiP+I7l5HZOocvlnxVvtby2rj
CmOSJuGB8ZTRqFSlIYXufuPfV1rkM2BFoA+5JsCCIDrTOPRbEilVvb+1idjAF2Ci
P5Ka6d5175yAOuRCm19dQaPO96Cj7vdc48M8yB1f4iSovrMk4ZdH9fupQl4rQEgN
OT7bZOVKmVlXJNL6MEV6msyGwjW2/WzCZUkdkea/j4GQ90BUWvw5ZmKwsItr+3M+
1W+332ZXl1gE04gVbXeZGvKcUkoxom7N3vFPjRUctUDl40rgcDM71vh2MJbxSXKf
yGuQ6krgfs9XXTVTZIR3Oun5VUVmp8QkU5TAVZjau2uCqWI+FlcEmlTydzu3Kuie
rEfU5u0FmUWtfFHzbEG/znoMfUdOT1dGc97ZK9KOfTHBaLbf/sJY48iRGvkdZqII
2O7d7MY7qqDC7BJFWVm934jUxr3KF6jKADMENGbwmZaApk1LWnI0L8gh2qJe0cvP
BtFPiO4dVTmsqa6zsLwBplbIdnmJvK6rj/5cx/+2U2Z87TIcBbuhCX+90aW9wCwB
6y7b1dzejUwQZX5rPxsf8At6Pe5okjksbabZvH1/RZjEjv3Qw+QRXewRJ1HkC5Aj
sJOei/ePpRLNy1y5b5n19SXN8qAX9Ll/VK3jioTlN9Dr5+b0p7Br544UxToxYXQd
dwVOg6H4NPDaqd5XJZQNfkwytKLCILJNMbJBEvrJpn+7SyqX27gLOvL8VxiV1DsK
R9tynjWgCMS2csbAEDN8pvPTv53Z7qKpWAKGOkSAs7ElGG7mmeH+kcmnll/0ORU4
6ZIyJih6qcVrCcD5t6/Sp5pAnbFks0d+1ajqZTV3U5D5YSrl8pwoHXeXwUbF0agL
nxMvwYUisCK6ZREM3p38LIn3s+POIHDp8vs0nUf25IfOurxzTRaFmw0zmtSxWe8m
jHLHTdKlU8ixKWCdHcBYUkTbnZWkyXjNbbUsSBh+BDdaU+bSMbwxstxks4mTCGSw
BkX58C7/WRDJU+fxsFCCwBcwX9036LTCPO/bmgcDAVmF+3uZ32BVc2lk8BYEM1sv
+ex4fdcdp9460IaJ/xubkaTbJWTEyENl3J730J8HNrNpMbzVb+O+/l+0ijrFAO7R
I5mJuO/T5OoxyiRZYn4S8HwFjGkJfW2hRIVFy0ICTXcGq19JkfnWd5rwtGb79LAv
6iVJfDGjbMVa2VRTYSqM/8pL7aPI7WEABG2xnbYkh0aziplB3EBBTVl2DmhSfM6P
mBbriwGDhSzRAy1ieybUYWf9qk4Gc6jAlsPVg4hYqNWvw/c2Z2xaMoEMXWHpFIdC
iW1mUrFi7yKl2Qo+06JKeansppkvFu1p3ijmoCYO9GoJdjQXzIWIGc5Ge/LklP8b
+idU3vHB9kgtLu0T2U0CIMg879ApL/ScRyi4BHp50MAsGeC8U7F+6Zl4rZh5tE6j
5m8MSQSq5wYCwyebNusR+8tVaf4r/nSyCGe1e4uJGg++w+sBQ7Icr11G4a7ZKfC2
ilt+7Cf/a+FFlz+gMWwA5TB5I7pBD3xasT2mJRMRtu540BCg+USL3B/xn7mLzHKl
cjVcL9K1MWN4TslMr3uCQ0YJtryP99i4GuWXNCzlX8scShCjt/QxPHYzvh7tpnV3
g2LbiXW9F9CbkvrRZw5kA7fvGFnbOVmSooYNrXXESupbdhhPF86AbIQZwn13Fy5c
paRaSCUKbU6DSz4mmeb0anIoZRVBoc1r+0N4Q/8DXKW/T30FvgK4qNoP+rtRura5
TM8au+MkdyjYy+Nzh2V9EZqgM/ztT1FlNR2daE939qdH9J3QfWYqY+7BNphZmB/C
UK9hugkpK33RHXEkJAaTRZ/gCurq/1Ea9UNoZKYIevbViUBPQwFCXvdN8AUOsXfG
uQs+AifwZropL6y3FH9QLAfdDuTB77BCSCGST+dosYRzSk4Vkk71O57wwj8U7bFW
RTGl4rA7W4f8/DYu4z+/2lCKwiJRh6EIVihRR3kLe3KFeseM9i8fP8p5AZljbOro
r+HabolyjxrflqDiWjyqIRRMmovIn5gznhvr6CDHZzQ6CW/iyN01kJoy09DbktLP
yyrbNIHkKQErCbIacAq/+cBlxk8+W2N1QXdpx14DSKQ7dRrikZISkJ86Y4jW2kcL
YI8H5aa+xKvgzRpnqMHPCStRG5vnwRRUiVE/L1bl9QnvG7r4dEWNziG/JFti5+lF
aiq7zBJhIz6QCQwP/LwFtW03SToc8zOtpE+IuCpJ6AqV/tmgTxcvkNgMCxewFgjd
lJHnV63xR61cyw/FXdKXlLZ3yAe4XW1SWbGvlO6jdL0yR2p/+ZeE7dkwHI62T/XI
h8OuWL7MEcGk0AK7pk9nlakpey6xsFH3YofNuj6YgG9s68DtPHVtS2oN4blTR/OH
xe583tryarriGPr49JImTL4neTmBGzLvYQc3KSlvRgQ+Oe4/aJPrQGej6j2nWZMG
YnfbOufZ7Sd+19xXN6of+vofPinMarY7xrY9e+uTwSVfL34sZ1r1XZ4WCTP1tuHs
iZkHmJFC2BvfndbW63+0ghw81w84IOqd/ev6KTsyV3544/zJbQDCXWHY8FRSYAXh
u1N5uBAI/PSPTbnvF4W1V6vLFTeb577MvVslwfihO+16b36mHR8bTwfrCX8ceQEN
JG9dXp67agJHSgC61F1fWRMCDnd1lp7pjJrCbIpG63gA3HqyGdL/fhrnmjnmB4py
UYrawp0xQeIoeZaO50QySd+bPv+p/nGnBPhIcgIwVIPGQWBf1PMqSNM9L6SjF+BI
4TUB9P5auM8/0iY7W6+WTC6O73bHv+aKvKer/5sK+SWX2XFD29qzQ5zJWGh1Y4zO
QM+FHRCcwuGctxg3BmU/m4iNbKILeyTlJDuWzIreMZKorW57b4mkjo38EvNGp52U
LSDjrrbhBFZB+jWrI1hp1zJK9tp+s5h5h49E/VvLNzX4gGJ6DRT5z1kQVchqL4uB
pCSCzklobCH7h4aATjP86qrlDNImezesWg8BTfnXd86APfCHLaXRnILA7CQV3b6a
ZgWVhkjgw0dlsX//uSkLq0qiqyHhDzrnN3W2OaXbx+5Nel9zhBtVWAbxmQo0hv7K
s7PO01R2iDKpPAWT1AYbr++7FDUmKLGVuoFfFTuRDSCxZjmTvNjvh0Pmkz/cQIAH
mSHdyBEUMPIgjFS4CLa6aQWbYOKTnckyKpNXTNjFiuWq9ys9XbwSquY/VpEUbHJm
OFwYPZYQ0iXge8lP1HqmyM8sNw+sF7DJQDN83unXHfTf7nLOQ+EkzNWc9Fpr5vHh
J8o5LiaYBJcXQ3Di0Q508G+qPCel5tRS2NGFKXU1oYjrlVwLv/ICI7Fxjae3Uf6O
MZcuAnwjkQLA8vq4ya9dqdmhdS+OsGEspQwTTsO4+3tAa4UlivUag1N9zLI08H0n
8d5A1ZQ4Fyr0gRqkD82gJnFHrqiWCZfdnDqTdhc2sGN9ElVCgfRqDSit39Nlif2a
gKEPtq7/rSBF8Vqva/ld8Gi/r57lYQqrp98kuus56Sv1qrPOqd3ff3lVWXeG/uxd
K/BGWu4AYStTqYhYxzBgwkHZjIgb925TNfTKluTvlMr6tEv4CsOhVqkQS2Uula91
qYmd9GYerd3+mNKqg1slry1Kk280m0/ZncenphI8Op5nxJ9pcnhdbB2xHRwEeAZ6
399W5bAJpaG3NxJ297c59MEItBTREKSTwUVrQt5hAqqhzFm5Q+dl1PFd4t8cxvp5
yTxmYPIIbC5aTFZ9He2efVNMQlgKUJl8lcYX88HrEIdAPerDP8KkmCTLSrGIkgGM
O5tNZLLj2yU4AwRqtPKfraz3JOE3aea5bc9hUiCEWUd1aNSCOQJMveu5Okp0bSqR
GkfaxcBj5u5PGuqG//PVmfwVww/WxLQ3FNp4wytTtzgJeS5Cks18eyK6hwXa2XrT
bcbUGdqtKOxkS2cBq8d28Uo1ul1ExT+Edq2i8ZaqhiSqlokvVFkFhv5gTPWS/FGZ
9BsiHkwUSuTJEVr2Ikfs49Rv/uLytlB61v5OXAyY6k38dezWohWTpNRIYXgGSPr0
q7P5Aq4XRAsU+g0F5qB4Af/HPCP5+Ajz0OlloQ+3/YWPjZYIRnPzK+cXxH9tyGfw
7YeA0bH1l7pTGlvDs8lZZgdHxN76lZ+pNh4bN+1z0N4JBpbG2Q5ZlnYyRQBas33f
/YRJYQpNBVly74fY08r/9Lothgfpy6KxqEsUexO3alt2qUSrUzKbH7HTzsT0zj7Y
Mqa6Xq4r5XJO/xNNcyIccdHWcTbdUXLzw6yHUCKaSZJ4y3ryptEgYnbCg5SVYwxw
s9mz1Xl+70g7cCk9rvu9euguws1UnhqegyWpvFRPZNJhj4kYjb4wlBBnKHMpyoBX
BKDAIbLjnrNuvBLHCUpm1i/+geJHXOUcYvYKsu4j1ijORJBUkkhKjNmFeLNFL+NP
ivWHjB4TIrpEvMnzz3Fb4QT1ZcdtPrKqy98mIDrCmhajdtiAmx3OSO70rpUUkyJ4
ZUMRgHaqL1mcOl4ZrNZW8DwxssEbZkZNJRZ/VNHY5L30RgDZLkzpfvtUlW/Iq8Kx
+vinIpf8PFTW4ABbJuoU3p5IBkiKJUfc/SmPRNozWWKIT72M1BiHli+DhXUX9Gyw
QV3a6zEpVOVhHfIHN5mfZgMljEalRPEsKCnfIYlReCjrZYAcUJDCQlbPMDQrSzS9
UZVIh1tDUfqYBOzPr6084ZSsdc3K5OX50WnWroGoek/cLcVsM8dcStZ/7jX7JXzw
OpK31yL04kSbBnkqov49v2uLonVB0BWgZoOTzbWCtVF4jDIX8c11kPwA2h5WmL1M
1pnUlUT6v1yZZo098bX0ldbi9bAoKwWrASTumzFHlo8lIsXhLVrjXMwcHeIxX86D
jb4QDka51PM1+inf8S0OKF1uBIry26ag1+gZPUtm77937CJi1h+No/VaN8hMoAuN
2M8R3MSCAmfr/OZG+oOaXk+v5znMNjJjhRVY/FwRmYSvtx1zrPuk5VR9/G0thnpO
OmdsvmSaZuEg7sI45WPrBT7fau8jvR35LFMF4gMeRcZTn2u6t8k/4FTcgxVFtxqw
lgGbbniwWlOuFG2NvYS3vvj2QlYjTsj3eZSZNyfk0F41HFTpJBPsWgZBMJ8QQAQZ
Q57w9DY710nZQU91ZGUeh4PMS+yrXYq2/EbgC1biOZ6Z/vvGk9XmwhybZxsxppEs
Nb/LHNAhyzrWd+3gLnYzIMbQtLYK8FAAEX1s3XVHrSkNyvEUWBMmPzMYbNS1OQfD
gUTtN5q5QEknfM7gMyVhoHv2oo9BZcyg+0GFlFfD30ly76sRzFy9QbeJB92mOjeA
5yEmm/oUFMxHAAhz15NQNx4Z12nVGsc7iE2ww5dHyGxzHVDGsfcBpb8WCJFYxTOI
VbmvUU2Y+yWmanwQ5XMXMcwUjbppvyfke/rRwHE3g+v+4cMSuL0QOukcKeNujypJ
MDdUz0h41e5NovKqrwrX4yEPpPDYlnQ/AsF9JNJ0hZ4xbU/EZyeWVcr+GCmFaMcb
+l/bpBD+1M4rbrN6YUeGE/ADeH/iQkAkp1H3CeQQgFrmM3w8swAb/Ol1n/Pr2jTj
QPlvOcndTWkkVsmKQ1q74N/BfnIX9VWuOUbip9AEGqdDseLKO6G43TJkoU28flnI
UctiTN7LuXgLyDrCyblM28eipGbXA6qdHeF43QwANhZv9uLOwVGwS9JVx5EKDdN0
w39hmuQ3xjDPMufHSe6WiY92AbfhPRYKsuSdFQ65pCovrz1p+sGWZYPEnlS5K0r3
IiOxaAqxNjZRNQ5qWCgO7a2GQCJZnrx+z4OayuKlYTx/u0Www7sEuGbPniWido1c
Ml9menBFiktzuMgOTrLKs0qHiOM24MpPyJULaP8W7bDsskEgjACVx7Jfejs4F1uZ
uVNysbOe10cHZa4Ll3F3usVESpviBxyfdDC26dWYQ5z9zjUVyhn70N9fs7606ZvC
7/r9BfsSaHerK0kFufMTjdlxaCKjsze90GOl3UxTBOW/vwoavO7alYxwgKS9dOML
54wQ3OxKmwc/vGep+4FwqhomMTa9A+gMXse8QdWLie8ghvq9Rzdn9SYNfxtxA0nK
IF+37/Un4dC+C99v+NMCldXkPysjSgo/2uWCMts5GA7fNJTKj6x9frzktyyEptp8
5SkY+00veM0QDUIN/+h1jwFdkYYCyHXUntK7XxmZb4KrzEsIv5VXFkfrhwwLBMPe
F7VIPCxgzh97oFSMi1BN6msHYDtV4v1r5yX0kZ3VaXPjoieh9cX7nFGCJ7L0BEEP
8cn2G4dqD7DHmCrRgRlJEOtyoOfKBwZCxTdy5TjPNXqXK4Ycj1v1WXbqVlNH29Bs
D2o/JQ0f/blajuHm7dlLdldBAeKetomaUZqUqyAKOkJ3xaKHYipBfqhgpNwv5qg5
rTppTKWE4ATySmgHj5fOZNOciaXXYonzLakmUtGzk3mLX+aZcaEuJG6lVHrEA/ba
xCnGPl1aFCFz/MZhAOh23/5ezUdr29+rbt7lfbPYscXSgBNhf+GIg33wOVJoDk5Z
XHT3qd030gXgGjgZx0ynVCwZAFYGAJtooYZOudZNVhLukdjACJlU1Db0+q1Snr0q
HHb0Ct5XWLL7RaKe8rwad8pbrjt0BxSBWSXHr+maCk/yJFFlfHBKyCh/aiyMZ40/
sOS8D6lYK2F6JjffOjqSIAYnnCF0o3Xp6fAgvADk//0GZfSP/2uPwgwi8glJFA7o
60tWdt8LOCPFLDfVoI/PIkf+IAS3a/p7XBSXJNddBT6+5XOMBGKz+bApJRY+OigT
n1GbU0nnc/0P3hIyl02ePNnoGODhJSewxIk9H3kbcGU+DauEGy1M/vO3BcfLdiAF
ongRQ2UTl8faR6VgxHuTphrRoL8mhKfA7uazJFHQfExk1dA9VN9Ica5TTH1TjrCY
DfqkE1xj+BveGqv1Dpf1x49pS5piIghLXdfq435ctGqTr+ib/iU9q41hm81w8RkG
OMMyYcHk4iSxiQaIx7GWsCAN8oAP7dXu+3foox/4aTIt5El7NIDJ9hzluw1iN+Rj
Dr9ufZBWIXw34R2ZIxMZ5EuuSF34ij623xC/aAstghGw+lppdo3JuqGTR7NwwgHG
AMKuRKdkLkdHMno41KwsFss6QEsYBu9LhnCtinoY/JVm6ErlxVPCA0vDsDX+okoT
yhNAbUDHchovOQhRvO0GeZFkvPT0AVwCuUHkMQppQk7UPNMZC8tqnbZrgcYNX3ZG
6SUmQuRm4Rl3OaVIoyOXR0uu8XsMU+jOx8IxwdOVx+1p/YLFaraio4Wf7Pd1JjOG
msHKIe6rYJT8+pWx2QE1yMUvYH3NmdTV4DxaakvDdd63R0TG9HNO32jlNbQFlCEp
N9UL8MhGyFa26cQhbPYJI2FfTDib0H8ZIHjVSaOjzNXFz6U7cTL+zfy2gJoik+7z
B9MLvVG/flGsyNZ4pWZjhXlXqHqmspMy9iNCDu7gC/gEXGF0q+1Wvq1HPQ/Ib1c2
c5nNUnjvSwjWX9PdXhEEDwJHMyIAVxwzrpYMwgMvU6XWfwfBcCbaDz7mNVnVc+wt
htZ/eeK+8ItoACOENZVE2Ddh8M7sFsImlm5DjSAXjwiAumy4ASGupXPjMO94UoIL
24SOBWNRdrmtJ1A2dMBnP++pwgqpc4PmTxGC+4tWzpDxc5yQbq6jCcZaym5e9nVl
7BWWK5RWGJF2+FytGyX/OY4GcpEhI/EOUbw+qnTAQNgTsDtGeQsx3MslAaRCqkYb
5NmxF1stMjTjXlamiVvJ9xRylPuOBB4y/sZ4SDIP2B/z+XSlVFC1ChLcbfqxO6W9
HvZnQvKiG2i7G/OiX6b+RFN9MMnVKnHetTmG/jF+c9T3vft0qGsECZ0ydsiW99rE
xdEB5YNCXX7vW4v9UHc0gI613TjosKjUStJI2ls5RiwVBiUkd+bSJUZPZzoSLf5m
N3jtgeZlqR42sExRb1my1Kh/Le5US2uPY9hC5O+CG/3NjeYJyELWp4iS/oykLgFX
x5UqZR6iqtD+zcLstypFrVYR8uMz/E1Ui23BMUHDN0hfzp81jedH1+3+pDFHAmZH
lEGWMd6ZUhlKSqKNb8hsezHWQRjR7GMpileuumEAe2PcLOiCTIsO3YwsyXxF5EGK
67i0+pipYSBADdDyL92HndLDpxqevusUQw7zhloyKnwHAwxyoBeRO9Vjryem8Ea9
v2m9CpJXS41g/d122Xtyk7/KM6xjcNHaVtxeCOZq+3djQWFhsktrRvz1ULQ7fW+Y
/Yq/46AkpKcx0Ng5NhJrNWnA4EsoaDgrIslepVOZxJM6CTzD4BnMswH3SUCE0uKS
Tv3AojOi5qNp1uQruZWkvuTZ9JGLK/60EuXDclPS+rjmaMDJ/3W4jVvKlfx4LAt3
vxYqT5VknUjP7Cw3GGO1KtaDY5IdPlPDJSdtNkoXldN7oM+W5hAKmZ7L8Q/KgNU/
UQkoBgVD2ejsRHXkqOA+IRVXUtNVJw67dpjWQdwtmFmHpVus3EyblB+pTOUdZl3I
3DXpOKnZCkF3paqlVnUO4MPz1wzrhZdhhhM+u97DWEYX505GVWkqxH8TguZ3EOKT
vtSJmdWgTsBP6ezlAMInTwY+xv127bNZU/XIuWb1uhKmZk8VBIf2lAuPGc/ZUxFU
tSbVCiYvjhnXDkI7j9z/MhbwLacAX+t2GZzAxWg+A/xv3XBp2qYfErf9mr38Myxt
b9LObuZ3xd00pHg2opYqw/h/EAuSnibzNLrCwVnUlVdMYkKfHsIfvRaDsjslhOeA
26ouLNl9Da7jJjAwNo4C1ZK+AexCsCB5ZAN/cw81CXmujbqbsQzBDgtbXjmex4Zp
R78j15815VZPRaoNk4Z4T4j1DRHELY0KDzU+DwjMU8avKa/+TGsRF8lmmmBuND0f
R0E7yrsKh83MJw9FdkS2DQskE/KQfOcF7jJCuY6tc9ans100H+u0arvDMAsnbqwU
RmKviotABZw5pbIO3l66bFaGLsMCqpaBWmmJM7ySkaFi+aq8KxAWVD2tT2xhvKST
60LksPUwRXHtJ6YLGNMR6vozJHMoDhBg/1sXnf1jbXPod9HkUAKdkFlih23GSQAs
IFpj8Wcpmm7s368Yc2S/VNX/rT0/+1EwQUW2A/VouBqg8aqrBwLl1vH8RVl8cHsP
BjG2ps2a6qNgooy2GLPzj6UkQrPjnWfcohdna9AHpPkpoMwMqPoFlyw0YdBjAAa+
Kl4Pk1jSz1KW0HzYEUMpxOId+H0pkP6H5kojNQ8J3WEgxixf8xlCkzn3XQG5nYVl
6sTX25tli5TQQ9w/7/KbHa8PD9PWAVbSv9RYKPVTEWmCcBzouAGJ8tbL4QXKcy4L
P20jsiejW1g5fIankHEHdVVvNxPsCtqOtoN+rrL9vsDuk/54qsHHip5572YPDzpL
SWP/9Cj0l4Qjnh30iKoRhDFifVpGywc4bj6n7Gyz1PmT/j4cGgmjGN2dlmVQZtpY
yX+ELxVJPqQ4ufrXFkHaeV+1J6f0pUkGoZYTh9NesJVjKKyIiFyQtdjkeOkTeAod
y535mNzBe8bX3rXOxoBwmT8D+ZggZfhbt8Gdl8ARtQB5lXwHAU/eKXk3hsDT3Qr8
A7u/K+z0Mv6C7Rcyb2yFYjujI1S0rI4pTpNtr5Y8pW+63G7Xbf1RVlxipUT5fJAa
veCX8Uc4Yi3h9jBazCU4DByd2UnNFKcrfSmdi31I7+qQVJeZ7KIQPepj1OyJibcu
VU6tmbm0U/YunTA8LVuFV1SZyI9mAGbqOo/7mYVtW5qpz8GFX38TZ/MJ3Lpt1y4w
l8hviOicRKYvmjP0gcXM4wto2XPybj3+/g92MZEaalzjYbnVM2CKdtymvsbJqUZG
1POMZpGUgrQePr0DYzI++KrBXc5AHYIPpBOXWU+kKcFrp4yJtkG9hb1QJY5pD4Ae
WFbjnu+RnGG13OodYqFP8vxrMMmT19OdRzrmPN+I2hitPBJujz41WTzk9zIW4jgc
cMcjVz2H6OWR77OQMnnlC5S7rtM4Ohe3myUaLXWY+iu1PqoaKD4jjtaB//5u2d+h
vKzXuKp7nNzbu4SYsev6AaqI6tVlujhja4OyTND5oFrbTZP72yyQKelsn9ac33p5
hWciRntYsLUqQHPbZvMegvCSY4Cbh8YhF7/RY3xBgUkvASRPDTiRD6iaL0U+YwDS
xJUo30IFo9XvEw7wv5c/LbMa4FOYMEVlzrpaeSx4eEfJ+Ew/LDDWhn1StzVe9I1W
2ojZ19zw7g+iAp1ONI9G+u7TFKKDyh0JFa6Ts6gm012YHvHQVLW9murvVGoUnaDL
ycdbFdnzXOMpv++PL88vDroJFCn4xo8I7ZWprrh/J5kejoFPE4j67dfXxVG//2YN
4ZEGoHUhTqdY+1vUe4iGkrKrJ5smt+Z9Aaybx9ZVR6b8fuxPGBQYBhjL5aehUiNu
fBu9geVBjG5Uy+YBWPkwjJN1Y/lvXk5F0sT9XZV0GeMV3sh2dh3sRwBNgCf7zdty
kutZQuIKXwXCA/wuXLuzrnjPnN7cN8O8xo0toTYyH9XCCDKSesgggY0AvhgWkmxI
jLNpPgCt+9RXXLvoSX/7CI3InWW1ed6Gw5VAEZHbvktKptMigYvlvhw4hoUWKCsS
L9PxcOm/Qd2oYvVoMtczO5iTCewPyExD8aqAeyjehs0CW7Vmi+NYbLPBrFM/FIee
ksJFEhrwLM2n+qwLGNpw1iAqkrCFxdwTJ44RST8ZR4s+ag2pT/q1UkpFFXSpUSZL
LryGE4UxPv2OZ78IFKDstAFDGUZwTmxDGf6TUbH+SZUnA+33tiPJJotQN2kz9RxH
lfwvoSWQIattBQkfOny/dHId7aofq49/pzGBPF+ScUb2r3rMf+RSE4C8dKDZi5FM
/dU2vlL5mt9/d76Ord+7oNUGATbyzQfBQD1pQJkuY7ySQww1Dpvhq7doi6Dy+QMe
LpdCKbZK1uMd7LhZcMztupQR33FfRW8/SOFMRLXZ+VM1dSuy8Th74b3pt8GPA4Mm
qOFc7rRnlPbkOeK6jz7oixxdJd4T1RYsev9VtMaILumvbQrEY9aXpMStIVg3lA+P
tehaQMbqFUYxjxYvAqrxRfX9mZJT+ZhBZ89d1av33zghpb5qk9Io3ngLtV4QIfh2
NpVfJdkAHyrpWIweKBvAepmjuJtqqxjTqZ9qis+x7cjbgOTn+rbVgCj/pRROah5t
hq7F0AIYPXa1RGK/UU5iNBsGQ/UewhRG0rAVP9xsY8rw6yP9YATvEGeofZt5osM5
KWO5n4Vj7I4Q5dDPA1psZalYcGXP7xFflNeUf5TjcMP+n1F6mzGDIGLjJI8Z6H6I
MO3hE1bf2iuqfg+gNbTn1Z+fVp1J319SfTXyWF3dkMKjU+xAYD/NAdr2RGRnyBTe
6MUkD5QeWA0+6z+QHlyhHhHL/n6C0aFzAW4lX6Pu2lEkliN3v+e3yf126D34TWaG
nh8oQ7OrsFQr6LB77su3UNz/DLku4a2NYADi55502ERqgGEXEZUGL8vsd6gJZlNg
c0rDEk4dMLzYP+DUwOy2YbP3c86/pCUdRMVV4/99zvAJKaEncsItPM9bdiBtx+hQ
rOe/j2yyiXfdZOQI1UABaRliXEQk6BWniNo56v94uI+R4VRijqFu5jw9c1xpo0Uj
3YInohlj8z3wzORQDh8x0i4SOent2K3erlAW2ncOugN/zhdXPqtrn+stqscyYx07
OsbSG+s+PFtA8MdxfC9lTCWsdLkSB4/EyE45DtcLjgHoG9RqU2KMm388+LnrWJBa
buPwj7cNgqMe/0takmPMloXe453blGtQum0GY3PRpghKWy+KSM1GRVuY1PWJkhj6
9q8+Ode7Qm4sADYV1TEP7uygqub/rVdbrhoFowcwnmTHAOTaId33WIpe7hcFAXUX
lbilpuJRNYKBTnoiAHkaArZZ1btiH36/RDYEkY5PFWsIDYGT/uN7ffbociK4d6eE
84qlOJWvp0oSKMsHlBiAe+NvINl5TwEKE85u5GkvKXpofJ0qFgRlNp7a/apJZxcI
3i/Ooe0QZxG0NCKBzmBcnLub3gX1pTKvDRnZtww5Ym5CbrN6FkkfGStVfRIsPwS7
u/dqRCxBn0oz9QJ9b5kJ/PWoHzo7oov8yWCvpW3qzpR2+05laDFk27yL/o9bymmw
ajrpIDZNQPG/3thLurlQOb1e58pRXcaUMO/2jQLmXxERfcYOuIZnHRCfziUvyu7q
a+/ZjZ2cfpF5Qphu3JDE/Q9F7pbujLd1s2e4gVJwShXew5ySwkRWmoKY1lvDG34n
zcQ1lE/iUUJalJDA3jYLK35rnbwi6ECiUQNutW7CVKj9JNkn8iJzHilWW1cX7Kra
5FC70O3uuAbgcmSnvvTrhMgmkpOMq5q4rOm0tMk+Tce8r6SvzmeqQja+nrqZ5//f
pG3bp2sqb4nTwPgL+j8c34mPlPc/OV4ehTgpSgPfdB5nXiRvzorI1vDUtIXoLDKl
M1ui0DGp6boBZrCS+krG7Q68C84kTqUXZHvWviNV1tGlAXyrOfot+WWcmC0Ky6PB
duQfoEpQnVJX+L/wgJwI+IofRhmWL1HyAhPGpPsukB5Vfh/z8x0Yg2i7ztHjLh7j
7Qd/zvUO/FMd+nDpBFodLsdsq2K0XjE+2s4M/w2MgtaYD9GnAmISsWTFbNnPI8WA
t0BYRlZVeMz7qFt1/ilCRLRch1GXKj5OGlELfDkTJxdn/NnJf1TzBtCW5IZDj/c9
fFwFe9Q7vJYgGe55/gZ4o1BSUFlPqNt7H656sPQd8Gx+N6L4DIiDMYaGh+GrPH2k
sRGRvbeQQKN6sx1JuJvhMB1RMlqsd+qffzkuE8V0ZcQSUMe06LtK7pem8OBqcsNB
qZKV/vdcYvZTRifFzjWYDaD+dL09GT1kYtPozJx/p2Ma75GU8KxJvcq8ijZnNFLr
UwK06PnV+3MN906VJ69bjvbL5nh7WmPuxvK55N/5fsqchcYJ92f8uf1Pqx32eL5/
LqTjmWyyUv3X5CJoG/3pih5eDbKrexBIgo2avrXKy8kcmqUh/8X0v1cm30phQ+A/
Th0Cd7Ds4PRXKNTtjilpEWbZtz07rE2xdzBOT4vxPiHORm+8pvXJRwhvzv2Lg6sd
CvGRoAsyY0nKePETMvebkH3AXul38eU8wOIE7Fvdt+RCLGCz+H2vOLjvg40J3zwF
fCQ74fsg2iaqTr/b/9NkpgkCwJ2Ubx/sC2gLB1vc/vpFVUOoS1rnBfjWlPX1GLhJ
YdTV4Ta0i8UANPSm0mRoNn5FSfyJykRG/dcgo+NxXu3rlpeHkq+otPoTmEZN6/aE
g6JcagCPgMEtPqZ9Ui0vB5i0/jOmgyy8IU27Bzbj0GVmJyzBqdm4pUKqG81teN65
eXAGxvkJ2Z2M0WFEq2rXZixU2z1hfdnWkNt8EQIGkfgLmet/j71Fw7AIG6lfzL32
BixVUzVl6Z0XLoVG/JgEGRwAPz9kyMbjFu2i3oWVQkwnRQz528Kjrr+XE+obdE26
ySrny1VXQc+Q8muPEXTma89ds5zf0OAc7urkrpC00Xdj52XSGjlEZ0vL/GvMnw2g
3LJ8xqqmFX7CLVmcCO4jqW4H8e4zUO4Bngb1PzJbZMnQSt47fddFPbWBdXi1MhOX
pQjqZrMAtKSBh7g/FMHPjLSisIsJb5W8XMVNhFSffJjY41Afx5VRIY/A/hrScXVb
xey4il63vZgXcB8lSz4GBubLkkhbR88wTbEC6pJzYu3FrB+/+zi5QyRanAB8J0GP
9UooaOB9IRub7zK2Jkl6HQ3PisBZcH4tkY09zBA1ZTq699SLD4kgiD9HwXXLYI2L
UI+bD7AMSf/DZBq0EowsUMhT4cAGf8AFVno5C4bIwCevjNk0G2Bw+5wb2DY3CGqH
pUQfYUrxshoY9aKtYblz/H8m3GMSxDAu8yZpwPTsk+nRsXoWMZiT1fMFYnbWwOFu
yqd8aQdtaY+XTgwSF+ou7BjI39zHNYLUQ8vWRUE6QczFdSdwuMz9pQfjL5A6lK/Y
SSqwyMZA/lNMkBGKCdyiwWpomEy1255CcNxiANVbnBNvyrRYBmX6oVWM7Jp5vsGJ
M3cbPd3kQTIWj2pQlGuMVzd9Vq20dZk3/w78CdjGkQwHaxj7iHdg8E/uKicaAnAM
5SyVohqjRuUErrQMbWBwQa2N2XFqKKnxsi/VgvGaKAyTdrordfb7D4+fwmUdeUUv
IZJdtlAKzZ9Hmc5E+n/zI3h/wrNo1cJP43zfcSDp7HaRNvEO5rxjif7rK7kgM5Rd
/AeTv2hoOTbU/h4txpkV7g8aTp99TFIz6N1iAoQr/b4C8oRcGFRj8C6hV+jK6JUt
iJN4Qsx7t9uQeMOPduuDJeMuZCvg2dUiAhh+Qg2ez5uFwKXxS9uOqPREn17I4rce
g5Vdt4BvZqWROGMd27be9yJ8HNJq95revidVGsy+NkUrW+U+xe+0/gytR+EqUHD9
5rMZ7LQfZAVbj3mqNfAkBB7DAq/bqSob0mTOVsTPx4rxvGnBQzZ3v/YaMw9mwOe9
MZN0lHMgoj/HERAZaBrtXuHLLYOJ1B40xqQx6g9k5nFQ4FBzrfepij/f5sIgkZGw
j/ZsFbEQDlsTFa24dWDP7xTBwFsSEMCDO/W/AdVmclnI2G9X13hh8zXjziWBHJIg
A0Prm0USjrEO5xMIBPRwL7xCOlNAgQp8mzexpldpG4ti+q36kzKaf7P41VqhqVcj
LoYyObDX4t4XFDzuuPusMbWZHA+IrWSH7xGTKv+ZLO3qQH6ihp4IHPXCVeejqiZG
R+6i5N1h/cuwswuZzWDj9cImH5pCymk2Dzxy9aXt4dv5TOFw2rmTQVzmh9NmBz0o
quyj8qoQekh0HLEIPnn37QDZ2IHEyueg6HRK8Kzym9WLb1/UnvuaL0QJ47K0YJkc
oYU0efrVGFKXiGnYkYlWBu6HGaJSmdfSuAhk1VYCLTvCTmbToOQhcWybpg0N+H+C
DbMG1+T4yOjSywD/yWNKs7UhBw14adeqC4vae2wZaxx7+1/AlTlLJIzn6dF/KI9F
8Rk4tiTFlnZDo7vvPsFGMdTJ0EyMMawSj9GuG3HZcft2nx+KjbOSs32Ev2aSZl5s
7Cm0EPe3LcKvfzqOqAkBeUgOBe9Fjd8uvMcSzVBKcvO7gS+YdOuaNcorc8/Qpe2N
f8xA5XrkDRevgMQHZlhEiMfGomoKMcRTQTQt9Tn/onJoxOC7zHD46NBYxlL8n8FT
dAfHEVNmwxbz1tAGeUVjeFWcCnMo9cA0xIZn3ZFdSxPa8HAqHrGLEsIBYpVsCUbB
jG6k/5iCjDmI1wMpBe/ZrFiFUlt4wwjbvV0b6/sm/CJ483ax9NDcDx99APSFiboK
r8oCPaFjEgdBg1QOiVn2c3ZyPfxp5M9mHJAJaCxwatMRTA0oDcH5eJhbLNGF3u1t
DBQSgxXAvi4kBB5PAOXnr/1v1jBxMD7r2H7jC3cuhOk1YhCMpkAI9KjKIslDuo0I
iqJWlVTiaD4H1Ri1/sBlse8J+NX/VQ/mEFfBA3FjyfQZ9p9oA5gSjUPATbO0Z4uS
eqxjdn2U/Doo4XLVb6x0BY6hi0NpgmgGYhrUbmWZ6EQklqvx1h/MzD0NeA8CwJnR
3ddMxpcSW7/SOzwM+rIMhPN/blvt3PeVuF5Q8sOoH2zGVWzCMqLgH9l/X5Hl5SHt
i+KT2IRF+Sq+zEK96ml+ncV1Kq6QAfZp6+BVuXJr13xSZvWzTQ7f+Lm4qzmaHOZH
dzWg/pW+GhcqT54jdu97R9XIzlBwARKHBB6CmqGALw9hOAuSeS3B2h7pxmXC67S8
OD4tzunrrUxDgZAwOG9YDb/KHOR5iNTVIHnLxpekuZp7+uTWtFApX/JQ9vzg7xNE
UZUxb/Boytzbmp4PCXwhMTjLwFQwgUFCwsJFY5Sj2duN8bnEnphybPPWmaA4dje1
gRwTubtygxurWQ2IQQAkBZyqAfEijohBO/D886XGRSfx2h6QkGmOFI4QdXBm0dKx
HHDTDPyPyrGJiYHgJhRiXbpkW0gdLigwhEEqk9Dv9em8t9d5onCFjK8DnInZhT2V
eTfNM9Zp8k+E+Wn7AC7d3ROKehKONulEhbQVz5vL3PhZUek79NnAvfaPj+fONfKC
HhMGll6KluircemLQJ7POq4ryQnB9lR0k2MEcAe2DH1A0ib1cSxt+xwt6+O/t46e
WXQ/ajYcc16vqJkvfiy7pLHxFX6yQ46SCcW3OFr+cN8UP4Vqj84qGrpDtcj/9+0u
5RhU1MusfRRTW+UFOBnLaztc4yrgq9wqxMgLYRX7yEam6Ah4TPpxBtvpzNKop3r4
9FMXmiKFS3WBPeFGYKufS84OwJMqs7y3Uw0WIAhUklAA0Zk0IJxVNZx73zY0Dx//
Q5CmZpM6oI+nCuWvAtD1iQWLZfDGz0+duLQvj+MKFAL5FMZSn5N/0tCBpN6eY7L4
a42knwsHgkZBkQmd1h+6FOK0FY7ReshzhI+fCu0l9QoUZCtgQ+7MDJzY5CskFf7z
pm1+DVLsr5V4oZ4VIhQPnEneVxnWPDJHL+TBeEpHVWLI9oOfBRF85VWS7K7XM4TA
58HQ7S3R8Rva6Uwb/kgkf+TIGio3LNylS0XqHmfY4wHiGMbg+eOHPfHb5SzVApft
914JyfFJ0KkJmOz+i8xqwvu3LfsiArEh0h8dTUp1Usg42WNGIlReTiiU39iMI9oE
PemDbcrRGYtd5WU95U2lVobqDIRAiwL5mpLj9FL6tTEH76+JqLeh4G4sOlueS+J2
FqLDrZ/0cHX0Z8y3RAa6hMOC+lukrpoZTJ54yO9HaqyyfYbwlRq3Ls6gXKvNPkcs
fDOSLOZE/NXrZuqINaZl08Ol/GgrgLInIT3V1MRJxSIwq/TJJDZFTRRrtqSOuPyl
T3HdIwNQgbKFiRBSKKdWQQBdt/GXbrFdLqRBQFfxZjKWLUcaozITBtrazLmZMQmQ
WXf4yA7YgWcLYHpsUnx4Sccg99OcG6S8Xe1PWipYKVKBoq0y3kfYdfapVs/Qh6tz
W2NcKwGf/DA0nOnv0yLcxtD59tSwzjbM6Pid+te8F8mOGLSj343u6nbzC5tbb6AH
aLGhUn08P608s/qXaNjvA3LxxyBKbvkbM/6DR7ujlxDY7ctQ96mqG1bZC8hhAyIB
St0HaeY+0nfzXsUVhuLXtHzPE8OOPMf6LVeE3SR1sYp5kLfdO1yZW1bd5JXv4RVa
Pr45SnRpRF1Jj3jhbPtdmcz0tWn8oq+jzL3+Rl2PZ08G/LtYVqxx+Ki1iy+xdMvV
yWDfUdJ95KJVqaPGDXW7EDldpNt4IuAc6TX7KpQo5H+3UowX85hWRd7NyaBArz4B
Gn1oamC6qdxekSTY2rpH1eWVZXTEeghrb2ao7jGyRPVrctBqhpxanQct2ZN4l9e3
y26zbApxlmMBYz3lXjJUSi9Kvdp1D308a5lxm6vTQbghlGnmGuao2ArcDbNL+TLI
vG2dRbGyKjOy+jiwaBNP8c1CaVKCALQrSagrI1gfNFvXOLvoYw780V7s1k9q+779
jjZYEkhJqxb+zIAHXv2gkup1yZ3+ZWK/JAUtpKvO3VGzHMjTyiG6KrhiIJmH7ps5
laGaOycpBkCV9p8xZ4u/lSIyr2vDcMAofU+IjJLB1J8z/E44iU+spvAMeDkjJOy3
G32dzXoPdNB7pr2OA3VhqrcfF8eBuw5KmOWqK7r3LfF5639yVWvS5yY9QTUGRG7v
i8vCRfRCDUbeyeURCaBUro+SHXK7AxvpotED71yViaYx3a8MsR8ngrPr5bl5hJs/
r21V46a+Xh1tUt+0Pdd7QESa+fQ0FaPI74+PGAkXkVQ1CSa/Eenz476yDnfyV6p3
eDB9iOyqAhAzHupfUu2Ltcg3BTCt+11K1q9238n8FAACu72S0mfIB6ibIk8AoyVS
G4cAlCgcd7ttt/sqPpPURi2dl7rTdku0o72odxaNhwon+CD5Ii/+jmz94vwMUXcC
vqKQ97o1mJPE1cQ0p3ZeRRVdXUrzuDPaq6E5bnfCShGM8LnIJKdcubU4cC2hnq0m
HQWLl7AtMwtp01u1ruZnWQ4MSj+5E2uzgmBU6FTdgw4PHpb0Nx+66/g4GkNEP/H/
qUEJxWwhMfBu/ddsc12d5eGkfSYLjMMZFRJl2Z/6G4UiLThZKx6IgtHf+jzGQpA5
WF0y5b0wZH6RkbZbVrKbKI/4/XMX6dhicqKxtGzhUnFRCYojOC/e8bZlrBv+hESU
atxlyOvgnFQZw7mvM18hRuPYeP4X20wG+eOcsl1H4hGBPPNaJwNTPdCSSYBVR+t2
5lR3t3sZupq3jYh3xBUccv71H2Xafw83RknQOqfRxtAEIf4AHnmLLbdhXAXxrM0M
Xnk8HMBS3nhaNx/fkGBwX3Fztp7jUoTwkSAzbECa7b9VyjvFbRq+nG9Fy9gM6Zc9
0Mc+w9F2exD8Wqor/Ue5QZjylFb4r1ANF53BZ8mN+SOXByDJlWb9B71zPaPl5b5C
Ymrd4PgWrsySFT4stBpRf/srUT0RlAr01LgyTdAN70JWqTAUKpgde8HHM/zRqxgq
4sJDOOOgpxJmLsWBvjxSUtqs+R11tmS/TbDRFSKG7uN3YoIpLb+T50aagM1rEjQm
zITOKKy4NBtNHjWLA2c/JxuNecSZ2NdAkOsdLuiLLVq8WD04OvQpPs7crTD0i4mT
ou9pOwIUg/F8sse7nTeedyg1Afxf2Y58pkt5uKDsCRASxyaX1xFv0nP5zok0IvFh
nyx9nkJomUbSB9JXXc4FQfJvqsmLM7sPhkts6aeTj4Ta65a+N2CekwAAGFOTaekA
lNqHkQrUiZkcNxm2ct2Eq/M6XyN7THpCP6C2DuqFoSWoff7A62skFD1ttLYLGabD
ziQVXu+ZQAie3qByjbZjv6ajFebMxBOOHrGGIpSd58hMIFzCWLxLMPZ1rdM5EVpg
vHZPi63aFV0Tu7D/fllacJWRDPMRqDFY7bZcVVSckjZdgY9DuMUXEnYw9o7xlOiU
ToN2JWvQLp+lfJFZHdgGt63gEsHtdGkhr/Hy7xHpp9dvcSRHZfiXILctK7e+kocY
hoElvVL763JfODDfTP+HPHUnXnmiUQNPNH2ryQoWVKp+L13bmu4mibvPCkVbeT4S
qahTNKA7C1Bz7lj7RlpdJsPM3Q6jmskYgVJtkHVgfgN5R1cvur/jtMlf4LHXkZfd
1eviHWwfA4EVjBLLG1mlUTXT8E1tjop7lWyrGpixRAK1rfcTqKdOvWi9KjqPByxc
Wsj4wk8qnjVuK1ZCuAt+bUPWIy812aH7CvWIaN8Dxgls+eqBvUjntdJh+jzQkpvU
dcOpP8wFnv6m/jszVoXmaCqVHHKePYCCxBuFneixjgzuuLTbkZD0YBkpIgDQhf3Y
hIANYuHFUckLAl39CFot3Kf/PaA7z7Xb1rIG7R61wG6L1wLtgF9B035NHx3iFmoR
IyiA9vQyocK/ms6VipCaG52jN//qRo2tE4aVbvZFQQ2DVH8VTmLze6KyGbwGEu0K
+q2UR/aTKtV7zem0U+2vHZm5lOqL2ZMKJ3/VIXSrh9w2DIBjoq66p498TMHwrArk
K0nxEOEYblWxDluxCOnzbYleVAib0Isa/Cw41Iv+45vMe+cjgHH4emoalAlOTyfe
l22O0+KCJeeWlBf6REy1gma1o0yW4uz+mabDJI+6ArcrlFDMbFMPYizMEsRPmmHj
c+AvO5RekuLbdBUb3KxlRtpiUA8Z4hW8vW17UXRzzBBWLFwcymQJlDI+UD8z0uWv
f9OGAei5jZzkL9yE3qKSgE5JDCiVRu/o/vX7wr9nL0RJ1CkBHXu5bqEdWLhN+69C
BbnmPBFYeofNsF0tYjaFssgZjGxXqqt+80USv5Cu/qg/vrE8Av4C7imYxuEdd3Lh
4h4JZcsJWPClkMq7F8XsFmckje/JitQGVqQgb/Bt+52RcV3gzDxAw8eIr5MYbs1G
ge2uq19MF6S3sZKtUSwinobogdUpb47wfp0AwzpeGFpghRCqCkBASMvfII5EFgkB
CFxBbEJ+R9/jNPd1sFA+x3WlVvRZ96+t/evS9Izj4t00sN8Wd4Z7h76RD+OCiRXN
sbT+Y4mLmvRvzL2GKquLq4M/qpPGcDasKFgZfODvjX0I/90SJq/bJy12e89A6Hb0
PKBP9A0wd9123+K3wiSfa5lhHjhqiRPr3UzaoaUobQBAz2ZxxZvlkBOLMMYz9/Vv
kkayh19IIkSUj7/Aeimu55Y7JPRIgX2xs0/yVF9HwvBt+e50IacvTdHdlBh8+E4/
BiouITbtD9LFKIV9fWv34/Th5Av40hfSm6anySxRQicJVvZJ4iV/bfUnJHORa/Yi
wU4KEk91tw6pgLXUh3cyC5Qk4xnQP9zbcITJnDO0R2u/WAKQzvQlt1/WnfvSR8WR
6PJDRXxVhCIqRQVC9eCaW0AZtxJfkQD3rHdKTngtS7C5Np0QF45SHeyzXcAe9x6I
487BWRpXCjjBx9XN4i0UvX/UkvOJ4hJiWc109RK3h6ZA/AOJq1Yw5GKabwGZtNeS
37XCQcXz0fTWWP7PU3Yj7sCL8CjMx3vKI99E9vFnLMmH0TxZa+wivBypqNJcQsC8
cYZART/u0JqaOtXzNJsZsbSLkVhGEKDPrztpH4znwePuHgesL1V+2Yy8drOJ7/+2
Ds/YdbILapEHB5I8pjuG/SoH6P/eh+fPD9T9VBF6E2OpMf/37LxOSrlwRwlBJuT9
jnqkPxrn06oRFsBnFltbFgbjURrBTRH2Wfad/GzC4o7iB5QSNEc5dLlsapqWnEQT
F4+JFTpwAU3H7v+Le3HqRz4+AVTV06SUOxwb2S2DKSGORByWfRT5piSPVwPN2Vns
6ztVKMs5w6NN31XHg5qprAcdxVVrHAYMu9FdTeevJ6sAg8BbuF2MgYaRSyQMJZm8
yLL2g3aH6Y7elxLQcoqDVvlhQn7k/Xe5Fmvjqtn+DRxMhn8/619eLtuOPOxTG+My
ST5AgKF2JAf983vZm/qczJrKL2P9YyhoIzPTtD0w/6zQyugRg78pZiD7EUGkQfEy
ulkR514KVRv7rTpAh5mqKgEceMHjuWKE02Oyn04jzNlvdzbWuaBWopFT5DxCKgT0
EeY7t9epTqKZ1b1xvh1n+6zUfxJmFWkv/7eiVuJUfU7TSS3Z7qg3Y8lYzovDcNsV
Xa33F6pYorwTyHeSPU2Zt1c7Vfb2coGpGrPQc6JeRcozK1m5EniHM4lv1WnlW0ex
IrOwg6rIO6xAiC9Fjbv5D77Qu18uvxvTjv+jVt/JCVGUNfY7iPimk2QYOXTnCYJh
qQj/aEqOFFXc38I9MN6r60cjcYcZmrlV6HcNHLjmXox2aaFDQol5VWEt/P0yQxfD
/VMiNwoEVy8GkUG7Iw0gb6yhXb9tpc/CgnD6fpwqpXh123/mJPPSRodt8vRhC614
IdZ8ZjBOJd1GDM4sZ1zLdqGbS2dZUcEZxvmEY2HFlFZvkADAG2uJsKgWhbk2Mwng
4S/464cm2a0H0ImG5VgCYI8y77x+0g15CIfjhQkwE5NZUgEXY4gGP8C6QnMxLWfK
1I1V8zJTdWYUuDsm/awJpUeGVC0j/YbI5hJ2/svqRmZNxpO5uOpcU86xaOc+gJa6
2vieoAQrnqNS20dnF0YnMl1KqpHv9HvHPkDmzM6w3cwhwwOBNnflm9dUSX5+PvYr
XDc0YewdtqQp7iJDvCRh57ADrO3QiNYRHU8g3spWPn7yPgLHbClsYGY3M1UfHGyk
ER5FOkfDnKdcL3X7V1HLJvajnIL9omDmRxB+QzvRj6IPoemShOq6EfsLPgT2sFMP
NVNP+rC3fzexlrLsANSY9wW3SBUgKxC0VEcRmwreVWRvuxHV8Uw51IAqGAIfYjEb
snrRK1PfaPPUD7/aep2TjoIPFOzFnBK92W5K5ltK48lPfIjCxy7kMr+BNrtdmpOu
On6pmIC3VtYJrWysYDtee2wZLmc6uQlw97VhZ1Cogd4e/uN4w69GOsLmTL8uf27z
lIVAlkiwQKLqVdj2OS/ptmum2xfd4Pm5M5r151prz6aNJ9uB5JT3MxkGOPPdYVFW
lqxnQtomKUnJhrmo+ca0MJzf0PKJygk8H1KN3Tfz0uiSRdaheMwjOgK76HmCpGly
WioxBIHWJFIwL9HuBHMjpSlZJ78Kpmg4GB3r+/EeLQWrN/sq1k9ZT4xgv5v6tDL3
w65HHJDAhJCJm1WUMOf7c4ecfetfoaF3GiKcIXZZvNRBThM/n81luKRNlbRJ1Ajr
nu8eDpeLR2VOAcul7ckX8iNmBwE5B1h0tnO8XuV3Du0RweqKl9SpyAdbX6eQja1z
HzmMDmr+y8N/xvu7trne802NYN+exZQVO51SfbmTI88ZwfrVkPayYyBFG+Rv3SN4
SGX0N6VuaqnNT2J3+J0SShYjO16qfB6SnNQqRLXkAKJFU+f+bRrVoGaRq3Ak+zr9
72TdOdHKWe3vfkw07Sax1KH/p2SU5+Pzo/HfgtnoFCvwPH2yumXUPlQqRhqsuMIS
OChwK2iuakOwnbxDVm/v/zmOz0wEvgukUpt4jBIPXu1Su0zzyPFoC+w2rDWTTjsh
rEdNS+3+28myAisbXYVzw1DdF62PK3esPmEWtVkPZl2fZZx3rPfRzrEEG9ZFRA7Q
8KJvzSqFkLEl88ozgPAej/z97/s6Sr2WYQ8WUlNaNSohP4EdmBSkt+sy77cBycUl
3Gvji56kViPyw0JyUd0q1fPGQcr0nqZao0csqDczEvZ5dHL+DZ8uQkzEazdrHwx9
iQxNQ2+wyMAARgf+BfjBOqJn0N+G+Nn+DXT4+XwSwfxikjjZ1NN1BN9LUsn82ED2
kkjB/SYI002gZ+uR94RFlBkCl19q0V3+vMKoPXOpOE7omQBNKODOw9ZFeJByWogm
ntePnXxXjTUfCKOcrgVVRVYedyrZCvMl+ovqn+QXka+PE8XnTwMiqhFniM+y9L4T
bdoXsKlhGjevGtGCvqay5P0cR/UXRWfpij0Ua6VMGWcKX6uMJDlsxR41tRLyOC0H
sU73oPUuvUahaWX8a0nei83bTYDjrh4mKpxUmS4+g2vNBo/WNr8cBSYNHyJTlI+6
qgmJp44BGG+kWzRkvYl520ejaHE44ZU44NVdQMxXMLprMeQbd8mcBFdG9HdcykML
eL3LFW03w7omO/sVjInDtDAcoEEs88p9MnyvrI7i7a95ckYfPEDaHJtldx/tqOo6
WYc7/CGlovCHaBUNePv3+FrKPEFIXiY6wA1ZR9aesOaHNFZjCG6H1iyR54yncRhV
L9Yu/LXKDXNrwjaAF/aQMtHbwWKioUNtx8BdgxAr9+hv6QKBuZ7/wjMjG3swZRuh
Xmd3nfIivU+u62YPF5AyiRDFfG7PNnE8vFUbTE7op7qbPar0xd6VQlTQpPgw+63B
ecUSMfT8J1WAsUk7ejlQdKetmTnJSw4bxPiiLdVIMQOXjIGmz5kWCC9JUDS2LgSE
lbZE9eh184/iZnVuGBAfk0R2uy3dCDSnL8Gw7qrJx/9RwwIDcFcFzffS0cLG4nPw
IM9po6r1HvtwSAA3GT5+c/hSy+SGc7C5ylPJ45kUHUE7MAkbV/WQOBYu9fQU7UIY
p5FCvZViNDQ6cJRi5lo6gHZ1dOtPLUDwBT42smF+u1nPU0wTfifo2ycqUGlSJXf3
+PdHJ4jDv9QmQJ7rTfWb4BqaRFOCUo0pbfNp8vLz75NOE5a6HYJ+cJggVvSC6Ybf
F3p5iCasG+zdbszgLntyrkItNdaM5oUh5Vbf2YUqLYbiqP3Jb0OAG+2//0heWgWn
swJEaG71ekHFB5QauX1Z/tdXsJFZ5f8oDt55Y9xoVo0ke4R8Wa9ZmVSD5rK6GXhh
dPDs3cz3ArxLknpR9K9r/Lpf6HeaOK8SIl0Y0VogGZglVLP8lCeiQxBBZvonJzfU
p/hqoeInCm7yl0S3ChHm1yp9sycAKw2ZOYEPrzpq3KfHSbctJcBD3J0JBfU9+e6v
1BBKtvUIsuMQ8mqXYLCKEC7Z7QeNSWnpHdk//dDTaSnhPWjJqE57X4W91DkOtguW
EskLhaxS1nAD53bX3LRPE5L2n2+XwYVCstalWDr2SjHb8ivX9NfaXdGMlmWFUCn8
FlklTbLYA+LoSS1eOFW72f4Ck0cUJ300Ijef0hOrThGsqOEhB6AoGooin/vNSh8L
Dx6VnOQUhyrcBfh3YEzMMx7VpGsqG9Xov9gQEVSZ+GTjHLwc4wqcL3pQW92+8r8S
nFsxt/aep1tqBOhLwu7jLpN/RNx6tbbJsGRUIsVtizyJQm06X7SzmG6ZHblYZSKE
tYQOQTVk3vIf9tu04VVsGLWYExjYSMvgQpmpvkBwV5PEJFbouKpyPyMmaa+Ji8py
NWONm3ckbgTs/90sJ95tFWDGAiAuW38ta5fwuuH3r/ws82/brs7xPhXW1bPq9z3v
GpfDUZg7gY8nhv0F0OC+/knpoyPKtOC4lzuQ9wAOiclu9WtrnUfei3B8UdT2PArp
MrsLo0IiD/f9g9ZX3pBj7aXWrFh3lbs0cLur7cDP3e5y7FsnU2QNccyO462FfnZT
u8e3tf4cESlt1g/7EfIqXisXrsqNE5W7pxCLheo8puR0ApfkyIhsE7p+YYDPvplh
9V0z+QE9Z3fWqnRpRtN+aMlqI7MQzhGbWSdEwAKUeZhfDJdyfQoPeS7krFBba8RA
F0dzUBV5KBvukvgzs0kG/oR9K33KXNdNQjbedMosTOxdUkM0aLYtpDB15Aj2wxFV
ljnQBrV08SHrqOt69Bsrf0OLRKAB6cd2tQQtlJl6oSQ55E9h9xnl49SjKDlLvPyB
sqNwDXKtqFV0xYGd8b/7N2ISJxN4IgZ+OU7Q7c4vgmWncx8R2qhZ4eBIpV5NOUZd
/ceUihB8Eod5N7akC1W4vPhInbGfKpXmW0EC269z3618LwhHOEWVBwJfV0EsSWmD
AOJ2242u8ub20v1SMBQr8KTBagiq1MEnM9YywMHa+wBCXIMoeTnzFVLSdUXOnRys
BbYHktLagn0vcrfZY6ft9TcZJN+VCYDoRfzuR9+fSZ8/6YMtzAPP07Wb9lzPp9h3
Y1MDmGUCjygbNBwVTS8WlEQPCFCYtAE7WcozME4+i1jkRTPzrAD17wRmKySDenTG
GCvf5sJYH9NrmBklkHe8U4RHeVl7PjY43du5T/uG9eWB0jzZG+/6JYagH2VVBi/i
O68Ie4RXzoU5ENA2tH2fTlwqeBRKnH7nAQPPuNWhS0+fldMAf7Mcn3pus+LzU8z5
plK5hDqKpk1OYyk8ZgEzuRzeJGmP1r7U9r/jjKrx7mATkz9TjNGb743GeHf1jpVv
miRlWPq8NZAGsbYXzYO3BYhZXNEV15tVdzlwb2UMgkOVEHPoig4HAomz3ZPk3czQ
uWWyUalMt/jgTF1TR6RWMtyoJUamUq9+H686G5kOYYguUfSxnjZ1IhcGykXsL09T
r9ve4H1US6xxXhMvE/qNC6zVnwwTbMi+vSpDosZRtZScWi5ETZ3C/3v2i1NVHUYi
G/mPVeh5ZfpQsv8Pe6BAzPSKdOH90dc1lgS/QxUnHJWbIgjDKmPMNKBXoTUzClG1
MtPVeCZKSGELD3f0n2wNKoKMJmkaK7Zpd4mTgKqq7/y6OQI8NFWg9oZXaSttcQGC
d/CsVemD8toHlH/lLVVDzT35JpIwkRnXM8mMXSZx7YpZB3+vmEpO7sDt12MY0tqo
c0yxbGzxRyFSBhsLlBwS7W6cUnPHeUGqyZYaLUfjfCa8t4vfVtshBepEg3hGqX9D
bYX7T+dv9txV6n3fx3uRdNALaW8EGbPDA0GN0X8XjvumAcF0bAMngt5Pjv7nqjHt
UfL5n0wFiYQDlAm7OVLgyas8+RW6f/FO/N0qVm47atkkbKpnl9cCmGnzx5wLIyOx
9DqeKFD5n6QBzKBsKmK9eO9bR/dvfC2XlmMd+jqn0kYvXwhJnfoy00Ye9kN+bREu
JWXp6VmUagNjPsRMbSZ04/ZQ7hVsMLxCadsBc+W6/pJJPR6wc6aWYV4Rj9lddRi+
IewGb0gUkWgoyk54TVx9O4cbrQCtnOf/yFYo+8TxPVn6xpeKVQi5ykpZBQY63qzx
eP2Y27af3oNLni05yj2bW7umu8kYrJc09lWYt0aYkq71/TOhR2AwL2WG+pKHJGgU
S1wDm4go5DCvq2LGXG1EoGQRnJZXSerVnxDbBcKM0AKCRREg1mgzvRzHHnWMCB5A
mBSpWnz7NZrxdTs04zyeIN0yJNyTOTM6v7mx3qFaWs5lN9r6rRomYw3SEXxb65zP
zj4aiJArGVN4ighrSroSYS0WDk++OaG33ACFsMzCi8BgOkw0QF+3KUbix+LooiZk
K83ztYhT2M9su2vS9LqUHQBIc9/l6W/6D7JuyH/VttZ4k6j1qMu7jkXcOdEnHQ0K
fDkYWgGefyQjSgoA5xlBg2H+0Lyw/vPA5i5nFVsL1wOUNvk1QgxLBH7J+wLBnw0F
AQjemTtnEvj1bTgyRYUhI3DvGRGicxMN+e0a4aTHa/oegNstqZ5TaWrEbz5VncBm
KBlM1NFUUzc+f0QFVAdAVg5t/mH9W3aLhxiopHtbgWlUCaU4VA4AlOrpEXosJ2Sy
t2Kgnoedt4OQYl5YjKvodNefca51TGcUjbxp1lbFPzr0uvebodI9XczwpvQpW8bh
4zNQ2EXXnG2rtsYAViY2ArHNlJfdRBj/EUfVr5ajluJo6xVNcDfEAD69cpipnXMA
lW9llVhLDbLCh/p5Ce8cAHm80HchcKvt+gIw6AhK8Z05jRQcRapCC7f4MGb8OzGv
Z2xk0RZqlOgdCJbmHjCnXC5NaRTMK+1FV21OlEsOdNhuqq3g6i3/3U8scEnLZtml
m/pqzfZJ8j2xoM8d1H0IoGthyNuLfqeYhrx9grIwB2DgBX71LS8njL9c540hIlN/
L6IZk0d4lDYhLyCRlS4ceXO1MXeZr/pIQW2V7FaxSsaQaX4HqSn0Puk/p2XbYxe6
LJGFKtAHnTZP25gLOyIJ8pOG/Rzef7c6siza6f+aQ7eUTm+6KLvnFl1PWxRDAR3h
JSisAE/fN8mX2QX3IyHRXvbFv9Jg1ltR5SBhdVsjUoVANZwKhJ0Z5leeEeu1sDO/
3RzgGdfUf5XstMEN6OYhPA6Br/hlBI20YppcN1ii/CoVhgm41by2ie/0cDSn3PqW
M41JZjEhWWp5W1XNzIIUG7ziC3j1vxDqISuXnuP7O9oHNy/U/v4T5gTTZvD4iZJN
5frcul+sXKofyc/DkRmBRDaRP4UfYqxFp65g2UwWdlpyd7oPXw27+viPQ0CV/OQu
QIBz9T8LCChAUX/luO0lURRJ+OY9ptFPrKPLi0/1ZgJGuQRhsXZ9t1bckj+KFfiY
lZIFYO+kKT7DWUITkrEGTW/A7G/OmLH5/Q9WbGqfbXrSaEbXmliFCWGCH7VNnhgk
fvB/q4vemuJUm9F2Bhtmmdcho2PEI26dTXh2Kr0LhUN3VypNzlMB2leuWWaj1fs2
86GY7QV8aqWv7xmBIXM7ov21YO9ywYcSlgftC6A3ANxlV6wqwHrzzWYstDJkjAzj
pMi09oYQz9dxJygdbD3Bk+6vnn7lqL8923mGS3SxorLCDuK5LtJ1YKx+5sODO34R
bDyJB17AKqHWGSvbeDv+7lhmsmEDi6IfQVZuAJBARJfNDw13OwEAcEMKTQVBokcl
esbgyDaX5fnCLSCiRS5fFsiA8CgTB7zmQumFspALD0Q6bP69VY83hr21+0ZEiwj+
xQjxZ8EAWcXhQ3Nbj8OGikZ7gyUsk7O4teer8zLgsukniKSN7ibHgjlAmfH8Wcfy
PPyvMqb3TDpxKV0bmtBlpISI0sYzXzbdPPrAhZY/Fbfc7EsZgbNWqEzLiAkb+wD+
QB1yBGXdzg1TrpgMOdebFOiQDyhBBwLyQqntj24Km2X9YrDteucOxM84Ho8chaEy
V0q4qgTCBmoG/BTtfg/A4MmH0iYrVrxXk0Oxb7dp3gNEJJEns/SaH7g1ONw0bN/p
5gy/LYlDeLQ07x+hvs/SA6kfMF8buZ8rX9+mvOJfvcKT3HNjX82eelAFGt3QcKdn
zx94RNFX4XcxUT+vRYjVgCR4va2QWQrzCHyuyqvlWWZ1ZGDN+ADq3JLrg5/mLhSu
DPUdr5e9IDFnPfpIJDtYHl+ujaBuAbBL40uKeOZYpdI9wk8dzMpugNC6O0bnlntm
oopVtzd9+6qpm1QQ1KBVUkx/XAEoVreL7KgV0oMZPfmyZB7/sQ/qXKnzV9/K4T7i
jyIem80IyQwdRGj7Oi68aG05asXmzuLzP2KvvlvYOVs0gX8vaOdWl1FPpuvVGIPB
VEePTDadGtKpRrSW55Xzyetts5Ybd/eILrxBmYnxeLe7x82qmOEIZ3QxhGD3q+VZ
Q6gYBowq07cVx1o3vk3RvhiSPZqTCs3MhBpxqJOhqQksGmiUXIPWmIXl1goHUM66
s2EvKWK+VRbhy2mmQJfTEpgM/fhLo5Xp6v5N0YebnDS1P2WEQlKZF4O0Vn7kWmOa
LeG6u2wEm4kkY7bNpUyDFlHkwOLA9T4YNauaAZJpX7mi/uG2LST2YlhSzIHT77bA
HIFSrh80vxdUYlzt1SpAYRZnF2GOWAhJHZc0peGd4CsWKHSRFKundbyFf1TRYSZe
GnugdKi+RDcAxxVMn+0+193MJTPwRRHrBAlkNbt0ThwaNJh4kuy7EKMGQQ2AKKis
Y5QD95Xzv8Uzl4j8xlU0W4+L7+yviD1vNYyorMm+06YAKVnfPEHWeNdsX1v0lwdU
sgIesCNQyCfJn1kOG+6wPPViEyBUVizRT8J2EJ3hBb4zip5DOJGol6w+/+XEzEUI
rBJKUeLIvqydAMYG/2Qwdc89cNWELXU7PiMIOTtNRLl9YSzKgpe8KkOxItfE5w6A
H2APYv4QlSL8ZQ2DHO/h/ou/Fmm3c6HCWHEB06WbkdSCvTwAyu9zMMuCoudPtx9c
1No25k8AXwjd8Y4x9YIiw92S4XMlATRdq+1o+iRwma0K0C30sAWaw5WjAg1XR9f3
R0Mk1y6JzIZRhygy2DvSAAgu9t2MBxTup4nCGx10sjDibDF3f+tlxSGyUmaj7PM8
P9XMe089LltLEiqrMDSQES3GzqMeb7ZZFv9AXlZPZ07+tL/hvVq3gWbs/Xt6wIuc
z6yPoaBfX3FjeEqLKQpsjR3R15cm34H3aVUf8e6xiOtlIHhofP0Ex/h1Yq334gAz
PhFQuXmRAgiAQVoUMP6K/dMjDSzX69RPVSROvDCYaqSAjYMB+/TAyB+L/yJ6DhOe
DytWq0uQ3yY6Giag6YaSYXpaKRz8UvYEPGedPASMl3Klao9jKNocgf/rwAs3ek/l
46ZaKhWasKK7cyA8Ssrm9ihonRbGPbIa8D/i80Az8VggL/foiCocw2Lw9Z2zapv9
spRJHXrJHz+If772AC/s5roSJhl6OlyZMILrmVz+uz34CVi8gq10+UuuQ629xEDB
YjRU6ZGOomUOqUXViN56/u34gt7xpJzlC1mlR1sXOxyEcEZ8C9cBDdEeN6t/ABUA
OeVMjre8NNDeWhQmI9l/vVa4j2yv5YVIeEW6zxv159bkB/4Y64C4ukv3OBRVUdeo
s+Q7D0pEsCG5hcgtmZVosj3+Ct6CAU2Peovw1EjTQWSsbAdAur3kgfhmjXW5RVdz
dWSIknOkd/+V+L32lUtKJetXKou1jcgIIcIk0cX17zy06xpQEpAuXVYiCklDCck3
PmtlJeePrbNSTdxUgTQwtI8lM9oFXld8PuxcOigeFIcAdF9UBebUTSMOz0bfybTK
SUM5sYCF4qbS5hU/OTp7GzSJp/qImnqRSIN+5FKJ56n5JGCMtYaD5jqeT8bMgzis
z1pnC9QqCR4VP4tGH1kS1SwV3ca/Erp8c5k8sURv54iE4ghtTvNfVGpIaH9t/+p9
oXVVp4LlmhScLAQ0ejfdY45J1dJXEW+xkZrAk8lmtmuiRbdy+KLQeBwRML9I+m+4
0K5GFMGGPuHVh9fimiPn34+0A9GIhrrZrFCtN6nsBM9f4mnvh9yOsgXVbTPLoklg
COTTDspZNduP+jsA/NgwW6qoqhT0DeFgIJBGNu6Uk7Z6CMaoUbQ406JmxTzpFYsl
mCI8Z7rdJnOn+EDAPH8irsV62OtKbKB+fnTaiTpNUtO2RXacvl2ypzVqF7og9M+G
R6LYCC0GGLKIMSeX4DbiVFC/C5ogzSUuu1rj5Qh03LWtFGd+0CcQz9LmZmDeoRXH
n1xWMnuZ1tSkJ2RcxUcbQ8NxZ1wzKdLyuiXZetpzQnUNFOAZkCtfbJatvsEzIBJm
4ux+6ehRoLs8w5v4qEv/djrY+PW1K69VB4x/fr11ZFvucz13OaKNMjN2hhJnXLY/
/3soNT2szuHrpSTTCoegy5QSrxFqcxHDLrZDHeRYKdYsygYpzlKEuqQ6HXuAwVJW
B7sSEaEC/OxoNDHnweHru6m7uKZRioiw//G081EwBFIhRP0caznXlJi8BXrx8JAV
+sfgEczxixyeqy83qZb0RGrfDqWc5sD/njVYOMSqeeFGNMlqPHHkHzLSxaYgf7ap
RJ7rGAVJUmodqdYjgUw8bwPOtJCHtaZHZ6y6hN0sZc/1WdHCyicA/xc9k39Wx9om
CMT6OlWGsNLeF05LMvIK6ECETH0PO72SwShLfNMX75aQ4KPpaNT5dw+6GZQyEFc3
QwFU9Hm4B4+ZGwAaLHEYIb8i3fzsOfYLcENEmEVrD/5VK2/ZfTUzGTyV7+N+SuAc
5tC9dinaKkHb+CC38WazVclt5CZUQ8sOmR5bF59PeLyLjbIOXqw52PyZlLdRC6XD
wAqzFyWhacZVFhb2kWnwZ6qW74wjiW8WDxLXQ8QxiQyJmY7KQLbr+BGATDqV63fe
PneJkk8rEwBoGhLrGHkKwt+HZRltwimJ0jbuk2ttcVATnzB1q1CkDTp3l7ccDfnl
AHGf4Yb5GmelUzIeXccBdfLA6y4SQ1zaT+sL4/5a7/EzhzirH3aqbFs5p24dKNcm
iA/OE5EWGjWBInTW8LJu1zec+6S1NkfXDubMzd5uXEqGVipYRQ+hLEyxHEyxChJi
JEAww+oPSUF+gjAjm/pmcX9Agupf6ogKWfDmQE8B9sRWEpjZmihJ+Yym85xGqCX3
aQA1UhJp69bHAEI2AF4OMNk8DazvKdXCiwVl4WlkqtSNAgmlEqctjvx9z+TtMfQ5
dLAJJkR/Qs6dWYHnO2lkl+XmlFg48vz+fLQndiscUylxTFRz+R+ei+oBjfib14e8
FXJuiro4VLW7vmL/Q8TqsfnrWbtO96k6D+eHDc9Co1upGR1Y2h3rRtSOhaF+ioVV
1Zrf0xhL9xtQSSjPLeCL1jgPe9p/AvV1TCSv0cXV6b9J13Gh/5WOCQQyKg7dIU/O
hVG6gP4zVRQe2rA1EpfPEPi16gw5zsg1MdwkXYi50bNibh2A1iNkh960lEkXY7Cy
oP0mOnPsSh6J3kl3p79FMTRMB/mZir7uQvcVzTYLxgJHp+4+SnLfoQto+RK4ivNJ
dh4q//MN/B/zpAd1ennCHHzyr59tQ7YPz5cve3Jx/Lx9MnwAodHpPusWcbKf5zoG
dzVJ5Rq2dlg+RF8tN+KTn9l0OHIJX9ze4Lbb1W/y7pYdeC7BCaC36UW+UPWYihM7
KYFislV1MQufUuArmkahb53MJlOuRXyGu589xThTkBnyuyMZV62mRZiyYr5fPL2j
fAR0vwVVefgeYy5Dz84tlSo2rfDAhHRKOm2MwUvjPs4mLMvVR94ror+q4ftySVCL
ENRLMEeuCgkqx+VDkPXLjsGf/PaDcmYUkkYY5goR96txOkj8x72nKms5hf9rVgJu
5Jt/HCenOq8DFNvTlEe8KzELr2MSTrmO60bSEAcIIlb//UaaFetvwHxI6B1i+WWn
+5D+4PkRoBo8Ywjlc4Y85Joggf7WBD1wfmZyrcKJa1QxY1YWda6nRXFDfzQ8q+VD
Cl5mvhnD4HBy+c7spTOWZ4UCz10iYJqNKSjIM14SklfwLYNKa+JYrIYaA3hiJfo7
yESnzfvX3GxCgTAmIXm7RYzxA60UDfjMD6CEbgEm3Z/A1BF6BIMHnePWdaEjWJ4U
GAa9UxZy5BtJxIHDEmpsgPUT1n54xJKnqudEWUvDiMR1OBsdzNj7zvbhplx8v1xc
VhOCivNZEaRQNENnHEPd5EuVoF7Xz/qdrDESfyOzn7bX5RW+yWDzDiBLgCK/RlMA
f0+1q5UYtq6EoMOkerSphUG+tOxY+oQlsKshU9rMEn3aBC0VtswF03t/ns+x6A9Q
1GrBV3oC6hwugOQQAuq4a6j8TjKnxvXSE9AJ2oLO9Z8HwFyNXxL65AS8f4KP0Al8
U6CsU5LPq6jc3S4VMmoFjYjQFo7tQ8UTn1I2QpUDs1dtoABbzE4pKT6vm9Gz7hhO
WBEPAFZExgqOgaXgLq7fLoQiTO2Uw0mj8kYPFPXabRoBcgQwXP9OghlBWqP4K4b0
H9bNmPRfUPOs1FDAk0Of9vn24ICtkcy1hvPZLC2C2ItuL7Y/V6pQxJaKSq3VGbjh
rgThplYamdfwm6gfTheRtuzoe7DKJ7p0wpbjFpA1JUgCkUV0rmL1VPS27Sn/GpuJ
in6fwYai3aIkDotnolIJ12QT8bBW+4dfVeq0qkJOu16VLeVNoAI0JQe5YMzFP8PJ
xRuk8WIpbSsXKz1IFfUaaeOiSIGimOq+u94KniEzNYZSfwA0e+Z9mKUf4r6PVyHQ
bKq0Eyxen3ko+ea9QBxR9T2FK/CQiOjML7tbNLfP+MPzZzlaUeDpIFnJk1o1v+7s
lkiMsPbQ4pF1BKzL12KJg4NPo7MRqymhjvPcKZFJe1V5Vrds82hPTPXnO7fRdUyy
02reC0c0nsH/nICKGCo6l19TX5a7Y3GsU3MrvN8edBWMzZ8xD4tHE3GtuEORiAfq
8BmYXUawzf+PJbUy+U8d1wHKKUH5PJz1iVKv8NQZLkT6wJgLsD0FzlQhpvt5b9GM
iaJV3G85DYtmxyyhqnZqFBsUL2qIqoWji/AbnC7/ecqMKevJ+WLEc5PBpkFRKnzo
shXKdh8/ZImca1nNozdsl78CjZsmjekBkwjl9wZncKPWlcQKkHoGrvoiAllZRBzb
kgbBQkJQ8RkK2oYywWl5aXPbO0KZSu/nQbsocpV0sGBYBsrPGrv7DIUVlt+5QBRe
DxxRQGMRxj+ZqRMfQnko4TPZ0BDp8DkxuwspGJXYEpcDg42RxPF5Q1mDVen+qTdm
hz0L8OvoN9WcQ/HZ6Dx2REqM62APL3wnjM3WT+TnIF3vfOkf0QD4C+64tDD8qcf7
U+2zAE5pCobUz867DNkwg6Tjg5VkI60ajFsKr0/wfbkX+ka7DkWeeU16DaULOBdB
bANIGSKV4nxhLaa/GiLRi1JmVk0i5cSwSP28tAkP1s0yzNYLMz+0HAS4AP9iJa0v
5OLW+nLabUOxywOojSHD0F+jJVUtpR421rOzTedJvrKQOO1E5IyVRfO+CQw8fFeG
lGWg2tKgxqQTj8m24qZvV5Gp98I+g1CmIe87GjoSu0wd0P0jlHof5hu7wEqDQkDC
nUeqqsMhjsuz6ohqqSO4CMS9Z6iKZUuFJCC4pzp1P5yO1Y/Wb8ETv753q8t9WE/n
zbK7ruiIzMVn4KelxqYm0DvNquEXEZcKv1XasBQQPZto5+wwiWMLgESZnYOj+YZ6
dsaIdRIHrSNixF7ESvpfwsaGQK4ejUufreslGKanAJNrtIVlYtA4V4FCSVO43JU9
M2imr07SP+ITlsfpS/jlgoVT4yE1Nu13vNqXo62BmLPsr0DHVdkzx5BsU2pOGy7e
A4ApQ30Ra8/Q0vaeXQIr6P+0eRDVHSiVJjTWJSyrZVgdGiZ0g4K35IU1pZdegTSO
C2gx1TcBz4LYZxLZuHzFzXNiCyhjRMfim53xhm9wnlRj5un3Y+nEbjPKokXypu8j
IoiEIREIMjm5mFkxcFqDig7VCps2Qh8iUPjbV+HHbYyasaRPo5I8l4KRh5nSgeV7
FIGa8flsx930Vs5IB97wpfDU5xZoxz6D6TAU+NZBYYcPXKLtt23VA+VPv3fU5mAC
HRI+EpKZN+73enbGgv74aDxweWAxjpCicalSBJpuynqAU35Tv86fit8JLjVn4Uuy
HmpLGUP84/gbcLyXobKjHCUC58DYJA2Xfo2UNLfTtG1EHifk1CblpSJtkAZrKMjs
dAMG1T5dbgsx8y+DnHtmegPKYFP85pbTs0kMfd2gPqfHKVJaztQITowK9+SeEVHa
dw73I09YaXGjBTqBe1pKdMDXIHrIjQxWlU/W8yjBBM1i8gRivFFqQviNghh2rSVJ
vFqWxDeyn6OtBR3fi75721/LvjDxLbbq4VZCDFeKWp2B+e3KPlp/7NFP+WjUKest
6URv6Txcmz9nZK/+V3LT18jV39JNRn5JWGp7Guc+wqDDQYTxltEazsf4YLNqQfPH
jlM/o5vgAK/fPjzHetQmrQ1Et9H4cDVK6WOkLRhUGBQolPMePLvDPGhlwqfX8Fra
3CNWQNnp7jzO3hRNV+/kLhFxIwkthKIxaDWBR8cFNtiLIP7t2Y8U87PldK9TwTdZ
Jhw1YQv0iJyUdCBjSiQkJ65Sl3a+bd2WLS3y6QSciC4mkLvmfAzZfgsMkwIlcxt7
PstHP7N8O7cyloGQr8LHmXXyAEpT4rsrSYzrDDC/GcA6Jm04LE7nvW+BiYGVm7xx
04v3g1uTbgm+axLw/Cd1ae8oubcz2dJpGkqsx41klQbMFuF6q8FpofWcEmPODkz+
JLCDw5SnMmG+Z9D9yOckNAMmL39mNQfdnHX1GWZ9qRThItf4udKx+kIK1Y/ywfcR
RcVnsw10w9hbr+rgpId87VwJYQVdoDY7DJJfspmmwjxmWEWqwg+dbcHNLtDSh8Jx
CV45n4JdRrpFuHQcKyF0TMjpe6AOo+tasBzzHrjrc3BFRzEAg4KueJQW6dsbSdkJ
PvENAoF1N7qu/7jUa1CXpznp/xUB2lKPWapmJtPq8WZqOufBU0Usb6/QASKz7/AM
jWtVRJsROUcPfPLE6tSCiHas0Kdv0aXmEWqxty32KrEBN3Rs11DI98HWDCS2FmkK
UXK4K1YM5LbTNvDAZzShLT1APyGChQFrmhm3gb2IdRKFxUxMAJHnoWT124tdZ6n1
zFgzUl0ZDSuusU2QIqid8hhZ/mMH7gkY7j3lzQRKVRGse5ETxuO+Qhu8Fm5puSrM
eHz1bq4P6yBMquLysCLBLjt5TUSmQ2728e4N8Ce2clWMOAY2izMdSm+SnzTpUZDQ
LpReCxSMA6oExVWPCSHGe1+leqmaFyFgkVvlm3y5bpE1G3r3BPM85tjjMACZyGR1
gnBggqco8IsL/HrQn6J4Q1cro6L9+ScJRmEAli7OcgofSIbdKbpoOAtkVQDvaAWv
06V0lKYFIZYoIuLh9FvQUG6EqKH66UF527mphWCU1zUBjSgsY1VHb8gskDnUBk8Y
FRkT1zRgzi67nRDNhEDboEvhQuSQC+aOH74xWUhHz3tr8+8SsLF+hP8wzJnGDrrK
RynyYjpA8kzhodzB38i+Slegwm7ea0Sei/arGZXC62ksRRr8McNlrGPEhFfWASnT
+WPZCU0nLaks8feB3iFQVS/4GgYbVEtXguKUax9Qx1//3lnMJr+TPFYfl+TVt8mL
f9hrMtNHeYMjOsv1SggudFKpwO8IfRMqABl54eaG3IdPBjVwlYyaqcSKNiZUOp77
avfIm7QPnA9Bm5+92lIPc0IMv0hbqa6G/RoODMCbudxHwRvjL04DyzI3MhTKB254
HtQv9obLJXOPWEujqu2VRIyJdq0vLNzQ2g/aZfJhtWVeedmDSjD/eV79F9ex01ao
xvH5SmoBf2UOHLTeUEPC2ydxHsEX32DQCuyywlHedldy+pl2yaf3adNlzyCD/LhQ
0mHyVihowYjYI7QmJ9+d+NEtc//9CPhPkKNjkmlyBQex0tMJIGKRpxrdPdvGswVt
9mm5Mv6QS6XXX4IeVDP8VS/fkumPCI99OJOrzHnoP2dTLCzLlJkrE4CB8vIfS6HA
67zH4GQlma6liYdjIWMA4R86Ph9uiT/SX1qw51CtIBbQRT9nH+EGpu99EZQurkbh
RJ9Opj8KVTRM135W4/S6X50Y09ZuHaUgFu4zH0OsiJA2VpVV3I5XVRGCUojZW/Ck
gv9ycCm/jm8q70dCc6KSZch7vmX+HbqEjhvWqgtJxCAs27X0V3XVhX1YLQOnjYLW
IKKKXykSKdhwKmDWPASWdnZhuSViMl+QvUazRcUkWrSfmkjbHPg9uKjecU0PEdB2
zuS267nj8CFy/pUsbE56ldLG82mNACHlQZScqKRvFPeRxSd0huuCm5UrubBUL0DG
fI1MxeEsp2ErAPCE1HJ+swmxmZyFXeaXTHj9Mkg3sGvFBX94nIF1uoUGDMSLD+os
n3/ttlcU5SRSdiVyvXVA+6o4xgwD661uWlpkBwkWgELozJS7fTb/VN+R1ruqYXf4
BUrLT6fdQllL+07CTRTZsh48soK+e+7a+qdaYEybT7dYDq2ULM+rcWop4k82h3NT
jcRQArqKXYi3xojqmh5GdLvAXxJddjDdaryIBaf4Kpdx2LIHWQauHvnfPY772OIx
+ThWYN2+OcJVOu+Xdzgd/EQBg8/f+GyLUhnLvHaeAQf9B/TKnTExgAcpgaH0HOS4
HhSIThldtzamOQ/6A9Wln2U5/CY56oaLDb3cd/YxYvMwuDOeZ9V9WUPlv1ff6KJO
Y7+AbAHpZy0kdgo+kG/tOOmuHis/2QkRRnOvv+Q6wqOO5Tx0xRUmZXMFbsccA6sf
XciUVFNImjdqXnRK9gPWXenwZI2aqF1sDCgx/byWrLxVmhMW1J+lBV9aJj00W8CJ
RwT0SfCwIc4X+yQqEDd2PgSenIWGHPn7VvwzAmQq8ZDvwVoPwi00Rk/EWCHDsBSv
3CSF+zf7VZ6drBAo//yXLy4LS9tsMK8f9MXmHcuUFk8dyATRncWCmrruoxzeb+ZL
3CAoxjGlVnaqPg6hAEcSnPXjioAl6DzHmtrWXp9weWEu3CtiOnJweWKHsvYIuvPj
grC9eqedFKeDRhApNSS0JgOIDPhdlVNGhBkVd83SV5gjGfY0a2c/5nTVTnGmOjWu
Za7aX7BPmOXM8ro9PooFNvVKKTsDSVIbObxnU+ta0fTdDDyJLYEG2ebKtOixlJiz
+g3VURPtg8qmiDsTqnmP9s7Of7dwIYpikC0UGOEBbX7lTxmbkaKvShHlQ2Gqdgl+
6Rr9dah/JSe/OoGoCbwEIefFJPrvH4ZaXsedDaziuvfNVory8xao6Ng8EbouxORX
96g2X246JflwzzgVRKt7fgWiuBKCSUddtGupSzvjX/DrFMo3zrXIse5AKsebUi4d
ebb9Oqm9EZLZ+Sa67yFQrYu154whr/keGRwxnRQaI0z1rCiSuRsRUwY3YKzUkPQK
UiP5gWbXcWNkd8qsuCgJFV58pY3d3dsmcSQsjcdnh5DchU0u9vxSKYLysbVb+7Lm
gtVSlBA9ARjAudlzZTpzs3DLIiIywCpLZfE2KcaN7ZI/zUiPv34wmI80yxzuXmCn
3OEaUcr4w4KRJ73PddRc7bBtQwgt2NQT2JNxBtN+bUZQ3U8eJoUGWq/Yvd+pPNfQ
4wj5KDk2m70WbYkAqIR1mUMaangFR6ixmMTHxZOmDrEzMRf/VsfAO+dthXpxPGOA
t/ecwx+QCxZfbiR0UOT1eyLRSQ0CMTplnswwYl9V5XI69yuHOxExNzUcE1GX0hte
+o0GIb3BGma9sKqg2j1Kac9bZTCDcwC9Uh58dnlZCEQNTTJeuCSxySvJOMuS5DGv
t1Bn98c3l3T+EQwF/oEXndqkjTnPRX+IyvYy3RLFa1J3s3sjDub3xhcs+QYTXbCM
powLa2YU0WDBmUw1zL5yGNilGkPmCV6dk0ZuYa/jcy1bpqB2Pc++mzcCpDE76B7m
JQAj0nnIKrTfd+iOA3YTUhA4Z/l7UEI61JGstsP2CRyUf3WWnPrb1oq+CKzJzYMT
Oj0rKT8aOa9CL1qjbaS06o/0MJLbZJ45fsr8aR4CrcJmYUmjielh5eN69f6vqQBf
u0ycElWbB5Bp1sIhLPffZuvP8iHnFAm0K1n8kTAXHqfDMF586vHVUKhxAads6zAW
8e+Z16Tjf+dEdT704NP7r3Epl18QoTpAhYMTFsx20K5DcYaffs1DSFtmlB8ffW7S
LbK+FwoX49fU3hCFQWADMfUGVrFGH10yHpZQVBiQlbas/KdYrKnYXKyjpKL4a6qi
Svzw6WM8wbj4qM4//QL8xESvDS/c0GOiSqG3jrxMjY27e72EAIQlQ3N3S18I53EV
f7Xrdb0GPDV9d8WU0ivVr9dfhwlj0uddh2/YifA69n6NB8eMNLcu27EmN+s4fvRg
4S0NOc4NFK0u6wQikYnMmQVcOcTTS2g4kMqQHdRHOVaHd/btmwzaxcNmD/6XOBhc
RoLuv1q362FjehyHqV0mqIB1X0gyVVcx4XNhlg6WjtGOwEOvsPOScS3O9a8nPWZm
ZbQUgu1CCT90JOn//E5gGnag+FCFv7pb4cbLqQJw8yoZU7I91KXrOdfvIB8Ly8cc
9FFUDEUoWH3ilE6ujRYrT0uqJJ6DnMAL+HF/SIiOGJB3ezcqFvyCgU3ESUax/qmC
LdXfqxbip+x3gGA7ZsM6maYGJ3qzPh7Qxiu4ZJxmm3Z9sDkOVZMDhMnYPtTc5tfF
COYRXR3dcvGKimZvu4KXeuwEseK2u9tKCCjUy9nQNtCygbeuCEXtzPmgebsydX3P
oPKcSqa1EmNbenoHCMn1MDQKRiDqbIS4ljm8sbHV36RR1pyYaKO3OGwtrzQ+pLxz
+YG9A2ZydhtbFCX68uvDDv7fLwS+tMvonwdGLjFbuEX56fwU6MeGwGeTWwLONi2r
9gHc9g5x1/I4xExRTlOC6PBHcExwnltiE044Ce4PgH6IC8iABJbtnTxQOdBmHL0R
VfLFOztg+lBbm+HLl4xwUZrcIxog8TkoYMJLoKwLWlTjYltuSYgNAs4U11Ua0gLW
s28d8wMTTnuWWb6vTTAS6JnOJELuYh+GxtHsAPuiS7rEJ9kVmQUwhl1X0uNZDrgb
ndKw31vqkZaiux3OssuYRtpaaIY3Z37hIEb+T20p5LfHrX4BzJJ2qiUBLNGpocrQ
FlQbsfuxUwZ1Mjxroxe2zkN0ng6ifCn2KzcO0oTEHgDvMODlB2gVGlNdfNPEQXGi
55Zs18VYLK5C5urwSo9opSkFqNfDOJJLy0Ypg+YkBcJqjZu+YioN6Ij5xKu8CEpQ
j5KAiK8tDM6NtavHiSST02aFj4/qednXlYfg9NfTemDNopfwCAtJCv3WNitnCXhs
9BYV6jH4Cjc1+oBBKTXxzuNNhaAg5oP1pP77JbNKCK+bHaLWT1DHuEfBf6fgHex2
mUvkpgRbpPk8xlLYpDNVOALmFlH4qPaova71dI5kyDvieONFCaCYRxEjrFD7a4AM
rPMqA/TXo0wx/TE9WtibO9+i2d5ufmJfgKFSJf/UBrJ9jPGcA8kWqoE+c+9CAVNe
OSjldBA/X5V69h/ttQNlanzsDiUI249KFHVVusFvmn9bQL7VC6uUYqo/TtfGLEyv
V+6ffL8VVOYUxqSRVlElXbhzy3csojqF59A8oEeSD/q4lB3t7RHNT7V6OctatJIk
DlZS0IwX3UBKZsAFPb1G8oBVhjmGNwzTR3CdQ6rrtuaIZBOz8NmHv2qKiAA/jy9+
bl24MGvAKtnVB8xNabvi3LIMOWdc+C7kvlxGCNCly3WoN26odmwZDSPYPcwJaLMX
ylxPRlfGOJktd8tbP6cFBks9b3XsdJqWZnqZ5pdjAhqbpCNSQfauhZwvSFVmGWD8
dukUO5sxq6m2xIgUCVHeKbikfVsQHjYo+a/9Cz2ho2FYBFjsECL1ozl3u2zK0d/J
2wKfU1f+IoJnCPLfDZNtcIVj8ZfHg+I1JfmJBiPnR21N+ihGsecgRQ6WuGLU9GP5
/iQ41Ub3tnSe6hBLf5KHMxk6pxAfEOhoumFlITZDc7zQKMmXT4MRhg+LxY2Ia86l
WvOTZpoyujxVsQov0Ghe4mRzU8V8WiGY25Nf2Q7Td2FdOao5xnjgX9MhxuvozRr8
9EuK0XnZIyiN5LijDix6XpYGfIFBYPbPlP9BGpXSRRyErcpMKEEf3pjOcRVYQ7Mn
RpPR0APXDsXbInM4dpfXSdRvTWTWofOMUu3yeSppAahexEpFoazQ1lKLeCRolGui
MfPjd4IgqdS9mCyIJWTDpFhdXYJMeXpWuxs4Qs0d7xNawjLp5qt9ELX1RR7U+tvo
45VEjqkccKT0S/gvKt/UVuDBvq0W7gyU8JApIPNh8/K9TgqUIt1S8yeoItG9YeNY
3IgJ/aYG3xBUb1SK+Qw81bF/Gf+ERUZEpzkwh3XqFXHI1A0EnVtVC1GNXVsET1zN
2GLBJ6W3JRGa/beJcyQsxoden0g9MMGL22jhjPo4njWbsYl4HqQ2W0nMyrO3/nrN
+tLZHk3rjDjdlrR2s5mgHFcN6mfdvpZcvYsvMsKwz2+y81Oqg2AmvCogYNx+d/kW
kw8CNVy4C/ELm9DNmNpXRG12pRRdTpHoGWWTzsmvZQeZCvyigFY3podTKosTjN/e
BjB+TJThCMhmJffC+Pmd6XuWqFr4pTUTzWxW6pRHPP7LlUitTc+smbrc11gIZkeZ
geYUhYDG8GyQwTHUy+uEw5hyo/7U2tR8NnmEQ6hCT1hC2+hfi+u/eVwigRsEZf8N
l8rpNF4du8U6Sz+5K1xmjZy08zZQY4QvQ94G3VRnjslGCPjdRqNxsoecE3dYc6/X
2jMvv+7Cl0T44ufywZsnDkfB/KaEQuGgtEtPmUzz15W/leWsdJUQyAuJFVvEul11
tKJiMmovpyvkGrKs4CvxgE7f4g/krWvbKWJnX+Ll8X7iSM15cCh89gMI90AFfm+b
qXhRgQVIMjdSm8pNpt44AUGGHcJvHh66aa084XLpubWog7/r87fjIIZYi9QkG2rm
95zWrbiXNDmdPlI9riwGQyOrWMVPlH0RX4baU3Sw+gJqCetcKR6ggSzDGfN4sn/k
pn00SQ86cLv2kerXMp8dj5pPC/I7IsP3jIe6BF8VE1UeNPng2IP3ojz1BDt9S98A
ZFQApLMOHtURPekrLUY65SrmKWSy49dTiMvZXBKjwqcy/eqW/bd6IqBfdOputzjP
andixauQK4i/6IXMnYPJ7ap9dkNLdYKjeWaHvnP/4FlxToIdv86V1U5nzjD+m4tM
pTUOww/T/0ZqduMu5A479dUiagSEq0rpeWeaoNRufA62x+NEH5UimWjZ7ePFW7b8
N4XFVJbh7nytY2mqTtrgy74Got5OJgdzuYYX3ikbMXlhY2nOgKb3VBrO3LDmnXTI
0B1ye+BXSvYtW5lqGbEaIiBAdqtBQsvsgJjvO90YH2lZddt47IdA73OHcu5vPwtF
45HBIlaMIKPtButEy3BO2Lup9MZw2/mPNsfox4JRkZHD/noZAGGDCIw3EuNbJYbR
PcFqsjUIKM/a5Ijx9znli1iK6pqpJG+Ux373tUgI2LyZ7+Um/nlEMxG/VRtSqoO8
YQa/B8GqSiy+Yw7yaHZ+Qp23aXU8c0YFwtG7+aQm2AGQKg2oBMFeGghrqmiqXog2
m0ijTy6BFywkXMa4jdkTfm85aS9G/KgKcnHU6iVxafv2OlhaEogvy30MXPHKijU9
crPdG9YivA74JyIDm0JmLd7J/BG1NqfJ4K5krou17SbjQjTWWyM26Oi3U6zVgLg2
iw4Y4po17MIKw1rXY0WSuta8d0/9Zfo2kMFDJAZPj/psdlHv2w3hrK1BBNCyeymp
e9GIw7kxvNPEX9diq7lpdY1ryRqZnL2zyWtS9LAfonEWwC9hdqoEUtWFz0r5/4hd
DDGyIA+Q9Ax5EyRpRuNX1ho6tM/E52wGeWoalrj690+mNZHDaukqOUWRRPESpfg8
OrfNeZ6JVYbXQJZ8D4LX9+dDXfrd1sFvLneXjkhRVN7fINRQIMLdtgiP+skBc2WK
hxoMHMEEmqfTW1jdV5Q7HHSaYfeFV5WC5m7+igatUuDcHapS+I1K5y5mn0+m7cJk
uVQq5AuTc3S4b8LzFlWvGT795c35ChmNVZSTtdQGdsU0I21JrKKob+1QXJhlhdwK
wCMLLVAdwPmoGNjEUyR1VoyMW7g5MMez9bxaL90DdIkAWpA6USrTkFi03XQ06GnO
yKeJIpiNoT3has8pJs4kcC+p9GQf7TVFy8UmdI/uiLfB8P57ue4UiZh29NzzinVw
MAvR8w50Jr6i3jHKEC7srkPi0v6Tlp+CB7gjs5G1Wmk4Yyho0uoi9ReQL80TRthj
o7CeV4T6vYRqWs2Eo9qv5h0QVZDaG0QgwXQXnWzPiLFptVY6xTduJkD3tOYb8ER3
adBShxClQ1G6vp6ML9TCbxCmjz2zVDyClKPETTTYKNcd1vaJuF7Grm6g8InHKXEA
MtOlllZVDFEbN182c4gxZfm3cE40ebz1g94Fab9KxoNmxsitW92q9rBqixJWAYF4
jkpesuweKAAni25nqJRNv/eQulNLGrU/f1K7cyzqDyPG8L+InQRoS0pJZbpPhYiX
Hr7t1ToOxedL9BXnBMXEJnVZhcIKb45Fsp24f49nc86Hs4gEfpNCAjBAUnKur7rI
uMLIAHXHGnaNA4g5tWn2q/DLeuNRr+BkT/maRe4ICZPzi1tzDxSyli2Xy6oyHHZk
XhIH3ijSwh3WhYIVed7gE3HemJvXR5m4YRdC6Pcmnmz5zwuUxm9dDK6SwfIbbwBT
Ai3TbqvhPWDzWA66pFb3/YY2bH7KlB1o4iTq0wLwLcY1uMtvrTeifT7vxUSBWtwO
hqa62inppSeGeuUus7lemBk3HyaKqrIiOH1WsPumC/l+qoWAQswDIJWA+kucSqMM
OsgJFurb/HwOkk7E0RuxJIp4Nu4gK7d8IwglbqbV4yXsSugyYIASioTAgQyc9bPl
dPth9sQk/aaBMI1St4TwpSVaayScAxfphug9bKI7sm6PiuYfNhj39oxhfRm5z0mI
2FsxU04qyr2b8ED+cF+8yEMjpu/GYHMOHbke3t99GI4MRSDeP+2Hie0QKkdGNFak
RR3B9JfoHUMgmh4NiDUmTC0BlZduNN1zf5VRQLU+dOMVvc94zS1QBehYP7T26RDX
J1DfadjBDbrtjKEklFRv4NOmZT8ERLdm+KlYuaUzjAspWUVdLGPwIfqRwOBx6M2V
RYSxhaG189ZpK/L63xBKFZtHs5bGD7bN8kaf4fWOIFXJhKX4GpDnApsKVRedOueS
PLvc8tDhc0TsZ6d7XAm40/T4VJjmzl+L5KeWCtLTlfBz4QzoILWtF3rZ7O+EEws6
38EFaAfRmFnNG2pePuWz6Xv6O8oanaoOl0Tf93sBPXbWfasrQn6WiIPgp1ctSrZS
272744iOFeT1+DZRDi3o2A3LiDVPIuVvBf4aftY/CYy63Pv0Iv9GqXlbBjSV602p
sapbd6jYWfoa6oiJpsJ2ti2VkDGFspv1A+BTJrmJvD3wVD8YFj43IxyX+pqmtJyr
iQuC0VH7J/kQz3DQ8xLFSXFEhiHDgRFcVjoZ/ud+qdoUXET7K12gwAkbUy3X5MeI
fina02vvqzOiUnRjcLWSEniT2JZwQ2bZEWaUk9L2Sb/3A67luO96emcasVVP+ZB2
rCAfPpKU2NH9DoyTnR051tXx1kNtP8gpTqFpLGDxTBykplyvVd173aB4mLda++Un
bb6A+GDEsu4MwkRocQNMsUV+bmzhcZTeL5L2pRshvdd87hcHhmZMORm2FfxfSxDH
M9FkPa9I1LF7P1vUkfA/VmtiL3GHYHgG+Upzm4uRePjZPDTGYVSAg0P164kpMCcI
3/ndkZ8dz80UckDUEDIzrURlfBFEo4l+9kDFF8Cl2fVW6E3AzsKkeDdk6NE2TePE
E0JZxCnokDUAcVZEbIfU4wO70M5e3ZlBu8OKnfwYKY0x3rrEsjLXkFT9uuUHdgYn
jonFVp3jDjtB3d14Sb+Rs4+jspJtUbQlH4DJI+SjIWimzMDvFT8mKniEsLdWAbbx
WId28tw/zQ1SF85eP4hn3Is0qVN/gR74MjlMRKWrX3u7k8MJSziuVYT4HTho/7lQ
vVcX1p/yQdqlpCMa0Zia0Wts3/sxB2MwsX4dxERPdkDnvMiSrUxAqjJMD6MCNrgG
GTtGeP7oZmHWM5KrxN3zK1hWck2+UroD+BWL+VjQjAN6kwyLYGbIBeJ9cBTG2yPY
mG7KUyLiMCwNyz1SdNDGW/0v2/dY/lT38DtCno68K3lq9Mo8y1veERAzV7TCXfq6
41WBge5fIWlmJ3DTTMFfT0xusrcLsYP/7ZA880B3jtAoc1MNP/VlKrjtCoycQVQh
yULfDkXklFAXFLY8pJm2NdtuM2gpCnatQGiIZ5ZYTZ1w0pLmnsRyzvYH5UTd9KWf
01hddpYoM6DzDYQKmkKI3NRmcEqrCMrgyAjn1LfYREpXtX+Nu5nrSqq7biVSXV2A
ntKFxhJmsGODf+8hKI8xB56tjcqnhJ0bkuh/JFPHPuMN5/Wpcd3Ikwg7+0dkay0n
ntIpK/ZAJVjq2hv03qkGdoLoX73TqrWGiGoYK5AFES1LGOLxeqIQry+IwphRoWy6
YUR+/dLm4dwgbSqbCvL88mq5NIEykuVy6E6rD/+1lzoqz10octX1rJ64pyDzJ3Os
hOk8NG43g7lib9znlSz43LvDGTVf2ZJffXH1S7KKS2/6rPjnzmQ0p+fuWWsoeTKv
dXtpm4nLqaU/yLJxSJqE1wscB6WgJ8swI36kp6X0BwKHqiUxN3lea4uXcYaCQffx
B8U8ApERHyD7E87yNe3gDhp+3y2t3un1H8kfDtHccVDs9X1ixFVI1lcq2E4q4DDn
K1IBxzAE0llF2XCwdbxC6b6Ozq26Ms74AA1+CRF6++5LHVRMLOXJzdqH3UUPJC/s
/hxGVKa6HEOIvUBqb2gBCgKfkbw63SvzS8e0zlTWDjgfTMQ5EzX9RsfptHYxJ7lE
uV5v0ydhDDR9sRirCGaU55oHWS/Bec/c9oUuR6r1QthcN59zQXpmxctLexP+xTJM
WNsh1VAxS8rnO2IoZf1Y8BBqY+Dx3TRxGoSvMlgjVcBoEuGI5CysUHf0X2eLve1j
wUCNUoZc0WX8eK9zz3eT0bouYEnjrhwwg5EO/8uRl8i/J3mK11AprdFQL224xYwN
f6Y4xDYIfEHQ2b8ChF0+upEfrub8tzDSFqTP0qwSLDzDrOhO+HJXmJ+w4c5UyKQn
913CEz/aRSPbRMPOemf2Jagk1YlzvdOLsCdKsXNsknuZSsg5lBt0K7glSIAkpiDp
A6ueSF5+7mSNSor/xHU6hVegGYJqDiBalO0uVIxUPqxp3OyRs1rntw4Jb3RBlZc/
MxxVZRWhotxLO/kLDq/s84sczuHfPTOmMpRpJZIDXQcSXkwP0sWeU3WwkeSlUxNJ
nUGrYssFD4ze0DjyNTJJak9Ue37Z3Gw6m/6yDjfSTHWPkYC3tE5h2usJ1Y5dTyui
tb/5E2FXWNzFVKI/y+koP7wUMPSXmdv/r909xcXuJOxve+jg1KVoJp9bdQq5dUGL
4/Ym/jUP/DgXLcR3Up0gSBf6B6lWU7u0R5ZMLJbb03qjuZjpg4llTl2phs5WpiuT
A0MHJBXrnZuqlFhQstPKsCOxyj6xflvc3taUzgW8pcREkATml1Uq4XV/TbGjr4ap
qoUCM6U33Zkmq//DWaoQnOKApR4TH+LhLRNCdadYSCCWQbS5UcmAcx+1gnSzSu4m
msecyr4kkpLnKVCWHS4P/T9RxU4rmSXi4o5X5jB7yNWbrgywGXiH00LKQiCaPqGh
JMXOrzbFtO4IgSNxJGgGGMGnX0xhHPGmqtXxUw7oFTFsb0vBKnNSUGwfh16Wow5g
R/z8eGokkeOaGR3jOgIjJooKT6CZsi0+mrkdWy8JbHjWBOl/Q1gFnj+Hcpa9B1Qj
FsWBlNWPkONK0mnKX/6/+SsdNfCeFNT/J1KzJvSIalGIbX5jaIWaHmMj2r+klQLb
n7DOjSKYbufPKBXY6HchLLwLEiQjmiOnGLmLqkHPudl5gRnJIya/W9IXS4FWSbrO
9OxTWnKdJCrWyNflBsNFLeez4i/RSqs0/PJBFRFV7Ldk4DQxfcq2jMBB95hlGX8M
30mthO48dBOSz0HGd9R61k0lQMB53MP5Qe6NToriopbHFgXoJPHW3M5zM4XagLjW
SCD7c87Sbz4w5v0zVdiCaUFlYs0KfvEM0OlNFpHOF44jt6ImlGN445JOFCoepaJl
9fVZZP+4v5TQe+nCUrExJ3PVAo75pS5Cf9R5SiSq/LReQuPa7/jtqNOY+elPa3Uu
ANZCoILTQZdqAdwrzJWRsfmTKuwWluEEutFQVhZ0ocOM4x/OLdKUepgdCT7gSKMj
DO/qE4UUoewObYqjfmtXH4XAC8rergh5L4MitWs+vdQqisgpyTjh124iHFPCGsWG
36k8lvj7LxoUvspIPPdrnWZ+5GZJ4azGzRiiJ+pvuogXZoBo8m+Jd2FaZfNEuF1t
g9fRdQdFuDnXUNJuJVz96YJrrGoPteOZ/5ZnOK2vy1i3pa1lbpJIkBr7Ol2LBWGW
MgJogB/H0n9JQyHkd/xUD7ylV0qhfwajHWqXkIeXROVtirUkAjLACBWmk/BVLKF0
NkJHFWoIK/toaQEPGWU/rceKMPupFky1yyu4XeUvEtBKPgMsKQlXTR4lfCndssZ7
wfGI3XSOMRe1OEDVXdwKNWe7+mPDj7hw5XKhPvsVvmQIEcULLXstoRzkkCmarJYp
2DrESJ56y+F+VLkwTKzx/8vR+L3no/vEAn+ogHkMIJ9MOR46SPVIQT84EvM111z2
o2Q0Q5Bsz9sNB9gX9O1AW4Z6WbiXzIuWFhRWx/iKltagVPHJ5acHOi0B79TaXGhq
8MQInn+HL1kaak+CMZDw14SGY0lCpH2coF8bwNcxWDdo7zx4Mw2kbttbG4VjJskS
KC5+feFvP+hmlzSVUJy+gOb8IWZ9oa5w9uj8giuq/vl4+nOUJVQWvJTEjdLsclrt
GKlJxRSqr+O6wCM7y623j/7vEzmGftEMErorygUdFEqjSf4neAk90urtBIq3n3fd
XqceJeZpDoDogvAJxSf2ARN7bytERSRRIhPChW8z+A4Oj0ETZ6IJNJjF4VZ8qWN2
Qy2g3jABKa1WY4hR5x/Ce/iG2dwrYv/DvJTz2lkKdRWjVV2g4ihDNQNowgoZoLSd
Yg1ixlAVGbMieMzRq7Uj12W/jOaXU0greGVLG495fDfywpIRczoMS+DPprGUc0tn
ZMOMRhEAfP9NSukTX7GjiEA0BU98H/iusgCxf0uury/dBEaNhcsTc7Ct4XxJUEOk
Bg/NGzzQ2BSwetO4uSbPEf+un7xKcs07FGOZqrew6muP37kqqLh3X0vp2yKmtaJK
BD8y6+GRzpfGd2b0hKB8RlipSYOcHgGI9AIRyruaQ0ioZvbmVx9EyZkEhvJaiNEl
A+UucLrNGkdCTgqW0FlZcVCK9tKmOEd/COs+zRqCd7RRYOIsckkejh4/ev97SEgh
c7hd5AN4JoYGFA1lgQwZ78TWz4WI713VIC/xPR4gWRBDlqLJKrfHfsRAR9K+iiUo
//rPAuLboUXalbpXMYcRFg0+MWNM3ivKe6hIj6S8LWbPA6Jbtb7dLKGJ4QBHdvvl
IG4ojkK+n8mPSEurOxyt0zsLJBGtjwuTz/+AcstApDCc8WFeOf9errn0mpMv0WQ3
wNnO/jzybGb5+HxC6OWnoCeu6IMTHALn5b00nNdC6eOzXMqVtsBC4gfUTpkuidCs
qeiNCwKiKBylwpnUiI8ofRTlq4/+dxJ15FYO2QtEPhcnqxS/9MSSlpe73m+WJa+/
L+mviFCsZfVEvIVr2QdZ0hdUJs7vRtdz+VxQAeDf0ptZVMBavQ08/xgq5nQBYJ0H
x+vV3dB2Yvvn/4yxzuOPRQYX+mEzHEGBoh812VpNrLnQtrXqQ1aTMcqZ6ZMZEMTm
NdfoGfgJmqj1biiVkrUJ/5NVXX1v74ZqYp3gGb1IR1LFRajxIAXMNBhdhffq+CJ+
pDqgCHv2OznFCv3XxhMTrDc0lZQ8xiv/WKKDfgGTvlX1PScjtj4C1JDM9fbr9Dv3
PUvdSW48SSn4bL/aZ/EiIVZ8fX44KapXsNK2/tD59KFNnjDwCdSH1w2FQysjAykd
/zc4JOp76UYyNZeTvOr+atS64xC6QHbRImyixzNCPH+rqyLTtYuapyJ23TDxtRlo
OgNZuRQviu9O7LyavWOKAIooAlwvrfQPIW7wX3ciso/8QCXVPFoLQNU5GCGkvLSL
ukQiZPe4Xsv/H8yuLBthU9SO3entiw+AmsmAUY4iRaGYmJdPZH9do9hLiFjDlnB5
XhX3t3fvvPNG0iFM6+SWS4Imz/omo8jPsFG6AQZpTVKDZsCq2EOnQwfG30liTaSK
yjALVlYquhbZev96zeEpwvbLqRjcS61sRJ4aeJoK4d+GZO29XBzHmSmASv8R5COe
jbEzKvKSponWYKEk0tDOR6EfI7jMlwp4a+G923jc3LnL7x10i00x31fKYJNQJNis
QojuDWQfOqV2g0A8CyVF1pThjZsrgCw0xKvxUBS1uWJKQQ8Q/eN+eJqqQ6Mt8Lkt
/qwG4OG2XeSz9lhFot+ywDfFow/dMyvfKT7y9+q+o8xzWv5n5PsyW+6IAMw1PBbZ
Do2qHThwLDjMG05YYkoLQX8HrbGiCe8+HUuoowrPyD50CT0NPq8edhDOBw4wNyo0
RtQKf5vLrwj3gfivVCHQR6pomdvprJZTRwTR8/yzbDTz75kTkWgK0zKrUZj77xvV
fGZ/MUNFfLl+48AIIaWwiMWg6XijHSJE3/2aHC6nVoPcw1fcI9NbZRzPLbsYx/UF
FyDfeRQyyG+rNI0RD0i5uR2j1HDY2+/cf/XfLdJEZzbbt0YvFaiO5TziekU+dhds
e6hoKkeVgu/kTTJbPc62BrYuAnRD8H/ykOi88asl6uuL6hp/vM4lCpvRn1reaNoO
S/eGmvLIsLpwN4rdRPWJ/GlogQu1SBzUMkvqB2KIyZjaKS9QeZY8nYF1E77cc+HE
QH+G4wYqA0ylic8XAL4TdXtfUPVkRuAym96N81YldrfkCXXvyU2qSB9KDK1SGSY3
m+/MtPRPuWsIhmsJjAq6G4B+wbtOrzyhk9xjs7o1ModKOEXQy3kDlOEUzf2lSiDl
PBY6OxyAZiOxDmQNJQr3efawW3Pon1AA6uAtF6bi3WFx7jqLjd3WpxFV2Lm9qhv8
2OIUMN3OPmZ7/sEpPDXdUYtD/vgT4p/R8He55LUxpt8u+3Rc3OucKCOfJhfg+0eC
fV9JryYypoaLUHgq8+2Hg8JSCnJJI1qNk9LcZk46W+I+2KlwIzr+pAk30QlPLQcD
v9vKVstzdepRU+7tFFEh9T7yUn1AAuzHWFw6HTFArpJLrgdw4o6TtjbGXt5dSCOq
w6TdO8DGK3i2znlpt+6DVWudLQCFhxuu0m14+JStQB77B1N8IXc2WPiT+t86lCdc
l+XmzX6jakjTcao8m4nZNn8vWoZ/IEogoh8V0OEeLL/ErUvsKEOIR34iRP0ImkHj
UIGR2t4Bh9H+1/k+A4UX027/Z/xd2VgRNllhV0PVfebbhczZjPrEFI610Osh0D6H
H3VPdUVdagonuMxds+y8opj4U3oGDOCHhIsLu+zA+HmUdjxn0DgEn+WKkCuU/Guv
Ne0tR4fH7kWTQUn5SWjdDsmFfOCtO7rpW34A3pK65TP6DSiz1ec92aLRhjxfp4Gu
pgvm872eL13892JLF0s0LjR3j5+ZrO9Z5dLasycL9eIphQ9fIc9bI6YKiibGx/qO
9sTa9StNQeq5ew+jjJywpXDuMiF3vmTzcY+YVkjCk3Ly60+sjFgb26EbgLQOwNA5
9jaafzuMRnzAkoUodT4axbq/YfiDJLHWPWK+FAz58rtQx2sfXEQXIsCwqrE+73rX
EmSXKc+xqNsMAyhbT0ao8F1JVOzKFxfS9rEZtBzAyxeG3P/+kIstqonvcZBdKTlf
k4Si2B/S8ZnEXCUj1TbakYSv2D74bKLNFon8exYopIVf/L3em2mriTZLooeOdIPJ
AQI62EvuWpOyd3qAheBcK9vlWp/qhtOhvNTz0/OFKP86QXRHwSfESxoXlMSUy3Su
8aH2eJdSkg+n8mvE6mmH3YltuPUjA23UwqDURQsmLsUqVYYywhOLl4o8+pGEu1d1
AoTgLIboTxkmTfO2upctTOKjawIaDSD6x4R0TZD8t7zLiZwVG3otKZVLjd9UhqMq
HyQj7yv9gla/A80TC62A/ZjSWskNxQ6RdjzXnUDPl+vKrhAzR9vx+Gn86eNIoYHt
EKn7Nsy9pWXWkx/BhmRfeh59v1e9Ae8oJ/Qxdvxq+QaBIe9TQpK5ngr2S1Ipywm/
gVSs+e5gvP7kad5eh6LczjXzsbP1tZARP/X/uC7FX1fjeiCSscZC3GsnUUxVcMSE
5G4Tac/Ji3jkv+MY81vjouwzCNoWYQBnM45zW7WR4olMlzxSRf/8eOoyORXtwVVf
YO7SGaGcnpAy1GPBT3rTP8gk43jsG8hTOCGQSMuASzTNeuS7cS1T4/USGXlWLnaz
02P+5js+DDxzLgrMfFnmoEzqDqsZ77jtv2oPTNAYBK9gNpLSG2CdNAqYYNDgtg1Y
NwjNbv6caSgC3MX5G3CIlPAI4IeMbIzvSJHDfyLjAmqCg8s6HKFRB7ccKflJusdB
PoJ+2oai3wvPt2ubjY/ux2m7dni3uJUR/FVDPSdmUH9ZsCds+//ztg7ujA0oAUjn
K16N5W4Jcx1rT43e2z/pCBZPsCjviG1rRrmOnT2TUXuAvYZ5p65Vq8v2ox2HhZb7
V1QyWab+MuTCihv85emyxx+0OK0l9dxAw4lYjlt0bIrMUo0U/fKU2RrZvwghYBCw
CzbIVEtUREl/Gknurta22/lLP6U92AizD8w+ShagElsZsApw1NdC8n2E8MzdJtbD
6lqtm5vtUQqThn5xgxC6d6P23d9lvAfRQYTDl3FmMXMtFTD3dAno4oC7SYzgIvln
X0840Q8DRQkXwShFyhR/f6V/c2lq83adtgveOwwNblFtuwLejQwi86/vWInagIUG
r6hjqyj2VR33/Xi1VofPgAp0TmzadeHJFNcO68X6LXnY3hbhTWkTBaWnRU9B2U5O
8R/gq709HzocdCa/Ee1n3ckj2cd0C9cVaAliAqSnlA3JuZ1FScAbaNkSyi/MuvKT
sAp+Mkqw6ZqshIVRs/Rd9wPr39DLT0pue/GCUSRDJb/kJGLZ15WF+hR6ON5r4wJq
u+cJVvVIhtyyHQMUKggbY+9Ok37U9CjF8ekve4kRsu9uIxQt3IHAfAscG8+afsir
aY+dIbOunBV4flutfAyJlvaL8pnnhzvzSa+58LiOJ9UN3BJP8Ja7Tb40O1NHZ/l/
EiOTESBXrIFMV8zTyQFV110Ski8QwNXFogBBIobujozMNLvvTMjbFFBrooX90C0v
S8pW+TbkeCP2x97Me+ovV+nh8qFakWU01JtGQJ0djq901bQKqufLW3+kczbv+EsH
ECh/yIxNx5gCOwm8eWiqhr8+61xZDpobkFjy55W/6XGlgRgLrX4v7Iuu7dcv94fl
mGH5PN0M5cPyLOUEUlJ1Sxs4c3BLbu2UP/hbZobni2XUHUgIEFyH5KTldV/u7jKU
yy4FPHHRQV33z3iKsYkrDWrPNW3vqKzqGnpMbhR3EgmaQq4+/OskT5n8Oi4RWHME
eaXMuybETPkB5jSb0otHvkej0Dx/envThGKkHGOtQThwTOGX8zMzZGlV0QDzJDI+
ADEfGRksptEkBuEQt4tCkflwJCit6vhXObq66qgeYUJpLWEMf/LyrTTsd5DWxUrq
Mcitw2vyisGBUP+ZQ/r8m+fZaBntJlAKCmQhb0aIQu9eapbf0Cb0ENgqaQh2ujLP
55r9vVfoVXVW2A+lj/3x3JAvFWO+Xet6F0Q11vJRMYM+nq9X/I5zlsjI8lFKiPId
onhGpyx3QVzlr211vHmYI9ezPcxeJFjQF/XW5ErQJt3ah4g1vMFw+pb/OqllCMgO
WTQB2RTNejT3GvFzI7E+nPCAqLvQa3u5ieVSIeqPLNktVq7r3TOvUAElSC8ssQ3B
16gPjE9PBTdh84pV027tdL1YM+ACzqXoW9rPlocFnPoIRNCsfmxn7bpNRwsZp4xO
slGAzG7xxUDCeaN2OJRetn83UsYveOBpeoFayda+xuGU4FnGf7V6JH2CNWJ8wbHs
NZB5HjybFZZ5rf+A5wALwzqdxJFs3QJ8bb6nneeI7wXxIpT8oK+jnY2ALddlDPgL
EsOUnBUZNVAFAYYnKsEjaru2hQpfwxuyd37E6B6c+KV1STl4CtzJH2tDwS1fLddy
9C5YUtKgWHzOZqyHTK9EAScvqnrMPvf7HdEOk5uxGZ7mr5+Whgyj0z2LICiteKQ9
brUv0M4u+kiU5OEQoWXq2wRZbVLkhTy03aW/nNRf4SY1kfUlVgZZmFTCLy5hIuNQ
iV3+mcGanAxvtn7s8ewFLUTLvEA29qhxF2olHfyVF8noiff7c3owbdbuu6pQPo7x
bPzMrJ+a5FL2ZO01MNXPOzCEkTDzhMtCSszkDnUbhkh8qLkFo4F+P8mXNl9acsUV
H5dF6vjSFFmH+Au3noBrrc/A/41bmAQzGNlER1RgE61lrAvmWjf/mLxNlGSNukEJ
IkdIkgwwWw72iwkXhD68xsn2dIcaPfor4boWXh+fVGfi9N2R1NFF5aG/rh2KCT3j
lSyXFhgfhrHjVXX+0KkFztkA6Ieqw1sFbdoQh6mhlWTck+HFBMFHETOg611/cWXK
SCaM7xnDWoMJTSbsvs6rJyFEkP3ceJOF5+3QY+bUZgdni2mlvSbCMOyWuAztK2oX
14sWDQTt6gojX2EoUX+jR74NqNUquE8WHpgfuBZ4jVrIQueqbKvoYsdbhkf2eemI
qcsM2SzUYzUTDeWJcbd/MdFKE9A2u5wuPa5QauTn26zK3dx6h6Uqy+If+0sUhpOt
4nJiQgfMpXv1Hp0BePvm9aXmTeEfGU6chUplH9Q+EU3tPanSGV6UqGnKAWtApYAu
N1zBKXoWEIaFlOB4DoGHg0x0mkkGTDpHXMtpGB4Y0vrQZBdoajv0pVNxIrq/ymWZ
LOVMOXwJpKbuaa07Tl+nYa/eUnz31Cn/naW6bFiRNnHHXJKj5sYU/Oo3W0GS8DlK
aEpwIATOUbmNQb6SpwE0fA2w4WqQCrk4mpC07/uhmMaEUz0+QRKGdJktIGAIfayk
XQ2AR8fdWBcf4VoFo+z8gECYftz5xrq/kXVOjHx36KMDdpDTtzP5GVHh5cZGmxKE
gNH8mLJNKZecYIlND7Gcq0N8e4ox9f1F47blcbvAMQHtcHcZFECZPF4R3rPKlIwV
pl656WtBK/8AhlcNH9RaaRG7S46k4ZM90Y0l/+K84oLPMtZ0wlN0OadMC9OWHzV3
7qm2/Ak67KW8AU3RgWLREvsg5lHPB86TPdJ/gHcw/FMOBJlyAPAax/2ObqrYc4uh
6oo6HEVh6U6ySlJJBVIKbOXRB1AZXbhLa/CMCMPfeYBcch0FjcEkCXQodffAdE4J
MKjxK35ivNmTaZWgGW+jHJHRQIviy647Rttujo4YKAbp91aS/tKNpn2pmfQj9Cs5
8U3v843nNMYktLnRFFdmYohhS6OOSeQqaw/3Z7fXps/Z8en/30an6w7baG5vGeu1
lviDaeJixF6zpjHB2bTPDs/vcMfF9ejgSUKfXAWNhWbxih6fyr69URWSuP1/nwXN
SFpcGmT4BXczB8VoI9skUAMWr6xFw3j+yyxs2+LLknWP208jz7NscipEESyZpPQt
Hahnvhm+QA3UoMheQD4bVNXZ+ogY7dwxdJU+nUepcPoCklMf4jweYzzgrLWA9mJa
6ZgIqSq4ut/uAF1tSeitFBz8iE69dJUv8g6VwPxchkDnMRh+vkOWfSjkn9kV1uiV
4lY8rndHUAGAD3V4yYrqUrVxStNTev6uEHPZjmDE6/mI4n2MyCx3ePXhaLE+PtoG
FAClKh1Fh2rznek0gbGqetI0TF7h45ulLQ9jVO0vX7MkE1ctUiwN3FeW7hqYhIOR
lOYbAhl3THaIdgRqRQndgxBIL6qieOu3ceQ/jVeg2MhEThALLPuI4ieK+b8lb8Ib
QWHULl8oQqGqlX74hpdr11Ose5WemTtuWb/P0f1MKeuMR8JkfYJcsdyFNhyZOwvQ
Y5WQNlxNHloEXSzDVlmeaZ5g61u0z1R1NQysCj7ZxzvCUvP46sT0gtYxwNCtvSVY
GqIWfEwlv15xqSPhk8D8Ne4T684Vm40/e6TxnQ2J7KkQ+4cyRlGhiUYAZ4JQ6oyh
iLEd7gru981a8U8PcAIRYV6UVzLqhpM6IpBl4n47MoiYynqV8mVSbCF52iPcaUG/
/OgRZn1eBu64hfFdNDcWgPZPbo0EjcIlLaHlQEhtKuWEQdU0YcPNRwRqSBvLVmiY
/flSDv/x5UsUAx3VBDu7gEoQXEPaMZKg22XBklr38Q4d/uXtdMjN1kdleqKB1LIb
6+2P4zYqb7ap1TjfviPNjGkotJVi/4Uk0XdV7oBKb3zfwsmVjDE7u05Zo3aHdM2v
Ac3bX23gsaXvLHB+NmRpW6sAXTgb50tq9RN9O3N/BEC8H3UTKM/gJOP9vOmoDILd
cfQe7InXcqoPMNmblle4dBq0D8m6WjR8/+edDDGnyHTEcVSqXfC4zBDNWuSoN3nP
Di58IPQDdxyGPhVCxlEBfu9noSLQCuSkPtpCrpPFOIH0vPghGVS5HMRTZ4bWA7tc
fO2FQ1wHiMecJoo6DhSmzPxWFhTTUgQzd2G+5Y+4ZBzDfljZnLIo68+mDtMAK0ai
9/yXeJpIRN4VH7YsccM2ceIB5Gh/+mY1v2EVdXq6PafSvsHSnxmXD/1crntRyhky
FvLj1hwasldFNyA1vCY/ydbu61dPIR1nhxsHfxOOHnzblrHCXFAhRyyKjUppIzcQ
flqwJ2ElvtlZehGFc/mmP7WkJE9Aw99K2sMWCpf0sWGauPWO3vGo9qUxzFVISd/N
7W5wrKJun1CW/nXUkXaitvYXu2EkVOervcR58PXgaEp0333F1FhQ6tUw7r62w0PN
n4VwcPiGrOg4ecnFOqjI/nafxcZyjNlsgCyCasniFRr1/LB4gcK5GQq2t5FOMpRR
2+qcWRhgpZGmxY38fZTxnSM8phw2lcZVhCwzOhJXuqAvngb7owPhmkL26sQHxjDa
NkLLxMTlIltprC7DA+ugDLRwACwizkttwpkipkX2UDhHQ4wJFkruIw0UO6cy4I2G
g84rDdkgxyx52Bt0L3pEsiZlSWzGYqjfhkeNzhvHBtttvJB+zCoojvUmKdZQTglT
3zA4Ws0z25QaWhO0W9X7pVBnpKNjx8HM6hlbPy9/G5pzBgh/D9kibMBqhC7GFqzf
SmiYEA6WPXaJKavLDgd9psaHCagQCwHKg7bvS2D9aVQRp4dgMPEmcbixJQuZObbR
IAB4vDPhLUDG77m2GeJ967Z3QMvvh18ZWTCWa3FSg01FFF2udi1pD8MrhLUJx0C4
/cAqTV1fD5Vd+dhrcOv0K1tzPYF3bS0bHvhGMPq7CNxdE01trRHQGTD3Tf9UHnL1
twpzBneGdTUDWCfk4OkOcDwJNjhUEssOQjncBUWdWokcSod3mzvpJeKLbhyy7qZL
hD4ABYegrpZA7Mgr8Ih2HLTjaVhzqINHK7TFTKgmTiPDHOIV7AExaO8Klgk1kf58
1+DVVMy+RMdW25CcXxPOvH6LcHP1BLpDOJ2/UaeemwbzrD4Al+/RMNnraDGmfQd2
WRUnNK9gb0XgLFWb0rLD1NKITfJ6FFmX8SybYjNyLGGNbY+KWd2tMEAORkPKr+Sl
AvWogyvCDNCZ82YW3reyCmA2kO3Bs1iiCLi/0oAzIAG+tni/PNl/Jr819MwxkvFw
mCcNeLTwbIe2Hb62R9wzDpgSiGHiCUfRbBeS7VpjwaxigOHhCOAMjiSsdvCta1rx
hO1mU4q+4zYZQ7f1mwzo2Q5DLNm9FYyf1zWcraYaULo+Cbf8Y6uh6YdmR2FTDDCK
ayiObzUqtfbiZBjjmw9r3H+HYsZH0q0PLbH72AQncFjQqSQgjJB9bLOT3UK2b/lk
lCCoKtetGKTdET/X0csyAYjDuo2F66Eeqp9/VQcFjog4ASjp6YzWiNJf0fbsKi8N
R9xEALTokDHfTYK5G9T6GoECIiajERNBdYKp0U6EWWmMUWIa7LSK+lti05ppSDP3
MZ4YdaD6cccBL799R3Nk0YxIEts/JMxONWAMr9OAiJEOYLUFLxEbrdGbKNKGjgr3
2JC0uXzJqrW61xVzmKSw2w==
`protect end_protected