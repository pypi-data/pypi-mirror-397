`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzY2+EFIYXUoRGNXzJ9ubqwb2XbFmENkDbJziflfXpluz
1VW788YG5KtXQNj7uMGO/YBC5cDOsDs8r94RnpjRLy2B8ync2lV93Hh43x1JP/9x
E11N2o2VumeOMrJiAT5l/HrY1mdvnnmFs4YDImPu6H5/Sq3k/n2WqxDsD4TNJyIV
KOzGTzwUrSCUTHfi2XzULORNHhlmvxPeP9FR2T8Zl6Uc7LObRusPSFEuFdX099yR
rVnkrpVu5wLpi9xY+Ac/LcPIreYiOErW+zTT9kWhJNHYpqqFUSh9fZlmYimWxIse
6CMX5KMmypC5g52+wDNVrIWXIz9vGQwQRTj0RVHulGxjmC+cDFHyv0SywP1EGcTk
GCBoaHR4AKY4nUa1fXmbw+Uv8Mtx02sfxk8rSaEcvyTPzPHrPdfelW0Oicp5St1B
cI/gmW4SBsO4b6OAfyBo0H9Ly51MaX1tGLNoz7tY8QmWZjGlpq4rR3cqzSa11mgf
eR3RSxiAvXRQmAbanaT/FwkXIHdrCdrdCjSbOA4oFDMxc3gRyb+IZPLfQIAH10I2
ZI+V6YMXZxr9419P6lMtYVq5bZJllgeh+GegGUWiepoxB+rMC9LxhSmA1hQCGJoU
MjVzwEksBoVx+Y8MqYQVCOOb01w6eIxRZTeYhyRJgIpJo92UBQYNRdt7Q0GmwIG1
gQQKb0UdxiJp0WjqykrIQ0rGQL5sxmYmyaRreoCfJl7cuECJpVy+mIw9K196k+dL
97LctJJPsssMxMcmS/ZWfua6kEIqjRvF/pG8CQoR9SjfO7I/9noRQSrEMo6K2yk3
nc7Bj+rW1nPIbyWFExYv/rO1/Lr7KBKSlON+Y0h+kC2GaQpiaS0OgHeskcOH5u0D
F9g05KPFjek4ORM2/KqLv/XuiOOXGrHuE3t6gku2N9V4MscwwtgIes1d6HSs0hh3
HqNE33Sk3oci+bhWXGG9Wb3CbU3VPytPUz59EUSvmO3hGgSqjCuUZFItOwRZQJgy
GEnN5JMD+u5tk7De0ssvR/EZToBsF3p72cgmboi+JzaRZf9A42vx9KmnYMIZ6qjX
Unn3P2/WizsgM14FU2kUTK70UNQs8uuY3ktiVmvbjuA/pKI7gjpTVTDFNh8NhcCM
j9+gUZfos99yzlQENRWEZ1HkvWGH+2JEQnIbucqC3qQAudxCmn6XO10qKuWeWROE
rGkl1zAJCG4XXB3VYDmCrNsTOPoocXPvageet/1OtO1lmmS+VEwCNebX9x9v/XhU
oCCNYVxTrt0xlktlaNfCE1N8adF16O6CCHBJleB36nFNKgKP+v0m4X5nS6ebiO5u
nUKaWKHf68oFuUrbEbpJbOXhBSJsN+U2DFumCE1pI0Xc7XgXyeExpJKhBOE+4v4W
0N/uopxOHt+IGvuNmtGqIRWtd3c5QMOjFduu1R4dMzXyj6s5FsmUb0H4OUcLWKxk
q1d8b6NJ+jHc9T4TSGoWrHT85xVbBR+Guc/8Dt8OMnkr8GnDQydMN/gVoBRVFQjv
kr9bquoPWrmSJcg4J1DOM2YLhBwC5uyyOC3j6u158CP+XVUyg8v6kBDH6kFwH4F9
hj3YHas+XxJolpWM6fBZtcycJbdeY0vpCfodZ8RTS/Z0C9N/gyA9+kCUIGZFI3Ro
aLmkdcGCosr4p6QOcXDnZPTBSCBTz7yWxWiU5szvhR+uhW17mEZeLnfJk4RMhEXw
p4MbU3MV4k5YUeiYTJ4lGYrwFHAxDU4L37KtL5t9zqXeo3nTTVdhgUSplwYtXwkJ
On4xFDAyPRQZzGeuALIVXzB4/PSUM0fA+z50fZ0SmUet/zEDMHalTn8qsDQQviyt
ofJCawWlCYaFaQG837SxhknfUZGvIo6PxqwQHVij0C+OLXTIS2CGjipA73QFPx6C
LjECqmz9SSnv3oQLSKVfl0RTygtsv8zOmwhDGJb6Y4HgJcHByjmAtjE541b4SKf5
qmmwKhdKulwv8Uzhjxr6qOfHX1B1fJVfEw/uK4TLgY5tqCnl66Zpq74rlWeSun43
4zD1e6mDQgQcyP7eutWNgZnYGye79IvHv3nrCSubwbM7xGJsPiIvry5Jj22lEzOs
asA6G0BDpVcKL+3HN9EoqM0l5YMul27n7E6ghUuArpGZ7obKwEAulzthEPkj0so6
2A9/K1E9TIcnu+rxDBSuYME0FqHfnk5dfaiL/o1hd09y5XgoMCP9ex3y4lht1rDW
lZDdPewEUREslMsUm72TDJGCs9KJAxVJv5BUhZpn8X8eFtnH91ab14EwUpz9QIHb
s5EvRZrfEU+l+jjEPe0SWNU1/ztGgr62t/3/vivEf8GmcqTEM5BzSVs634ImiKb+
Kq4pUiioSVDDP0AeYmFnWo+Bfpak9B/IYc1CR0HtNdKqBp8RDuOsdDMO640iPe+h
9mV3+Rgb7eC2SkdY5UWIVxov4HgPaxXYe/w7/D/PmMfwKsS4VXleR1vZPRHtK2NA
6UA4qzB64Kd0R2wnIKMp5yaEl5YQYy+GEBzqB0p3tx9VUGrMUBiYPp3hdObDyGzT
IOIE5isnSAdqQQW4IQagZtTO9INuIke2cLwmxhZ9dOEmLflUDcMQ2IQyheyabgsO
FoRI0qwXUJ/7DBw/0o/hozumlBps+02NPlEMe1id/M8ICtHYVlIzq1XZukHfqLn4
l3adYitb/1egq5MixX5tcRbCHX0lNlAxuqeFyG1aoV1CQ1M57Ds0YZcNyJa2/63f
ePjDb3zLIcM9YjijqOP5JJidDLNTOz8cdeXQEkRar3bwIZEffp4hGsabKYuytq61
nb6HR7Azbi0/qx62JJUaJbNaa/fq5O20uWS0rOxgULJ3ffhV2wlZmqBcmliq+Vyk
27ImxgUw221BovvBcrhjCEHgG2fCqllAJZn9zA3sDiUGYdj/952OaqILH3kzYko0
6nAhACMZXCiBKujSmQs8vr+xv/oxdyE/5gsF+HlDCiO1NYZQY+CYJOTQFgODgi+0
DowdKcsU7vhYb8LEYunmskLpqolj0ysHFlKEzLVcINkodqH4JUwLcHWMpgzhsN3x
LoKE8SwVgXXTM9hVphPCvaIR7oHf5FcHCMmUz/UWjJ+8PKid4R3cKMDdYcDkDVYz
QRbgOJgLgO0NyLq+KjKOIlfsq197aRLiLZbhlwQx5Vfho+L3Ae+byYyP4S9qorvR
HcNmZ1O+2dLNJVqmcEzf5NZKO0AQyj/5WULPY+2hAq8DgenlyyId4pCQqsXiSiMh
UrbjRlCMp+2GYWkyUvTyl22aM3ZLZfDqKJwu2PCxYlG0GXgsizoKfYbOrIzEIxUY
SSLiJ5HG1QRHS+JMqwALJNBOhYMwLlr5FWUNNcrTd8qiFSi7WICvuh4RGCXze5Uk
l1NcgFkUMbwkyFuIYwFuvJw32BGsj/ZeGfXUq4Tscqun0kz3lLswfZyWH07NA7LR
4PICZi/KKl2HmYFbFWufaF0nvFmyDZgbhTKBgtCmSb80X4yU0HN9jFkLfjn47lh5
VzDQ+8IDWNHXay+fwUMxx36vc/tS2wS/lpYxwOfyb4oGPatCglWP23wgUH7XGtZ/
rMMXRU7leRJXcO4Yz8TfuzGbUDEBNsgBoPIZ2j1hIQfp0y2H+Cc+X5mnuobgEAsm
cmPKhqjkXTXbcFHcUMzzTJ0nuYGWVE1JXZiY/SfBvt3VoBeAqMvOSk7EBe9LYNO1
2pvG/Sot3kKn45qtVm1tvBv8dWuBR1vnle9G8Mx0CS4fZ7KgPCTwUklTi+yj8A6E
z/ZlQlDioUeA6iC2JaUoatVKPbbS6e8oZbRbLDKOao/Wn4m/X75oEWFEIsRPIi3Q
Vb/HoivMNz/F032kkQPJXEgrd6ga5Rfj8gFQmE8JNXz9amrqU1I591Mc1u0eiNUe
H1EFqh56yRp4zhOA2fOjSv5z3PxDkBJlL2AFmqJJgKLSufCI0KE/sLsU+8QBX9Lk
3OwtyNnZRd9Xf//f3jHs/rSn40Bzolj4pXL8tnuspADLwKGOgrJTlaO3+iNzrPoH
ALvgiYsuv/0asOLmOvOdZ0h0TUDgKXWagngbCqp+ZnLMU2lt+8xJoK85+3cNh1Vk
YnSTytqo/2hUjHbmfqWnX4ljXkAhNAO8UYSH/g2/D08DRdwJFEe/9Ov05Bz1DFl9
g9aFyEvJCyM1pe8p3MnaliAoFqcnXbtL/FrtFRE0wS6q1AVFjqnggWE/8/9Bhqp6
ka7q/DR1p3Lwgr7es+XWzy2h39oec6ZOYsxsAYCeuMhqdxJivbDduiWKrNd6BUhb
EEli8TQdXeIShZWbQ+b6ZiL0HBvRFHd3GD8SYBNrsXuMoWpjM00g6dO9UbS4WWka
4lYAE7ML1Paf3xcGG7gY5FIFG0Dxnri2zQcrEpGk2vXSJp/x4W3/xFRggu98oh5d
8OyZ8c93X1Prxgz6whdMTgIL6OlNst5P5xHzqrsdIeACbEr29evzxOueBLvBhF80
xXQrtI9E03vh5PTsU2EvP+2+empSRchL9rttcfnMa84fFQmxALPTn8MdohOhnr/L
yTz5km40oyNeqJQIE/00muehpGTUa6MqOWvGdLCgG/03QeunDD5NQ4lTl5KoKVNt
CSKMG9k9Ir3Cldj8McIgIubj45JXxEq82BeklrluWVD+UlMft9QsKCBH7DBEo8OF
cD8Lrh3eBlxH3DYJ8klrDYfgPWMsYR30vOQDCy11uzhoTrrBukdL4irfQSSZuRSi
4D+3i9JDo2norNV2grBtbe1OOxYMk0yVttwNZvxIQES+Y2ZgsZeHTR7rX5CmH4jU
ZGF0JqPOqoqoifl+kbQRgkJRdz8/VaHFug4+tB91qP76qmSLabsHYa5BhcLSdD51
eQpBkU7qWMhckGGjQFCXCZBfALmZkUqb9KCqgsOvSSOVeX5SSRdPQz3lhXKzB0oG
gJadqQXaMGo+0q+IOZBKNxYF4UolY2g2CWmR7rZvMRNyQoLeawYc+FeiC2W0Wm2K
3c0uFWrgoWfoW2tK8M1Ly2pzPS8FYuKhb7RS0xjr8tbZSsDu9mkNh1p7al3UIKq2
fvnSWe8Ts78B5/gLuyrHnj//DvJdAoy7zn+2sqic5PTutsoidfXXkx7eHqW3ms8b
3c5zXnkBIX3rnxVDAylKX0gbCg1cDkUOEE32orlSTQJRWgJuo0dgNAJCScIUAxvu
yQjg3PLrJRcf7NBTy8Es6iHkwkg2MIuSw6LX0UdEifMcg90/PWTnGA37l4C7N3L0
0LZwxC2IhhBc72y9OnBNMYBd7FWo+iriZXGAtecG/TKdWcj5/WpKVJF3Tb24RIxl
wlDTM5Fjo2fuTUhzOYMwsnOAaEaZ3MduUQVE2cmgyt9zAmvr0ylkWZikLiS6tH6P
nYIzKCVFnia8KWJvB/ju1SFrrM8So9pOYJVLg40nXmBLIOHiPdDKtfvMVR+Ub5mi
zI8X1SS7MiaJKl7n1L6OIVxNba9uj89C/mwnhZ94E5sOjbXWLU4oT9ogtyldMWce
TAjW/4bq0R3B0uHXVhbyg0WoX21OY1o3OVobyXrzeD3bQ/oET2z1xEMEC0Zd+gz+
7+NPxNhDLW1/kVlN3YthhbH+bmNAZNYlIM3H8sG7QGxpHs4sk/H8sC+MTjKpOfvp
7F01UWsEv1/OgtAFDHHpXPsi0f7g7jqPSOtXlD7WXBTX73B8RMg440aFc2cEFDb8
nxqULe9HeveeES6II9n4Ubfsn11hgRMcOzv52C78/lkGeXKgKPIks1bhqvRaeYW7
ouROTkGxUMcpapjYsopmgmWhKv+OUXK6X/P+fI+BYEbKKggC2z6FYw9Lv8wvsX6k
pqVRll1tn0iw/H6HQzd4zabW5H1RQWtAzU/Uf7iAI46WAypWwzs4warnYSqFueTD
DhQDHCmiJfsb1h+M7QJlIIoeljZIs26VT8qHb4/R/pFIjJrCv/tJg2guaAde9zL8
K3o2fcdGXZednQoGtu48hRLhBGYRnthuIKH5FphCLZBKXSZN9z2/3hE+HvEbw45t
xNkUmTjgFViaMw6Trx8rWC8mJj+QLa+ZqDC7E+oJMimMPFXh/CIcTrJgVV8y/iCq
TwthPwLHxYEgXnIArgn/oeuPeE87qmzinHzqC+8BKkQXXqxVkueWg7fa4qEqRPlT
ihQ2I85XdNQWdpNLbw8lvMgqjnCLfhgozqDGtczewjj0OSiEXQr0PUZCgeEaY3Rn
AbIWmxsnXaMR54Zejs17WnrwKqsNHIlUIRLkF8kb+gRDIjYfYLYioTvxpflfGJiL
7q554AI+Jk19eD+zs4T7SKk0DxCicLRFMED+tvhYKpiLNjEcXHNyPwa6ymkM94M9
9svqXp9yLsFSVne0eB4TfW/0HOtIrSNsHgQEzYv8lPQbRAbROmX6kcmkZAD76r8L
ohQfUZiIkReIYmSsdACuaXknJJC7kiEdLvdJO7sadZobpAYZ5HXg2AcRnZFAe1Lp
plF4aAnZdIl36Y1MLhztx6MtmBoQcJSZwV3i65jGzN7JnnfC5G95BYlBpfEVtpxd
r/R/wEzlsUtfcWxXOV43BkJPVrORmjnyjtKX7WMEC0E2QT3nn2vFJSeip85+sxaX
ck5saJJp0BK0dKSCN2TcTQn2/jO2QBnfld//A60INtxzya+J2JxkarQ3l8DEbHqi
sp54Ep8OBzhmtWIPsbIO56dWBniU4rgetueU2K/MvvZjD0SH/IRWLUzuyw6DwINp
u6Wg1fQG8NZ+9wsI9DJw0r28YAwdAiEKdv/M98vlg3DsptJvn8Cd8GUmhgaWNx2c
xfOt8KQ+wM6XqSEzipqFxL/XGygbVW7dwzsYAPHuj9DJs9DeAQtMSzAWaL4oP1d7
ypFr1mijWFbeFlUVlX2+f1AK18Gdiu5q6IKhNP0PbKC3AI/MS3c1bftlFEHQohx2
PGp/D8XnsBGhQz3Bb9284UCGP63LGeqEaHHud6RYVR0jFOA+iJcn0QaOkvPuFzjV
xUCtvb4Yw2dhhjXRWFKQX890dnT04LJ3DXdEOFPWuqaWNv9oi+LdVnQOLLBniUYN
+C6C6iForLjISTjNx87S7hJqTU5AasvkdzeMQ+zzFQ94C3ihTyIcnDl52/krEXN/
Nzzy3jNiFmylVVJWV4SUPht9HNwyTuChnbYs6wCf4hp9nYtAU9NhbxQZfEI5UKGg
mdrBRG+6/iQn4ClPGnIlBQMPsBbgSI2QkcAZEN+jvKqD3rDuT0oS0oJyIK0x9UF8
D/WgHZBatfkiJCiplC9KBdPxxdrcRa8OlkMh5F4QrKdQbRRW2C2ejHUhp0tlEDrt
FJyA/E89gpGZDtfAILZPgzWeWyJ5PrgL65koSvQxINy14TjgEAu4inaYXnmPql2q
8BVhDmr55wsb9G7b0c6ADVA+iPsSDqIEnLRje7a8Ve4esMfugG//4EEtkx1YDG/b
UWHJ4rGWLrrF2q5uEbYwkh778qCoY9bw6vm7H8UY+X3rBwzvvQbxhSs8UUAc5ZM1
EjuDNwIe/psDrTRkbSy9lkND7FMMlLHT3k3VDDL7HIV/DntQ7BVktp+TvKIZ/nRK
JBpvywJnH2Iivi+OsTO/3gsPWSp35zIyPETftc+L9AvGpyRaQYGbEl1br797MMOE
/wrp83A/t2+JP4V4cUchg913tvlof8+RgfCYYLqvWhf2N3tzFCdvyFNWSEO7Fyvx
F5t887LvwVSxdJ2/7PXtJSSAW6Y/0mVqD+Nr9wwpeHdKyV80Tpi6Yga5BxXUpo5T
J9JRZgxQsi40ImVZnicDN0n5XH2zSERp7y/KJimPGK56yG1wHBc27GEMwQumQGG9
fOLMVpGo12hN+dUdWq4jxpg7hSV4ZiomQjpZDies2mkeVqp1zRlltO4ObFVms09T
qTyRQo2P7etn1jO4+FPE1PhbKBXwdsl+lk16hwu8B47yWhZAHwee+rWzuHceoDZf
9YPcaAYUE7S0LepR45YJNWajlqG8UkQiMM+gaAEQWrH2vnrWtlVzQJU/gyqFgH4j
hWeHGSBoyZPyzfHtFPBX7/j0McbeB6pNBfwp9IIa4uFjqYrQG80nLd08aTKY5r+e
qcKbJ9KZL0nhnvOKb2/p5/Qesi49F9jsY1+SS9wV0llrJvJ1l5xU1hhVpetIcsCe
E1K/m6zWCsab0uN0DquswgG1iqxxhNR53Y+0Sp9UWxnDhDACLg/cd6OngCxjL4ge
mRjl7gHxKwLYDEGN90hTBaJ59XK0gDXLjsgw+WP9YVyCdFuY8lokE9TJ8BauTWi2
hbmWy63m4AN6v31CD10wiemzZAdRGse+W8XOrKuKbwrJ8OVfn2j1ELQK/eF+IXwP
yvmKuYkusFdbpCMFad+wuKGDbmv3b66UPC/UEMXwK4Q4jdRkW/DLtgL3Jcb4dQLM
AqQ7eZrk6AoEtjhADDe/fGRU/IQJ+mFdbogoLZsw4Qokh8e56zuP4RV5H9RvUrkF
y4tghFXE1gyH3YrlZ3FZxvnrZQ79h2HEipp723tDwW3Rhn0wODvulycCaf9tY5FK
uxlV72gS9Sde+D2YAp6t2NVG4spqK6J0wQRVU1tzY978Jn5nV2UK1a1WLslP5KRo
fx8KQRiaQYqMUZKHkXwUPgmoVG23b0pCz7uoXIkDdhYQFVE/nWnyqCdYVkvK+YG1
LwrLaos4FOF5WFZSTyUMumKuDfip2L/8aktjeHRZHfIpkJShoE8cP782HvdUpVmf
EHbIIMiEhoWs4uWQ84IYg5upBJF+WWa6zYYTaq8yaNVsm847FwpuqvLamMCIjiAz
TQO8SUPnkuYZuqwtsZzaGPttVLSc51gowIWXWtNJBlGT+Rc0EBgz/9SAgEGhuIkx
enQTKfHXPrZkXK2pzrQfXA/1ciyi59r9dGKTfMgCTQ+KZupOsfqgEYJ7mKY9X76U
hbRz57ZaMyJXdhmu/hR+SYv4rMJjJZxC1VHpC1OiQyFwJ2Ntfw9ld9WbARCEvggW
DLKdVDoiTr+zqjFzKzr5lHywmNZ5MGH8nfa5wY6Wk9vu8PbhSlq2yHLbgTxgq9aI
m8st5uNJAv1sxBYLPH8vkU49pVbj9YHF+uO4XFi3nVNmPzijFbhgZaNeyjhZRL4J
6jIUUkQZ6glTNHzgIAjh4U3kOwYCgaZul2TSAOiYf1rvaP7mDrR/4WeKtdD5OzZe
tqov9+Y8PG9nWZxYbvkHXGixrXzwhmT2Fb+2/FVvNIySff6zc4Vd18S6otfApD5H
zcEKTmrhjD/7CKOksvE0TAT1WjbHq0tIkJ+UnTXUE8tHaza9EQ1Met4Up9dJW2/5
5/Yn4rt/lOOtGQHoO3n7inTIK13HViOb1++4iaukEyoK6AgU4l1uQwr1ZUvAg55Q
OtCL3yVuldambm20O5eyHj4jSOgzb6+ZhvYrqxXWcD9RzJ7gL93lU1dKeYQp6bZ8
ZfXMVIFfHfe2QlAREB7KMN9a1G1bhdlfa1sLLyguMmp4szZ+yQjCbtIObfofRy79
ICIBdJcioWI+b9gDZuDxhc89+Fadu/ErppkTsezn7grHresYDavQ2BiZFPpoM51U
0H2Awe15/gbsod1UAzsZiHQL7iZMaICRcRhWfKFnj8+8Y55dRYz75/517oz0KcDT
5G8wGFbmZb1EnNWLTXt6Mgh/YMaN90JYjexXNmJgSy4SYww1FZcsu6zFwpt6ljW9
BS7ID54IG7dHJJhHFQbEaLExFTkryMwfh1gozSouegO8BpOfe64dJYuWxrqdrPQj
Eky95oR/Gk/NkMBSL4P746c5cfiCTUP1ABAA5lUv/n8KEQTfbQhjxFhGIP8rzs8u
qrq3IPwyCK7u4qA0tZ8Qj0/aE316gfoLXuz07d9i2g5WV+cWmR19fQkPzcstSRIw
N2EKUv7dU4tdnkzMhLH5ZuNM5CaV1Pa7wuSCR8Kqm+MU6TpnnwJzX1ZFLVXt14xq
pTt3RQCe4eM7lmjtiRlqZ4OeZghYvAlODJ/K/mezRwsVdiPgbRkBjMAXDq1wyLcU
WAg62SRBVsIab1BhxgT40oWJBX5dmmskPuGhejHOelKxwal8Mx87dp1qHxvST8OP
ZoxQemDJKqdrHRKVq+CTexMiSZPFPwz0/8ZBgyluJxJc0VATs16t9xHDpARXjUhY
cYfe9/NPlXEJGD4Kc8mS+DOBCvR4YpeJWH1+V2S7EUInc2jc2KKsGDuMHE3SRCxS
7mBPShSjW5TJp3+YmwKmc7AdZVteawe/+rkTXhPvgt0aRIXs9GcD1hR/lFVkzfuH
sX5R9v8TDziM04O5SZAeciZKSeiILxPadND+wOX1vHioJgSzmRmp9ZDcmWuBMo0Q
sjqH3CihyYoTpVpE4c7Al1kNGIFT542ReQzfc40MMSkT4SvI6LTu5RW2cAHtE9NA
3Raqy2bqscDxW4Ux33QI0KRjbDkFqkVb+7hABFDDo5+Bn+8IASRrGBicXoKv+pJ9
Ie1eaJ7yIWwNU4WDcViKWXFwiknv20lWhI1JjLnfzSzA86nGsVlJCLlZcle1udLn
V1FBNLT8MQzQT0jJuXMl2BSDJjAjI7+Hgqr2ozRx2WT44hlG7kEjPiUQuEZ6FZHf
nXtSp9CXvyHTCBXp8Mf5dOL2/d2Hjvcd+2w/HyFkW/sQixM/bbRgZLEX/vIzt6oG
/SySZi7j03gxBQUdWX5mv2RNrz7fKN/tuUTz2ugNZ3qZAqZqF7OZKbhwVVhaeaqn
b+w+ak1qwO/0uKdicRBgYaIRD94laHL5yBH4RZ3fHoKOOWhR5QBalPrcdTRbuxJu
u5qZZJSK5EuDtnN3UPGW/038+VdgtrNE7LKb03rS97P+s2iCLr87ifVtcWTRba4a
jwVPVe8YAvDZn2apDlNgU9kEhDeNC79arIivLjGxvfSI9RYXcaDriAqyxvZ9sJAu
ItOrereWT/r1dVbF9Gf7RKPC2QLTOs2L7fu31WBCozEU55BLxHiuf3Q10rWf/HDb
zgoKwp7QAHf5ETm/z0qJlxyF4xIaKqETQfzsDMaebVycBwEZ1venU6avUUB9epFK
/xMHjYj385Ff2Zto/MqeAOPmW/VOxAW+nCw8xtN+mmQfgxoRl3xV+F12KP99cKmg
I2glNkBuDaDBQ/7W4gFqP67O5kQ78CiWLxsGIaibzKDcTH1R/dK0oIVntAH7+d7N
t/Z9Q/NjW1J6XXXs8HV50KRZVYyWoLpNsd6DznWRYZL/MKoBo8WrpA70OXTuFUU1
2jGUzw51oQEYQjtdC5nNoNQ9e+DQd3X24iKk0wYVLiJraWMl63hg0PfcqSq9pTBp
Zz+obI7zCtOGRSeY+AkPdh1u7ohWEg23piWW8nzXB4k28p8f1UWLaY73NWxl1z3v
EvF/n/Mi1ptInSclT8T+OG+fdPApG6Jd83A6RD1mNrIVEz9jGh+HddLV6lDRt9o2
BmTOL0x2Gbj7ssOKu1N6xTfxh3ubGYNA1q87nv2fp5vUy/xku3fZWIxDLNTPYOsb
tKinqBKTp1RZzCGPSF0teCDSg8wvU3Dv2eBD28YuDz5H5W/zfFSI2IECnFlbVC0K
4XVPhvYWsjyf5GhYQQKtL8K+jUlXJ7LDSlhsQpP11uspvAUfOMJAKndHijTbGScO
w4jOVLdOhQq6UR5KwCmlTQ4GRUpbkSHZU8D304Dw1FLs7JGbL0GOYrxRWO8jlajy
3qbDY8ZnOPf8SVRKTkgvv4suvgafhjZGPAAnVxdhvOq5/whK2qxZVlfkTkSKSLZT
++nKuyn71eUKolCiELn402Yp49Mj4j+FFlEpuU/EeULE7t9gRe7QpmXfYe8FWNNZ
4IRYvxrKngWxDO23fe1yLzAJDH1KtCUP569BHEyuCWas/UNfDsr/Oe4qe/goEzAX
KoaHIPW9WpToV5fVo1kbOTgnRkeJ06YdyrGiy46NulNJU2MayzPKPMk7RKUpcoSr
uwBsC7wgvbbxg4FoKsqYu0qtRBqVhJr21xq8aXnCC2Fi8BOs5/iXd5Hyu+Y6er7X
omTRt1cSLn+AWod/yXs6zH6GNxx+0UcJH8cAwAcXtzYobfY5PxBUd7x2ybCIpFbB
iz8fZvmZJq4g/6VPjhjyVzq2rB9POsNieY2VE+35k/w/5MJ30wLmoQMc9zCk1UZm
Y0qcfzvZY/F+PZQ1B6o/k1MmiCcPTHHAqWP4ZUFQGbt/1DMqx7DK4ZrNmdIEyoTu
0yEeoaNeq8ASeOqFY6dLlg/vmgvNenqQp7j7UWNwfqMYMvzgqZrwrcbDbk7/YU5A
8TQsH4mlO7dGi8MlxrJuDgV8OS7ZSGTCM8OWqNKr9UKDxoWs6rU+uYHnMiTk54kW
KfJp7D4mjUWp3g0IASEj+Cvj1q1xn9Z/ZT1cVoIB16CGU0FSSvn3lehyc+KHM/eQ
jwjdrgIJgrx840oIP8/xNK9/jhlEoL+MU7XJa5bXtq/IeR6apcadAnFl907uVLhJ
b5ywW0G2Znih4a82RIUAhp0mj7l387MA89/4t8lyle+qbRrrT/l72QOUwFAq3/yk
nwuc6k12JFiuJ1pK+taEH8bNwGWyG82utZ82Rst2SfcdCf2BBn4KLEIlXLQtNQFI
lWXrBteyxGrm8JwHe+MeAS1+X8y6mEH0HJHSix0w9pKTuZ8L3ODcSY+EjlunmtKf
flTSV1Ckm6OU7xxqhZOiBAvDI7DtiScTPJAnU9DDQ6mSy0GEgMcsVAfUXxivHlz4
KvunuuCelrBC7ppoILupaRhNweSATrzseOmSLgBNwIRPLYzZ9dY/mkxRhjX/IXoe
L4kX5RMcGiq9AT5UO2EVdDOcB9YMEiduR+Q1fo6W+Ay09rQPxpA7ELmHHql4jbG9
c1MqWppbWWSssX6uEJDqtp4YrElKnTCLDzBLArlvsV66fTietFwLsSBtkKuVIlm9
ZYPKrNgdCADf2ap/H966EJuo52zlF1CBqJA7pS4MwZUExfTdRA0Mul/w1OpPAx37
GRlbE+JM247MPyWkbXs+pUrX7lzqg63r2LUrX03jKJvdjq0GV1DOvDEJmip+HaoR
u0Q/Mc2HX7cMs8dTe83+T8nuFny5liQAsev+a8+PlC4gRN1PtMnSqQe2LmaW4gDo
n2rPlhPmxoWCUr46cVpCecAX7mx8lJZtTUyQ6Ms1wZjCHsjcVxHEVePXSNbNqqTQ
vuVsmRwM8ynazV3fK7LCuCphgr+W2sVctthD59DjdUXvXiLZgujvhMiwtTGomkJC
jIxQSXtXkHzsqoA0eANQndqW4f9QHiP3agZnOnZz6jEQYmuYp+mFSgfBi8MI5XoM
16DEQzR35ZiMVY5+rTNvKHuwDNkdSGC2nlrnL6XkmzRdRecb1yS4+0lVqhnT46Pz
jz0sgmNeXpuqgTgolOYLPcPuRDfW1Ja3a+MKy8Eb1r1HsYwuvYvL+NnX/uH8+iB+
W+97ilu9EhxMJWifted4xVxUR8QTKU5R4zqbBtJ6GdHZ6mSSRVXSMmWFK/rj7hUM
BccTOAJgc9iXA9NC9DOANohj44apqnybXABB3aBkpcUTx6+wn1Iam+Fw9hYTBUYP
CRM/GQzqxE5mIq4aWDtlzy8usvw+3Hh/tgO4ViwAn0An+zrBF9T9/FG5ziOXZ+Sb
hyOk0c9Bt3UCZNP23TBXb7+rF6dgrcykPs5ZFiYuj8eaL5OHW26BZhScCeXO+lpW
ChQxyEuNtrwlh+bwHF2DL7onPLxQY+tc879sPzgaUB5oDriqv1XAbbmybTnbBp6+
c6SbRmA19gUxX9F8r6w5Oakapwz5SdrVaxuK6lOl10TNR1ZCBdXkPimfsXICbASP
kfqnt/ABB+7yYx5K3M3L8/w63GnPODka6aaNrjyWokVuL8ILbzZseRD5e17oIpjT
zm/gNN/tE6EIu8fRlpaDFgbyvBdc/GTTElKtk/7XWEypPdpt369mUJ37ygMF4pAC
tBYQLCYFyT/wvW0KUKPO8405IhbhedQUjMnAfnvWdP3d/euMMwcbaVhqwj/i+Po1
jf7AQnth66361O7tJ5n/7wqvpI4iRVJKkyxxpLDRf/ENcg/zJPuwE7PqQIGI5fup
EPo1s94HCB0RHvdjkmjaG3453lb0tTeEXVa3JIqU7QpPXT5hZJnYGHMcxNniwRjE
m8sZ3saVOIm5oYW1JHX2GOD73vNP4M2htdtXbQ2qDpXHMemg/Wj1BJKWDD4K3YxS
aeB4f/L73U11J/un/bIU1dL4xSHCXpgrT2edKnDVfJpeAW6hV8Ohuo2qyaG/6+S1
zU0034yz27FfrIsS45FCqcV/lxGyeIg6dAYq3J7NU7UrTRnbvx2cpdsboTCNuW1G
nnDGc1S1ft6jkIHvRcYBfn6ZO0s9Ij/9qxvUqixXT9fh958nsMdcvVnW40E9moB2
D38B2rXGF7ju5NZ4FYozS/JbmUB+oNvJLGTxH9YhqdXsusJAsiw1BVmA2gVhwuBC
DlPiqTzUrFIWJaUGaYBlQHpW37SlxwnzJkbnep4/9Lvqvy+srk+jPEla4Ck0XV1U
z6aNtDoo7Z72eIRGqDDhMiOm7qJwu+meZJGbsITs7kEBs4Pk8mEb6codVuHb5FnN
FnczP0stTeK4D8YuhbxGYo1w5OIkGxjRdi7k5gxIiR3q4Z1OOuVlA5kCplRbQAIn
2myPyEHbJVk4PcmkV+g+c0P/h/vRjiNzbys8IBS+a6LAkjmJlYdXtp9bkQ3QEZyR
yhNErz6F1/58v+P8zv1Gf0JUVMCfvvnUhOl4pqvSKmIOR06u2cr25w3p0KtWCYr4
LFJd5tPfCnztgeVS/i3RBEJmQNqtncGQS9qDEkoIx1AsB27wJ+VAnl+utHYREAeV
Ac48Ho3rSZW2uafpLnDUeQfT32bh3XQ7dh9GcPGm03SHpI6nAALnK+5Y58kQu+xV
i3ISeaF1rJ4Kke17cBslvhlChe2LAtPAGi52ieuhJk6u9ZitHG/Tc1Yc4E1UeZeg
Tjc6gHCoCHmrBPmtg6DO1nZEnn8rIkTZ7MwCaIoXWRsNDJXOpREEpgTLyUv4bhFR
Cj3AHdat2zh6DdMCtn3Z/X4+uKOSoIpSiM7h1r6V1ZeBXH70R4oyfhPN5aWHpeMH
RTXgoqFwCOHBE7GBM4VNG81fS3YQVv0NWmiTYufg5biMt0cP33c0Epv+AqtxZ25y
cbY/CMShTOHmF25hZVvBH9hTKCv+pRy+NN/omO/xPEFtjseAlxxL1w3XYnOJ6HW2
O6stPiprAdoAf8i7LbCCZ1Gv9EXlc/+ZZdY83ywG5SpS6qx2zZO2LS2Nxm5/SGYQ
uACpVdCKF0pAsHcYoNkLAps3DXB2JcK0/i6vy6QDrCI0cHqOtzzziEBvAsNqC9cJ
6ohHNR5AWOxQfVDNXgsNXMyjjCIayBxPoOXf9ycMtBjKLx/QZKM120PS7Ve50RQD
CUAodO3G/ohjHsUl1zTpp03yr3sdhkAjCGFOKCz1GxkyMZ6+znBP1qC5v6dLg4hL
aF1pjGqRV70NZzk4+Ad5bNtCbEVoEFdkxOAJfDI0GC/iQoSBHVGsOz7HDSRncmUo
LkPw8BOQrSRarG5KXEcKm5jjjZvgPiB3nu7BV00Ev8j+FS9zEwkftcP9nldypFUY
+Gjrcl3D3rCivcpemq8Mo1oSY1QqxCYSgc0lvzq7FCfUDCoxE0L2SYN9sQ7Rlpui
+t4Aq7XG3SGbEbh6WLajrq9EA92IpEqFwrHxSwkgxjhH9q/DbcU9cxJA4piuAg0s
1ef9cvQcLtf4QHcheGaP/0LabEr74toCqNQ4L7BeQTE/Z9P/r4vGXWNqMz3gsspF
rdyjIZ1zzJnTAHFn3KW+MUG2vIMe3cnrBTjH6RgmfNxxQdLeRMhUe/UYl1N5YFvj
75xWSOQ490cgBcA4USXd/IF/zf5AA0/vbDSMHWFdnhctt/GZTztYoKAqd3QkABVt
KpFBSmINRqLxcAKwuc8qBw7oYkpLcN+VBIdIJdW7ROoVNq0+zkHEJK5LLwF+eY9n
f8j69l9ZQ+dR0SFRcjrsUtDEpOSppMbi2TCv75JRwB9AuZ20kPBD4DP9b3CKueKN
N4lc+WQw5ykjwtbkEj5Te5lHlN9PBstbaX6t7tEpEG/HZleKYD82vsLQN14ZHABn
GddUPBhEA8lkbpw/FThD3yk3kbaf1qmezVz40M+8WkOGVBFyU0E1crIpbmYj/KNV
fxZknR5b+VXl+TMC4WuP7xzsq1lNb9albYTZacIAiGvPnCF9dPwJx6IxH6NhtBQ3
xmkOSHuGtjbfzNJmwivq5FCKu1tipanj1t5aIepOq0Oib3Ixclwetjilx5Iu4i3E
9bCcndFk/lMsjBqzkE4LKsxHaaL0xzrgWQm+3xCxhKlF17dlT8xIPWkscsKlgY63
eA03NmcAQKsAgemiPdsXPo048jYKqW64rmijnXnbohsej6aWP4j+8T5YPneasLHN
eNvKFc2zxOyuLczpguqB8sC94Wtk71tQCeUxzp6T3F5wJizKhIHEB2yXW6cgxpiD
IkIYskYHRZhx+/KFdtc2hht7sZ2kDx4AOG8ops2BShmosF1h7gFeNNsyzKzoPBKk
P3DXfxLkar4h1vu0UfQz4pKO5ntvNNCL/X6BXykmQfgS2xFxphCxsy5/odgUSa9Q
PSlDNPsPIfbnK99prSfV5AXFfHJIkxkzJDseXaxUPdYXXkvFReeJ1+9N9u56IUJV
odXTjzExgODxe8NqC8p7TxWRlQGB4EdmDH2csGsuRokvcmT3cirBhRzXbd4NOjKM
HNB5xZar90PrMwVIlmViT7DiduKzoXRlK/dHQQTjQJdy7vLmXYx1vhMSYznLVkBK
bNFAOlV/jeD3KzdFIJH2RRkBPaqkD35PVqBKrqIzpireqYxa1sVBI4vAaKkfPer6
OH216Ic2xxlG2RlRG94mrcuxGlJisatVjZrP/yp3ONMSVTtkkXGxHb6OTyqUFPMP
3GanFivqIGGbrnXkfIBaSzJtzbXWdmBGzS00Wd2A3BLW+TOpoeYKlN7hlvjjyahL
vUmY74wkDyCv36awtcAKTeFR2JvyujAyooQUO1NWKUA/DhEQ9cqRZ58m48E5jYyN
j+fLgtoQF9FcfOM/9mdVZZOrUy58dnVcgbwCm/6Np7PiC9LoFWY9Df0EWXhlBzYe
7ZNn1qWIZaQUeXT9tRU+K/2Q/g+WL9cIETCgYIknE1HPyGEYn05VkD2qUfTnQKPu
ti4vmM065lUtPtFd9E+58D8xXhMaDFBr9ZVy44jeS2/1jep3skQk7byYgW4UdgDr
HD8dHTG8VTum38Vt88OdxUPLwv8ewoXE0SaQagMY2thZpdqUBOAtSkhkycm/aVTd
I8A/H+CPaHTw+6jhbo71CY67qD1REWhNQsnRQ2/WV2njO99YOFuxflpao2kjovVM
K+854UcauMKW/WOud7uQFOLOfK7DvCJp3v9UmcJHFRmhGHmBQnOL6hScbURU1Jf0
Evksz5qMbT3S1DSOBGxuHhQq6O0k6+gvIdR2ttoXydRqhP7dJ4NWeCZC5FGVA4hC
2FfHjL2xyyGASbXVN5bcAK1S+kXEd3kzYzWhSJAkHgijNik31WaPuPRog74enJGD
MeJV7SFViRjiXQfsT8mJwWAJiDFobAsiqUYgs4Dritd0hpARktXC6R5Zq6BnOb2P
NbvBxkG5b6orjJupUinuuSbfc14L7gzGN3CrGK9fyxk0gQjw02M8hKrE71ZhPjnQ
dRzYDeKYr/A8klfWU3GwUHVLQmpoea8d3Ezbpf+dcP4t37DSdIUv7Nwci3oCHj7d
io644ory1nd2D6md2nflxfkfSBK31rdaqJ3BfJemkQUHnxsm1HfpH+dhvjvt68pU
Er6cQx8FYrwkSLuA2YSgZFhlSZd/aa7JyrQfkuUszAYS9/Du93h2FpCAs0qMUglv
0+hf5WTzhqXTN18SdEf1DFAZqOsFVrzsfvbEtOetNN/vyAWgPQ4NDdNrR9JWG99P
yEVfzLcuwvCfNQchx2pxVplEhh5kWa6oukoapot4OqEqBrbl5zQF9n06E6wQlj+s
0MJFpAmGMiwhlU1YwGr1fxf8zwZOsNRsj1Ut3meBIbXYTy8FRtKc24NcmSjVMQHw
xWVqk1S97vSlbYMANrTHz8z203gMyAMil0R6QPbI19vLqbvJIRdPbeAzKs9sbnaC
jTZENI6iutwAshJnoft2csWG1q45WQe2V+g2ECH2nEVBDHDLkgWELg/cxcUtMFiS
OGpFE88lB8mYoBihG1XO0Y+94QnSspnGShD1+u8mv2l9o6jIdKty1Sfm53lWaef/
+91LPDZLW0PikzR6sCwAN8vvMrytFY7IwRncty+vp14IbSC2nSF+1i7NGlfH0iys
E1h1f2OIfzSxlLnc2F6cyXgP7iQqXFBWdUbwogGYAw6DcH6E3NYFVHWW7ncAThYN
jEKOyioaqSFuOhuZcFBLOoYHivDxiSfVHeLkIvJhC8i9NUBaGsFlP/AVQbXEQFld
58iTS22v6eW7fVAZmB486g3D12DN2upBHoDszCH+JuG1HcrgnI10PXxpj0DiWqKT
9KGf1J+XcM0oGHDIC+1QJWPYYbfT21El1ndTekvmQQBiM4fEz6qoYvSaEYTWduN8
zfO/EDUBlZxWId2VzVo3aTlbnubEGy2u+ii61J2Vkp0oOyIQSrztDjDUvkk2g63d
/h1fru5oA3ihR2SocN6sCCl9m18Rxdr0qSzjS1W7ZKv9lYKSbZFYabSiYQLgyP2X
k9XKVnKS2DF68tKBnTWxYrlxoBqrh7h79LlOyhJ4I8ERsGo7XffU8oDzGzL4i8ya
1XGZN3nHLKcjntBQDt5gFaACJouj7R5DxDqu6XwbFGo5ySdSHDkDe33L9cPxAroK
+DPgONMzgUanuPiDRw4/RerxFoAQWqnwnFvbiqLK5dPWrEhkpPYlV8UPF+zXAikD
jO5E/JVj516tPx9YZ03pPlTClktXxvEhnP4bu2u1kZiS/nwK4W6VY2SCVSxUSvph
FCT8+Qj1l5DqPbFOZWqjJiJnT9CUU7qSCVACM1QKGSGME5fvfHEE0rZgALLWBa5N
xsGZaemefUjHgy3lYKY1OD4awlqkMpYTjpw8gxdNynoH9mIQ+JbEnLl9cWSiK730
ktDMzlIPXUyzOW5wD95kpZY1L4WNTYw0nf+Q8uasy8LdOKSk0VTWJpWun6H2ijFO
srpZaPoKcaX7DFRfzw7UyzCwjwvQItQwywdbN/tzZiVdOH60GfuY1HSQin0mx+Pi
ToCuPv4BiVBpCC+obZX8Sua0ceTytZhB0DiA26Dbs37TQ1gsbmleeEZjWfAfbta2
iHqgKXezj6uEcIYWyA0tUv5/VntFb8EQdcKAUyo2x1ZdwjrmxqqPELLhGnpCWyc5
QPYhGevmbIEWdOlSh14ljkCyt/qzJeaLtx4zeEp0SA923gt2239oR8AUvTKMgU3s
eBSn7F/eSq+hY1V6nXM+q6yMf9oPzBFHh5omkreIOvyXbDhvxrowBrL+AFh1+oy9
diE4iZg4Nt6KhQtMMO8+OctXyifutDsAxmx6NpqoNgHfTdpD97mL/UEWpkZFhy/F
bALnNGpI6nHbguB8vtdD9hJShuHUf/kPnmqpC0VdfG8RHZakqtGVG7QG7jVDplDG
uxr/WVYkiKI395rIOP9QP4vh+u09izO7zvWKVVnaBnxYLUooJ3G2O44skcWhPCF5
gSzmfD9tNa5pP8ampxnf6yPoXvB31dhphxD2fBzdW9QGdEHVz8n+ydW4Dp1rF+ze
IcYlQsWinkQknQC4hrezskFwfH3tpnSnjFrQgOU9VGfFIKpXV80651CIpyoECCHd
erDCMQPq5VNJ4i4zfuScNHgYN780hHEk2lB5tQAwUzEtSXTTizbRMBoDcD3TBX17
hx/KASxGe2EcT7x341SdP0N0rn26L+fHZ7PZrhoBf0VOzI0eV4mRqubfpyj0Jm2m
ci0a8O7kkyse61NuqlR06aeq8u9B22z1ESOR1dtvcYFcW5350l92/87z9akznZqV
FwNMiYTVO72elfDtMCOyhY/ZTneXk8cSz/LUeVvXkygkjkWK/vmv96cSJz6XU7Ma
PuD71CErnDfgBvHFSg2iE2IPPArUFmBDYTxI8e1eA7qur8IkSbWj0YPA0NNJ1eSh
KBdbNHR2XRFyhVcVYRyE1cAD2fBxzrQSXWxmPkdkxyvEyJ0RbyiYEJUGNCBz8qvw
rlfyBa7vekyroVq5wWF/St91HYyKs32hh4y4AY44DCjASr6u+J7ODKfOJbNxyyeY
T9YbZ0K2bDuwT32rIcHQXcmYDXLIf8vtGeRtsajULtbuxFP+kTFsO3R8Z/zgTMaU
4t9l4mcC77ULUuj7lU/p6ghMuFglZUjtrK72cj8fiLONZ10iy7vX7NEYLRitormq
taSkkvXh0WLj17C44ngscuZvSHjY7N9gWpsIHBzWFOkRCKI/gkKz+RoRNiwYE29Y
IkHCIS8Xsm2oF7M9iABEhpPiQfyjdLkr7HGOvmkWNocjeSEq0XcqchS3JxvekYFQ
2jhD9Pf/xO+AchPhHjJAeay3ZJWLFfE78LdB084tKQek1iTIEYyBndv2rJoeOND1
stbHHZVfKgCNWaVqq3BZDjmIdG4mMRQi+7ShlW+rZPWRT3091mR7cLzW6mfrd5sE
tOfDzWRoazIdnd/D7PpT3/OMTiAQfI8mbEtvtfcQ3jwIRM7xCJ7FiLJyIr6488qU
Rf8g+ubhL1JOvkY6xzav5qBsPEj7onyrpevsI28AHr3JCMWu5pXJb+83CMMm/MD6
8Y88pzgJUMLCy2lq3Ge1KBlc+Ii2Q/10gCYI7C6oD8gt4BDoLw4gEdJXWe+gHwbS
Zq7QD8uJr0A8SkE7ZZ4iokzAlISiOeOkfT7omDugEvduK0UN4kV5DL9DOxVOU/MA
/1ZGBehoQzadUMiv8saHdDBNoDSGD0RJEsCLHz0oP6nd+LaF4i7wnoasmJl65fB9
BLSxvTqzUxzM8uoJj0QVS3Zq6/3LsannlkSKZlt0JGAZyBLxjkqkVW4OxXEmZXaw
erJyirdRh7CBDUOu2B1XnQANrpT2xUXAXaBdXZZhqtxnu5ORomkN4qPtHwrachKL
S9U8MdPvFcGKIlH76Nc/ZQyL/Fkv+fl3vRZ8notyzHjCk+ZD7XYEpSNpwcAnQQ0T
Id/GbKQc/IUvha1gFFiOkF58U4rZyt3htvpDyAdpkaTL1gAdDb7/DbGbZhYI4Ojv
Smn+ZFHlFE9mwmC6LXQCt8iN0my7rDLMAnkLeTIc4p4Xd7SN87IBhwMVeHIZOLQV
ImHmYCES0k7uxqq+s8rXYf/8dagmCJNrkVCKaVGWQmc0KU0UDn5qv6a5F3Qof1dq
etnG2PLC0AUL6P65teeS/gcB1cWUwruDwGPivBC3FhYPn9VP1YliliBaZPJaunWO
tfVfl+58eWQ9g6Kkd3WPM4hs7AQjkd4nUh1Vdyt6tpriVJtUhsbgygIBzEg7145/
PkRuWO/celc+RJVgd9WeYtOcHgRdaiyFvdrhOg2DODhP2VMFPHVWJ2OE7Q2zE2uN
AacNbPW0L6Xg2se0YORpPLF0bCVzYEe9NTXAoev2ACgqOxJcIMMFfmUwbpbzAVkj
e9RKniUTgo6cp0v1x2rdWpQBY5+kg48jALJ/mOYIH2WRnur+OKAPa+8RbVQFwWiK
lU4f8nJ3/ErlKX/k4+X4Ybt9moGRUzZWQBlCDBUfLimfQ9jnk0N4xP/Jyr+N9rxc
4ktpypsxZ4G9mSlILtupPB/V/bO3xRHOmKi0pUG0Of5uZ718OHHP/Gm5KVgR04Yd
GSijK9IO165kOGaY545wjXQlcqsNnSvAQBqg0FnVOUZ6K3e94UatZ9Gpzn2KDeuc
Xv6k9xT/dLAg7zfpycfsUSg9Qolh+ZRWqcvVT/L+3RYhpl+ej7nh/qOeGnYBGm5z
wVU4zhS2t7hJNY8Mm+F+VO8HEe5BalXA56v6L0shDMVJk0u6DJRMGsrfAI9HX6ze
QWs36FLlyigicDxrtMvYageWsZ6yG9CZlBqLoSSn6vGCnYUvU0pLwAM7AkXy+esl
PThcq3lLFOg/4oTrBtPKL8B3uphY/2YMY1iSPsLrN9gGFbUXsKND8CRhF/Qzfx8c
qvgxufdNwNSaa0CQvesV9JfE6pDZvXuzRdFNwak9FaLy+axGnb7CkbkL5g1mJVci
q7hIjngC4DYt7rIMCn8BLipn3luTS3IJJKYzzy/S/n5gXfJ2e/7Nm5+LEQuztWq0
sweLu5ez4P/De6S+NtcDiT93hz1P6LoVR5uYdRlBRSbW4eQMcfXjCDUYKSCPw5QN
ojN3UWzDxWx1Wxa345yXuIJArywQiiSm0c7oc6H85zpirPOoEwg3ZribXH9lye6V
U1eRqE/uKWRysCjp33GEcOeNG8JbBZQZWnG9Cr4DE7Xxf7kNEvB91mxFBttcuenT
0fl+kX2tVUwX/SGmtno6NP2cL+LSjYppNcXR5Gxy50WWXaYywgHk/tvRwQKoL4qw
cUL32S+J3K8rhfXRaeMGt7DD9H6xn3ynGi5zg8+kxP1et1gVuaDq7icLnn8MZr4/
Y8fAo64kdstxLJf4lHomNebSSnBI3gDjmSgCfWr7gSW1MWYboyq1JrWmyCEudmXY
RFg5A4oLUeMZPxbs4OEswh30GHb/EEvPwwEXf7r//dPH+vQP+YK1nklIttygBX15
bBWra42i7CIRhQzuf8pKx/d6fbo0tcP5YK4LnSVrwcL3HCQpuJatJGjBmIkuEZfK
AgybtrF0IUCEZDQx7tIuzjBZ0hg5sXg8u1HgM07n51qXG98U5ToAfa31mU4vduRI
/AQAvstVbM+0X6M3EMlnhmLEwc/VHzPdYuAhqzpkK5lp1R8uKO64f3KcOUNlMg+V
l8nUnWBpEEiL6FcdPEmcP3pT9/D/6ncLNPEOuuvV+4dMHYHiO2ll1vp3qWCbYRAJ
dNigTRjyh8UFvsdSw8PHz3CKeQdFuutT3/eHnYqPK5LKfgMeEtSLMeESnbdXB9ZQ
/TDER9dmCHoKx0wMJZV4pxXP6K63fdNgeV4h1EBfcIbdeEYMWnH5V076omHgyqjN
3HVwUuRqbgEbkifImcMVDy1fGoKT34+Dol2XxOl1I6oVfnhPekLNPDWk5NeVO+hR
HN+RcagH2h/UO+CHyoj6NCZqEOiovuOPfuKxjVBM9qmHRvefaRGeKj3vSWZIemJ0
7TrcXalcD34MsputfZssgdW//JQB0M8FtddtAtWFXGyR5w+DICu9pjpUOHkG6lev
eKaWHQmUdv9HdINol/xuDA5z3upEHSK5c4Z/2vyOvnoXbR5bfRcQsPPyFvzyb7OD
md+633NhjJ6bMH0R9p82ksFRpCxiksaTM7f3DfBc7fX/XcFweuivcfQ+e0zFhiNf
voaeoMwc5iLp5HfyoSpD3CwTPlTP6udhGEi5EK1FhphyNlv+ipHhgt1nrdJx7wFj
0WKrQTVorFcGN5IA3LiNSNi3CiKF5t+wGVUKvq7X0Xlqk5g3hC7Du3dYtZzP/pTW
zjruFIzkyalJyfEgJObFW6+H85AnoBHbLx3NrENq6AeTE7uy3JBNU95RNuHGNZCR
zBHeV1Pj1jeC3b6CWsfpZVqQoK/7C10jaCMjJXhrmHnNNtUo3rTKMfVf32j064Vt
48a32f+WipMLA5I0JDeMlVYciuatQQU+bVjYop7pIerLUrXVd+aPpu/GfJGwPRLO
QiBBXWUcRR7q4QuvsIkO/UZ1ryeKTVJf7FNkQfjJjAk9ACih5KnisOrSfIOgfLO0
k/t8Byp5x58V6HCa2qwnturKaGCUFydXcaAcv8lMKuVhC6dXCMZcu3Brr8PXtBmU
oBhlA1aWk8cdQS8/A050Ukhb7seiRWl1z+o/2JPE8vV8kE1AAEXC+KAkB7wJU+CU
axPAPXxOILYXBWmHsgphsS4MdWDZng5/7wTLPmwCz4MhHc8Gsp61dywU0WYJd8uQ
12spoXEmA/cAmRylcLQ6rl82MCZIX9L79F22wYPk4S8+RTelgmxQYUl48CgK3enM
4CTCW77yrCIHddR+iElDxiXMFVi6fUO/7+6Km10e8E2WSmRZFyd7icxQFrE8dIxY
cD7WJLM5V6L6KC6wq/r0KBy5FtjSn+K3pSIiCoPM0s459Js/fp8M6A5TmPZRZN+k
AnBrEDvgnV0G3c4sO3DSnz1QSPt7/uVGV4x1snCs1tu58w0rrdqX6IACYqTePV4z
MTFmjjP+S5lfAruGEYwN7u3slpmk/eJ0rRzOfEtNMkQ69VdZ7DrNPMvR7823ba33
n5QtQEILvmJk6unIVyTS47jBFv4Nae2EltDuLsiNwffWDTx2b96bZsTaqvYzT3oQ
eC22kukgMMf4SCxSz0fXLdEu97OMBOidwnOnQfBHVUDi/duJ4I0Ao1PidEQaKkm+
1VEBR6mSqFzKAgrH6tN1zy84dudcVNut6JqdTz4wSrJYVR99m2pDiQZ9onwcHvox
Rfc6NeZTuzO83HlESYmiMA+23PgnW7DBhbevxzEYmqaJ662Maac0BEWiJJkPgXpZ
qI2ayUQS0jmS8KdaB78yyO8N103DALuQfBMwqVGy8GIGK3LLUdFxaPpa85uTAHro
tvzTVIoQWbC2T4rDMUVhPMcBSgDoidzSWHiYcVO4dl3opOBrE0g4fMiTfIgILf+Q
IMBZWZFNGMCgNtg+c/e6Ec4p06OeFy2zSqQfoF7Vbjg7o3Y8V1dms2qa8eYs931O
/J3myKIlVPIuoPDwsWeiXp1/ZO8zY+b3upwsC0ZpaSxvhl1iJhEC88bhewtOFmi3
S4hW3rsLTgEFQW7F4t763wsfJo+JOnb6oBBuAcdf9WjyECRO/zlripaZQg8yQaFY
pRZIgi3nQbKDU0eBFT4wFT2vzdio+sitccFRHwtjZ6YfQtNREjCCOiX5orLtDQHn
9CT7t7FrkprY9DLPvX1fxuNEAtCKueRFsic1s4/yZU0wxHYUZ4BWQm/iq4MRMLFk
ggasAIYZZrGaFkfoGvmMuundn0FjwSRdS/BQoIqNjswb/5OhIatPaTF1rYo3FEwQ
0wivlejHFDvjNgM3CoptHuAdvf2/s5QhafMydLBxLWRoIdhv1LMfp9itu3H7DJH8
Ym7jR1NekgB9r25olLqRcxwW8wqaxMCHSvPzG6+yp12N7/td/saZTP5soI2Uhbm2
DkDJdXKydI5MuOfB3ihyRSnIXUtJ/63nj0k9+Cv3Hn9OLXjuaaUkQ37kpvpnPpTv
9kKwcnTS9JtBVl5/EielOOVGQX5iKwwb8sIsJV9fQ8KEA3A6cVPuQeOxcQgKCWTi
c5v5S2THIlctSUPnotFr72DrLbU41SVJ5L5OcTTgPs+i1Kcw63cUiU/0R5hSYXMg
N1mq2RnZyV4xXin3X2Xx5I9N/q98RTW44/2hxHUlR4boKEswG8uPE+yD1V+Xwmid
uZN/BVD/6yWI9JZgqD/ys58vqShnkDAOfXQ5BDeut9pA2tYHzlk7SDZIF6//VVl2
K6O5SmbI5iisAOLoYbj2F97FSSTVR50gxJqnRsgaWBJmRXauV2fSR6A7+2NzqnFa
E3lDEtW7EA/yNFF2Hr1ebII2Vd796dXZQhj1Mba0NI186XGd3oX6RKjGHQ0rBZk7
qkCe7QCciaUpmqJScuuL+gfZl29Ae0nbn/eWP0FCZdKpWlCs7+WxlpIXFdHNsY+R
tZPAb/gYQSPzPqc2FqfdcOX4P53VY4uZBYts2VCUtfIUBuZNc76mZKoUp4ci091H
cjeENBTUmwPnd4AtMC162lvTLZirscTJV1Z8CSRBUaL4E9rJl5P11p4QP1IdsRT/
/r9vo1MMr/RC416joQggGr6oq1wPput95w3OU4FuAfpTQY6711NcN+NWltjYG9ec
Rtt2l4Hrxk9q84NpU06xiVBgWB1SplCHIFXN+ns+C/oZhhy3n59EGVGz4oBwWo/x
NY/z4A7VrWWO7ur97P8CDOPawtoIfzzIXylvp7W0L4o+AVsbeAV9Bvk/uSkW3Yve
4D8EZQS06PuNSA7GIrmNAtal2Ho8+R2CC9HFp8KIuAmtCPdQ9LolFTke5c0tHnb5
VIdATRuKLoNzffc001IiyOpg1IFlJOzc+49UAXBkjFVVjRxprcdJC9o3miGWRd+y
JVwzTjx6cUQjmblOydHpv0mSRqQuyMb1DbJgWKkwt1YiCr6ibucG/eMZTbn1KAgY
zj3t4P6kH8UlUN3Em773SNL4/o9KQt10UeN2lgBygD0hZjwm6III5GVL6l9UYGR2
1k6Ocl6GqBmklIM9swFcwTpJHJrvRqTPusJPZLmGFmATS2bK8p0wUebuU7SQ34K1
2ENFdmTpP8kcMgK+YtVinVEhzj7KXGYdeSvgEc2O2Jdg42GOOMzUs2cSVpaChTu7
e1YtODRlCK+sLxFl8U3WEa5+nUHXrgEs3y4NMX54ZU1OcC9H6ROTocMnOSOXLga7
vX14GSEv5dpwck19sWZGBeqxdCTCMnoE9Nmgpm5iOcq0SQr8d01kHfpYpF29tOic
sGXSp0uzluuUsPwCirhIsT94XqjqH8gaPFwAx/5dZ2tiuvGYMlkjTLVVbKuWjuHj
wUnVKSzCG1b3/5ZTakKd07oK7Ze2Q8VQ30w9uLFDT7Kll2Ekut+xXDtjK+5bM9Kt
UfFVDf/sqqKR8rEqYOBJnPgNGjJsCyW9P3GpuRXoxuNjTyW+iD0wHVl6ifOFmCAU
naL1FAWTv1tlznL8sdHe8fvO1u5PCNca7IdjRK4VrUwylS1mce/bua0LKmKCLDEb
bArC10zjD0A5gPolNw3dW/EdO1XQMosqWo1fGECdqDYF6rjFKGXToMy+k8FSenS+
QNoQABWZe/iDl2gplDTe6qdDFo++2G0NIwEqvdmbQOnygfDzN/fmVu5ujVr+joMw
9M+Fick7uOcGlXdomBIBp/slmYqGF4I3NU1P0JzHP7Tvf2w/g+3aagjfrTXWQp9O
Jt3HmJ6mZMXsK7zPNBSZTgHVNxg0vo1eBlqG59hshEGpJ7UCHl4pjpwqu2xtJC+g
0udkB6+xMokXWcd4AZwem1SiT2OytMytiGio1RLtDcx2qQc8EfnmFkg7JNRCqawU
sB8w58SfKyEtu7Hu37XTnEgaNw4PCI/3F53yXULkIlx5pf+KuWase/K5yUWdkghM
bL/iinKvMuvVySLzn39f9r/gWAPpNfpREg4qUAq0Z/z7RgXjlOxxpdJ0b1Rdd4y0
RrsfIp1EZCM+40Gfr53a9jUaoTK3IcIgcegFB3wS8xgjn3lV+d4rJNq4VlGGTCBZ
iREVl41oIfXHarSchdHxbH1uO6X1rgwgqYuEztfvZ5zA9682mEbveLTgxAOJQLgP
aS7SQJtB0FokQaZ02DeqHRw8TBAaf/2TFmEJVYaBQMmG3QsvmPzRZdBcvb/vVsT1
Ofx22FMGinMGdsKPW60+aJo7zvU+zxncpxHrZ/SDC0EBWpD7xuYwgEY6Kj6fTNM9
Y/kPPAiQkEqpRqYdZj9MwLinMnf4dtaoPkmPHP67SNTl63zucTpqGVjcXlWXzjGB
WF9omEOBpOqggeq1htPnygI61MfEUjkzcZTCf91Sr2oihRx88xY7i5VjVHk+8ApM
XvyUL28bk/hjlAaBVmeOclE7FGjLJwiOxVYugAUPyBrA+9v95K/1aQBellUzNbmc
NpVW6ho5hhzZ6Uj+2cnSdshJBrpcg0WCL52zoHYW0QHbTzdfudOzNW89F6IFdsaS
3W+LcV86+6aYPWvJlvKE/D3TYvV0yDFvoYtMDJCBqnfe/4u70wlHEWK+ls74BZzR
L7uyJ1dbfwl4huFWzwTAVHxCmbk0/T0OtF1QPH6bu2ThIsYrI9Cg4jQsiWsy+SiL
e4CiA8eIKAC/Un63CVuwD4VcJzA2DJncogBVo9N7/cTG+4Z3KdtG937QCSHkRQQS
slcBeRbQwZMM8HK5WFYMRzYLXFHYKa743Z1VZar3Z2GCzRmI2rlP0KQG71vsPPqZ
JpHi1uc8uk5/zrNSL/kKZwUGVcbR1UuWe+x3GtOxmMLiM8Udr1r3hbPl1otN0DGh
7Sb2/11TZ4bCImDxU3Ja5DMb0gYT4lYC2/g54WVAY7wOQscbB+vKm+oMydwrXBse
QTqH1IUmq3i2Btn+DZdcXnyICIElkRJQYwpjDRHcZ4mPuzBT2OI1MitGbLwD3xiB
lao98G5DGb7vd9Ahkh91JnXPRNBDGZO8fcYPbhRUkzNnlgLBQXEC4u1p3UjUzqrU
3KxTIQKKCvI0j8OjMtJn5Ca8Y1Bm1Wk9BcBBLkD0K57VjCs30mrjY4LFS0YK+uWz
nSfWjS5aKFnjOT2p5BmdWMHoEdpFpUladM3vygqNOKYec1LeLG0aY810nORJrjHy
zsAH0AKgLtvoxxp0htwYUz6LVsXNbfzS9stR4PDb61pElfN7mhUPhYiEky+B+Omd
w7UBWS1xNOiZJ2ZZ77lMQosMTav+XjM0qTfZu44Pm8voWkcooPjyqtKu9aqXOIi9
asl2DR4e6EgtrRKYgOiGCtxssEt4BabjXIMgMUXt5eHrDQ6Vq1zH1xTUNgcxXKvU
SQ8nv+3luOlJfzerM1NAc+7oOYcvh7SRFgZXLLaC3nntexl3/67R0EwTZTUMjJsu
vbFkajusa90IGl/VUbNxh3nd13Q5oMDF4chm256MpTDDYZzriha+MeB99ksCwaQm
41P4yjAqju5r+N8MBt22fCZSkjzPCP3y4oXV7153g9W50Z7JO1sDOw2ybgaMl9Ix
zMFNrz7EZsdyvlvDRn/ok79CqRC8Mf/NDqNYPOUv0yi0pJ6sYwiRiiiuKtNnf1ed
k8oLtjlXwCcfC19k8s47r4JkzpO36WWKVrUrUcExAXGkuQS+r14tWk+tbKFLs9JM
AczQ9B6kkVjLae4zGiyv49FzdXz0oDdiBTdjtrWyO/EMIzUGdqslBRanCRqzzipM
/+p087DeQ9jTNL/TQnXIgD/22XofcheBac/Z1kdGyWjP5I8kEzPZH0Ap0b2BUeCE
EFRPK7u3O8xe6VpYOy7NcdA6zF42wWZxJ4PqzgDM+HQoZKHhIxTrGzFLgIuONxy3
qaI40fgpwNQ58QJcG2fHfuy15vuX2JiSpitr3KvvhhAfCGZtS9qJECToma1yG17h
r38ZMkWP7BRUB8ecoUyLxl2wfAcjM8YUJ8XCYvQBsTbrFf5KlDtThgzrEtSzp1Xr
2pdd2zSRR2NEjCJmjYFYaXXG/Fz6hr5xrLdbMSApHXbJ7it6u0rtHfMDCZlkelWT
hI+nCWFxeOcMCkL3Ax9Sp0bfgw0M0wSkj0eRRLTvNBsNcOUOOQnDZjajph2htPxs
HFnRJLYPTjIGjdmUrYVuNKKtDwu27FaW7HyYAiIGlw+X6HtOeE3/dT4DDFgsauv4
s8Nr/BIFgY2M8P3ILxDlrcCIJnqO7B6X5YiaA3TpI2yBM7g6mo4u8p2lWMcoJX93
PqxiPDxj2N5TABC5qffOL+L3aGdbkKBYBRAEfO+DO0WFl7g6mOtcY6YlmTVjmDVW
Up+9kRtQDAieJdGwdJcsvto4kg+EKjQhxZQ3hbmxGGzPlhVLf+nAqBP+5Ju2ynII
yLVV7XBGNTHBy4lbJDhD3ZZULKl3fImWuzBVMMbR91Is/4tHi5W2V9NNKRziX+w5
6YBNaT66qq++kJ+CAyfolrmmW1VS6LLf4587XjlEIK6VLCQjSGTfeUXMwmKeVBFY
8Mbn6Lw/FQqv22LdL6eowMImL36ONU4P1Fbdc/whaz7kh/fFjs3Dp+HB4SnMcwGw
6/xRMW2Tcte2yjaFR4xScjLo0JfkPn+OrGGM+EYgsE/7+YraD1Pg7bbgoTpynXoC
vFdxLqeEq6+7ayVpRt4Sive9JKugAAtImiHeFKlXNRyrklKyplw3Dirfmlazj8UG
XzGp5Id/0cXJuwWkZThu4KnjfdeCWQ/mJzSQz8B4BeZMUpRHywdQde7bUWvRm1nf
kzuw2PbWQTa7Wj2lPZmYJFwBGMYA79eyFTihimIF6srW2hz9R507tPJL70wbwpZE
WR4/9gRu7dx7pFZP4IQ+ouhhG6jJkHhhNHzQ4kCvie8qYjNNl1pDhzV6GpQvpxuY
GQyrWZtuKHuC0ceiWfyugpVUBs6+80xkdya3HBw/KMEEruZgo42Ffw7xlvFBI2GX
+hZ45gny3PS5IKWZoPRBWChIuxQJC6I7ZLclxyU4kdUOZ4PmO+kycvwgN15FwdHm
eb3ukTuR3Fr6w5T6LMigSXUzhFxIhOnWCtb3Jqy2i+DvBqC3o3SvA3ZVVb3kpYSa
1DIvrQkz0Qz31vfSb6240RPRexSvAbDo6HbJ0SeStY39pkvCObN3MgjAtJK19m99
49gFwG1B9I+99flK3zX1sZGbxm5tBWFqB7aDdT7f3l/DeoiROOVdHBACBsLVDhNP
NS/Oa2M3BW28onOfptUAWKGqeSvgxgSosD+mZ9sRlE5N50HAJW/bRoveGMsjFyes
McoJRLXYumehEruqoW9R8uIg1TLBQPs/tIv9jcy2r9lklanlmhyG+Dwf6peG3Jj8
bl3XqRvQT+OkmuzQajRpspBHPiKWuFzYcXRxpTLWkIUHm1CNH9Mr0R6wJ/S2NNIJ
/hwDzU5RdcBtGAI0DLdoyL6GbNOkdTyIDhVyNRR2cLffpuRpZrZAKjCkjujiSFmO
qHUGGnNZCQNedDG6FeqA3NRLrkIE+gCVSHedxZkQ+E0IP6q6iUgvcyOFfWWkFpgY
bNn/iXs7pI4UtzTZta6p7buVZDsrgPD0ego+dHnqVyKL1cN3BlAQuWEgLt3nnZHX
PyhsueZCJLuCfnpDIMjpZXOf1+7XluJpLwzJrvnaVNhIXuPE+Wo1JZo1XlINNtjV
793f0Uy6KogdYJ7deKZ8A7QJ/fq1T2pRNelxhrjgFUIvP/+GlVt77iX0vsPN9iT2
sB4XQ5DHL7OTWohTaJlY6bJgQIK8VNpoopL0Ju8fUu91rru5IeVMgsTfHDzxYN9L
xozUlhmvxT4ag5uppMgTLjJwka4UghZ9BEBZNzgKgqM/rKFhQZhdXGl6uVfeXve9
jHx9w6avel0mB9Wr4xzPRuCgZQqBtQjaJLhqsVXX5GC3EvdpN3Q++XqXia7IMhzw
vfSe9GO1dzycxlC2xByB0Stx70Ba+t3/gy3qyWUO2QM3xUAEy6V9CVA0bOand1MB
XhYwI76AlIIVdYogt/bRw0LjcR+Otjb3h82GzbNMvtBwXJPqUdts7QVoSQc5AHKI
GbJQkvQWZoV4U35ziMnFqA0bJTcrOO5n3OEUd8nxQIRhKcWPDgdMMz3bjIu0Ib/G
C0NXyNpOcPAqe6ELqLgfP4/JJvyD4/FUFjNEwBAMcyWR0OgNGryj7esAt5svKBSh
Sbrhy9u1Ssi7GHAjozikVwWZs+/As0EeWW9uu1FdwRvU6elGT5Vpu+hfvZRcZKAR
1YmqKoidFLSmEc24xU4P/am+CZezA0ruYxQgTeS9S589Or8VIORudMPmjFpvDENE
Sxmgap/x9/vTwmOoxqxrPw6YtIcHUU8CFysaKXw0Lk0ZWYS4a4RaK5p1iiIp50Rf
ztf0/YF6wBtykjqVr0t4oDYph5ceT1YclkhBYhaegh/AS9d7oA5OUnynandko7Kk
LAkhl0ryEowPP95y6sQTV0LDpFwbpFBC7mLbPRRYo8wsoeFQYXJ1ZpFCMawq/cEP
RjHSzENemt57nU58K7JsjegYXyE8qdkuocpZgADf/VafGGcru+gYKAQ1jvuhx4Fr
V8kKnxhDGLJH2wRvmaziAYf+3qSIouKqB6LstMudsw21+Ix+hT7MUq0mK8P5UPDr
WDEzd+AoFU1F5y0oa6NJEPj+9hj+qPFhQuS7ufDuybgMldxANc1oMTFxgpW0B/X9
RZ6kCrI2JhusQRQL+31v5OY1zkJYXiGSLrXpW9pXKnEQyXPIiBpWPsmlr6h9o2ki
7fJ83D65TM8Fk2hlI3l4gr9GOGTI20lDTvg8w7/0c/CQErj9R1NP5v2AxQFAMdt9
/HELZFD28gB924vG0z5lcdh4/TGIeeqT0nHk5A4e7qQjHtobXuwWTG6mNVLDSecp
qZhLHte4EMydYzyqnJitptt0a8YTa0oxfqamGUzAJVxFOeFUgaeA0Y14GffbgR61
RaXhKKWsU8SVue82R9+9yV2lJN5Ced7vHSgaXxuNJmMy29Tj4RL+dIHMUD76lr4B
zqIleVEzhHqqW0hn56qSP18NnTT6Izjuft+qNj4Hn7aRoqpDkqWT+KCdH1wAkCt0
uKQlgGweN+QyVOh8hEdAUbWHsGC5V84itgUp+tWdV03PBMNiV65nxxfFANox9GhC
DvqiLT1X7XBc/Q7VmljtrnbYUahQqEJ+A/65VwDcG/rtaKhGiVQ+Xvq1kEKHmNz0
95d/IJrGP0yW7JhWPWiSJ9VNk8Iz4uGG6U0bDEob/zbLSQJOv9g7udy7xCdGKZp6
XJZdZtTSJ4y/zQnJInKsi1IsLNCdUUELB/aPC+738k91DPVz/Aa+rOk1w8MBe4y4
FbnMUWZCZkvo98NknYYhSARsKF0NdPfUJuaHaWBdkr1MV8jerMeErgdcctiYKWgz
SCHjTU4HJVryOyRybY6ymeKy7lDAiO+HesHllJPZqOWw2Wxtsic45el4yRBZYqr3
Aimq1l8KrtDxYpiW1vGBHgFzjJn0nSx6o9fBFu7Tpu/6UhNl4Mc0DozXb0r7hHdr
jzvZIu9007yR+Hc8DUG0C9HGH8zRqHyQtQNg6KUv4pqokH+CEqHSxWRaqn/2y5ae
mNUiZQlS0kRvYs0e9k0YMFnjaBeChQBB5dIrB7pFAPbcv6CIiZVE4hw7ZWlcXt4G
My7rJSUbbnz6OHZyNxvAtD/9gsfOBv/RF/P4KedXI0E4+NahLLY+hTDiLJ62EUUT
96GwqjPohy7rsBtsQogYXRAcWU3y2/VsxSgsO5MMh+lB4kSQ+LHNG0OlHqkf8dmI
yOgnvN4hRyu9VlnHCmiMjDscwT0t8/M4E0etzsiDhQ2sumo05reGlpPa+8zQa4Ev
emVsMgGi6AT1wMtFSdhWnsjNYJ0rUL7BuMMcwdrmIdmuGap436UlmvnKcSpSEOHo
jMWDG1GI3xdZi7RUjFgmw7TiAvV57GEJrbJs/E/JTEqkKikhL7Pqk0hJwG4yzg0p
LvHpSyQozg2RJYD/ty4m2Y9sN7x/2cXM2A8tqbmby46BOpPnoPq1H/d8QUaA/81O
HStj/p/um/IkB0t3nLNejgiPEBMYd7SEsmuRpXvbhaVY+1orAnX0KisUrEOFwt1m
BnLVOTKCgsm10WQlGg7W53KvFjEF292Xg48EWyhCteLKw7EGDuH9ESw51pBXsXeS
ZypB4FnPQ7EiICTMzdIFWySMis/g0gBDTOYWvZV2ZKj1Xn/AfSGTY2th1SGO00MD
Qim3j/jXfF9dF6nbfGDbphPfJX2kvjDxgPtBgpQ6llQXSzTejhsU2qK7J+r7pCsB
rWdo+NebK9bA4vylxg8Wj/qYUylpGtof1XTCbcnPjvE6jmKq2abZFxRDbmzSgjUm
ivdRyCwrkWoX6Ddee8ExpfoOzgvpe+ia7EiQXVKHM73Z/ooVjd5IVZt3lCTxsQEK
jsA21gf+S/3dlI0J9jXwd/YrJBlKgQkNuyqkE0IUoDvTRFVz6SPGaoa3ZJTWxdRq
zS6fItsSwOk7QaWEMbX/m5S8vpE/W4GUmqRaX6FPKP58L8Zn5B6/IzYqemXaClLh
u+ZXppXhiW3aenam/BnAwh/EvdZ25Y8oXZEpTYd6Uf8Z52sPH8nYVqqa991Tqb+R
y1NodQja7duZ5hKIAkm4doqsGMhkMozA3Md72l+GATMwJuqxs9wiquf88BpVrw4d
WfFKWt0lST+YxWiDmw94fCawkOXx4EAONF7pjk5WlPFpONyUCSGi3MQjb4+vpe9k
FL7monGwUantexGlYyafjitpGKrOxn+UqaL0XKx/yn69T2N86kYRFAtsICTtGVyL
+1kP71S88GbTsSEqVuHLnUqZPSPUSKIeHBHbswE1ORLiIZPslL1PeomGwU1Um4It
b+pKtoPQ3O2SywwQEh2TtgQRwnT/14xzfwZYwJ1NZp92XLjBzksJFBlpexHHVTii
ePgmWOt60yIU3J+JIIx8FiX/xcy3NHPgc1xgc4Q8EAL0jrDFreUHraW/hGA1qnt8
a9/t84i2bjFh2AYgb5X/OuF3yHfpvSQzVd4cPfm3qalZRh4gNRPkpuODnLuBSnEx
2rAIc2k/CCp5cKy8nF0Hm9mpiwtgiI/KToQWR8fM9w4cF1g/2nfaiR135b3uTEnR
FnHzPBKRt0UX8gAr/8JMqDsUHJa1eFxndAxvmKW+w6MoD9shxaqtpfOa6498g8ZA
JiFIPHIHctdmPukPvulgCWxvD9416wUuiiSIS1ttp3XYMy8Pe5RRMCpjS/07aQAE
v9ecZI+JrY6fa31/SbnoUx074XNkT6nv2mvgTzppCUAsBBYo836YmD5MCfDjT3Gq
paXiyDsQSmPO5gBEbib3zwDt/aoD3oNYDH0on4kEEwkBOfc1Nid+LOqawZkBC0Ox
09Umq/zT7GFOCzrJ5wTAGooYiwdEqI1GA6Rk1NTmy3/W+ApuJm8aopoa6Ky4Q68v
2TyevmPeVldxE0p/ZNrse2Cfmy8j2W1jBhgHh9GDUenmn1dnmO//pOElO+dTEqwv
iS2lqxLl+y7BqnjJa97HjID0opJcgP8Su5iitv3oY77+BGHcMwdJrdcC73PYu5tO
Ug7KWRhA//JTYleAigqYJSKI3HIQM032/4g7b1OvtaNaixmGgRubu18Q4oZZEdU6
7IVmc1LYQNGou2WetWLGAD4Vp9FL4U9+nmKQdMsEoJORfT9xqWsVt2GTbSmn9NKM
9egVC8gwdqZk/xXqMwtuov/m/x2Rg7iYpcJVI3Xyvf3kxMy4hTQa0/7obkPIQCT6
ypErlKBRqIgXYjeOSlPk8th95basOORkdNRhXoB0S1OMhdFOqPmFxlG3jW+LeU7D
h7mN7LiWHyLdDpn2+IkqMi1hZNgKxOthF7i1jj5VlEHO0G6c3YPsa1B/+PzUtU9L
T8v4Tbjkah4ZgJewXgVpSX2DaePny3aLos+AP4DhBwqxoQBbepTGAkq3hM1852Qv
4M0pkCqiFirH3LbCk1NBCwxoYDpxt2eGjBUwG0P5l64e24R+DiG7SKGcR4VWUOe6
M/I0r/YBGp8Z73Klv+0JUXkL8nPgGIytfwJeRTvReKgn+vlcfz3gnEMwx+H0U1MK
qZMWZHClLoe7Gpura6ZKVpPfkFQDZ0Cl83E+mRJN+LD4eK3e5ogRngA0fsexIeGV
ZwHFgFNLfQ6ct1/5lDJqWVIvXEstLu1pRuGcTv0WZWS+qz3VGm+7fpxoNa2ibOxx
vhVq2DthnbzI/l+1tRGMXzIEhz4LgF7atFIG368xukd90QbjbYezRbMZW84fYpXC
Jpaq39koWa9txX4//bbVA3Vxi5QOqFXHI4mu55z136vQHmC7L/4XDWAmgf4CGRnO
5rBABw4Lv2G3b5d+ZhSPyhS2dQ4uWlCVA6xMb1KfylHT/Xs0cHajMUIzXjv0aJUq
564mlzEE/Ud87StqI73f5yLhIn1JH5qtmJBA6G5FG2ZNmDPPZzQqqeYEK5J4JEDq
fY/vrr5RXorpej0Yn1sKX6F5iADk4dyqULcSb2yX9gI=
`protect end_protected