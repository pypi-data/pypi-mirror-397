`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzQ2ej/P4rBrQ1qSrxj0v8Hrjr19iTrKsfFSlKxIVapfw
NPC45mZnDakGiXXKUQZ0mk/T49qusLxBqM1nkKwyr9uAErgVA335Hf7zXww2uJFJ
sfspjuMyRpZ8/vygto2X2m2Yp/i1QQwdudJ/gb2/gHjQCXrbPIhbqu2gf1KIZP/u
CpkhQScm4KFy0vIfAO2bUE8D+5cUVby1RmbLHNfDhuHCk+KrWbthQYzh5WicVpXz
SVsGTJrPOTLYD7ZRf8C89SFVP4xiut3vq3FSF36lCcdiXGmn+VjVxWuBWmVaOjrZ
8uLs2RZVWMhBDjFcN0cjyj+w7n6rMhQbeOPM5G2HVAebIrSf1gUs91179zNQvNYA
mFOofKM5sLcASvOhiyfg8uESaAIUr1c688rcoXXLGlZ6CYu0QmQy8p/AFoXZ+mlA
+OKGtiXAzw9lP1M6+7O6819F1/iKXYkv5dSRaevz43LqUL7nQ0Knkl7q8Yzo0ZbL
NYM99UUX/wPoq8mjhdraKOUlP4Xg2Nat3LeycRZ61/GQIvJjWNKkiW6o0kcUS6bv
PFl7v7jM+53SCJJD6l0ldYGGxX16UdCj/+QJyM0hV9HP0e4p88vpn2ss/Jok7r2G
S69hAPYPTk6D4winRTGrzRaQCVOpUpyDZ6Pckmtale9mv/+Y2mxkCZK0U95dWVwu
ulK/rNbU12VlNXHh/SBsGNGemUG0eQK1RjFr9Khd4a+KosWgo3D2j/XaMkGWb+zV
QnEr17hyQXJFbcptJ1fgNVnij1iqmy8J7rzjdUrZ9c5CAnivG665/osObFzy7pgy
ryC4ZxqbpJWXaNgzpPmjrCt3TV5Dwe6hl30HeYC8x3CNYh1CAGobLsthOYtxqjME
7EVHm51SPykXba9p21Hmv67yi+3HmKlk2HJYewpEmpileEjPk/6W+gEMxDSux/MM
cdPWxbRB01ZqImsW6koIOhNXmme00BrA2pGo7aajs0KgS7/kBGrEKz9LfQ96TRsE
jOb2o07GDKZ4+ptp1gYT8SI2cSG/2FMaBxI3whIGMLF+QvAIzfnRkKHD5+VyODmk
PHKsBOp53BFiAF0fpTXWaqifk3nwktsukIg6fdYXETot7pbHXGzN4qPpkIwTqYQc
fYfY/6CAQFotCh6+pLVz75n3pLJTiYqLfMaq4OvLuur67OZuhhZTEwoeU+kfykY7
GNSB3dFzlppYzPAuZl1Z1vXMBmtZIUSl9KSj0VsslFgD4SJ11u+E2M8ouLPgLWFk
dUeSqAUvGVodUXuz0rJyGpcE8pKMadF9v/ytRUOwZpf+gDV4zk4kNSGIG5ZKQqSJ
xBNavz7ZjoZ6UYf1nPOhefUs0xrW1VMJGIYnwQQqZqLKKYbtmaFUjqrPx4/oR7gE
VBzKNwzzpGTQNqlDoHAA68rlVCzGsRp2tC0xrMOpsfXnIAqza/jHp0WaXViXut99
gV5XrdRj4Ih8tnsuM8Ci9WuKYMizREK+Pa6OvC+/tMY9/+cUJb9fNMhMVP8BNOwA
j2DrnP6OfmwCD1hwSLIins/Ci34Yzwmh7Bvt9VHrsqhXf+bfCLhSv8N04zev+wfm
zj8mSOa3nL3ZrM0bPwaCnU6bSxi725RujRcZijBBF9RB+t3lEVHp6ZhNQA7F9ZuA
BhnQWpMly7u+b/4beDWMJZq2YFp3/xf5st5i5SLqo26xk4iF5koaCluYTY2tc0Jw
bT0tpYm8uuRW8DxyqRlW44zKM4oK2QpZ7nCSo7ID10VlBBOfUJeRVrKClj54TjbH
rhJHc2yTJZXxXR1FBy4dCieom3aTaKIKw63/fnOijEEUxeLQyWPzf9wMZiZDto9+
8FpypH4OiVCUfDnVLoVTsVVY+4FN8qbJMW23TaC+K2g+A/5J1tWawP/GWG4lhCX5
XZOKoWgffdnadqb0jpuAIo4RkxouIiH00CEL9F+TMw3FlRzNsSxB8L5pi8BHUIm5
6zAht36IvdcyZNSXw6kuSJTAW9q8IcpMaHAIgWECqzsaiYbszC0j1VOXDW9D3i2U
0s7R1uk8N7cBZYWDCCz/4wa34HZYdxuL9VItcDpdA3NDwYfPr1kXzRX/R8nzvq24
2kg9tAJ8tfGogq7dNrnwnLhyrHhuH7dRfnuVk7v6gxSJU5ciGNfR9WtL1GgnIrAT
nfaBbUO0FhuQEKKMk/XCoNUd/jbSV4LVC5ealW7hAhTu9KFAKLe4a/ZWTpAJosv3
SNP+vE7xiabHgXrDFiKMUbeiJQJ8jpzXbiAzgdT6W1GCKT4ncMny5jV6yJguTmnH
LJOM1n55oZygq4TBwA2ynXhqv/u9M8p2cinLZS6y1xYUB63T6AAR2ypn9Ngw/z+W
qD/HfDl4y+j9eB7m0lWPSAwjXrzbUpqwxhYZtyjig72kTu94KoAkTtTpaCslVvYI
DamPGrSVGngxPngml7mBvpHaVl6F8FK40eT8l6QQwfeVHT/74SiaqxW5xOTh2+Be
MgoLmFHeUWEwrlZaIvYkn3BCZlAvcMLZQPk0J+muwb2Gue5y1KsKYzCCRvHMzJ7U
PcxC7wkVpN38bv+Esf2xoK69Tj3XUFQIHCIohd5HyqmZ86ANAzZ/b4XDdWAVQc2k
M6SXGb/zAM0JGK/xMz+QFNEwO6DSVcvI3/9Bf2JcCaBb8nY6lcfAFBXbCRwxr7FJ
ZYM90ALxGPyPfHVJSxVHxIiFQOe7eLf2xKIMMJpTnryQlaR1Oea4p2UPGM/oplUG
yoH/IAX1XT4BOtmrpJi/HzFEcN9vEdSgaCDvTST2h5WJYJP4U25gLkVdXvS8R3t/
xke2DID0O+JxrKz6/z2gDJkPkLjtnzTOsLAsjviL0UCbNohroJ4zxxPQAAdLEx/L
Jdk9mgBctyCHp+VEXgq9eolEcOgzxsxV/+oKVHSBaTLdjwxhIMZuw0pB6KlSjNM2
BXAdd5ka4zyU1Iu1q+JV6ko2ei+nYBGef2zh1PKEN7RBl1mlXfBV40rVXUj2+2am
hmm1GGqj1HCT+kXkhS5YnSAwLVvzkDjdCBEh3WtGlIFuWszVCsvpxgsWQvLLtbv0
Fed21DJyPx+KK8Xx4aZRyTSRaWtOMCX5mYCBO+urwWTZaLdDWuFblUUZgRmJVE0+
MP0tthcQIolPxJ9kXKakNXF4AtKaPqqZjtkFgCqK5YTBKHLZgylT4sLvGOkYiW5D
+jfXTONOoflDk5Ns2trIXIRtDTT0OMkarfbHmkFoEhJQGv8ptVEVNmafPbLVyrWE
CtuqbsuF8N+bKMIjvWkdVgxKNXgXSI5e5q74BpzlkEJKj/le0tKAwmUAlFGA3KEz
VixxSbMsBds5Wipj9qBP8Q4DR6Z7BwUOOKbxWMfuOQb8APOdDEpkgkqPTNbnAbUB
zz/moxihQbspw9sytC/0Dyv7WJBjX1O4hkdgYR/6RPInh8ra+1nhoBbML6vQSQ61
vK9FBBqQypE+2fjNIuIEZ2TdNA00cfQr1RfC3q+1KJMDf45vYBU5T46a/d0XcJil
mcKsZHj2xUg+9mZEULobDeYJ12FAUvlCXBDAP7XrWNDJmdIvpMHTaAEYw1uicUlq
e7tcl6p0/nBiBqlsObSviy8vueMCYicNah4XdsYFuUtPJME0SGqoQEzRZzTrqWM3
ENmbkiDk6tU88B6rU8FFBO5MtzUyGpZ6CRRsoj/ZP/Hyt0Twi1EQBTbT4PFsj1uk
+H7/d+1/6YuwwpdsCnq5wYLzwlTG97nyjV8XNrj9D3tOPhnDmga3ok+rKmJz46n+
k7RHxWlz7oo2rAVaGzbep99k67FppiRPSravxTRha7NWIHWCfvnuMHt/Fkdqwcdx
zKanCYAYEGnQ0yhE5/W7vU8fNyHZZxkV9NtWcifsORYMPGvRlRmRbKOReGTUmTHO
/p7IyyZQWEcptXcuaePSduJjImRS7lACaLImdJec4Owjz74jxYIo3IoxTnIXSxnH
y5q4+E44Lb3jP3/Jbxjh6F96sKUF//yX9FCrgeSYFT2WNUxXwdLaRxTMiim7YwHw
MFAREexheKC5uLxtH1lzslqeHkNLKhVp/74EJ/SE+1sjL0otsvCUn/7Qq5oeN/7e
dPu3FuUbm3f9Ng2jjXqcubbXn+Di4zLb0FfYFJU+xNUY6xYbv6X0GzhdxaPLaKF/
pHN8REuVkUdSVSO2ybK9+4eZIpYFXWllHmqv0wxN6g/1WlvD3YGkfvRTt1pQbkmn
Q9WX4BPoVmgnzIUb2t8G6U8vHOChBWKeCHmg0dzXRCzKcCx4sd8ZMj9z4cs5X7tr
fJrr5/jrYtV/nie9Ri3A/DrPqghoHFpL0st23HUfbI4sNra/Qc0ZE45ydCrBO6PT
H3qkfDAH2pF5a2m/Q+7i/HYIgq70ku3LiUA33+Scuf6fwaruqqHLPf3xSr1eAjHm
9XnARplTg4ayrbOJ3HI/obG64sJ/+lozXupXBpsFLFLWoZnSutgzp0H8XKE2YRJr
aekrhZ6MFx9P+qWjR1zOpXPTDA+o20ltXX/S4F+YjxuJS1hBT/HtlbeD4GCkM+If
CavM2fiof/UhwPmKzKN8AlVN8LBaQNQimbxy/ahgUr6RT1+KOrBWIjY0oZy3LTB9
gfAWsk9BAXGA7ITpwPePt6KOSMzwJ3FWta6xLINjDyOw+G7jr7UFbnxjMfa3Hx0l
W/3JA/db7Tt/oBFVqceRdNGRZpN/PFt3MzuMgMtAOZxnZxyApOtERN0kBRnQNKYB
esjAMLHDXcRLbyJ/6maCvFwZd5WdRTxyKviIPn3pilMxneHS+Yhwtyc//mtdRYFe
VC1NqKuKyIsif+LMnYz7uMzQ/qFFyimYhFMHrqxWvxQsC2cLUNW5Vd/YoUAEN7EK
BH0Vv9h2BuCBKSbIJcwYCuFvjlPNbBUFJtKfUP99nOOaMu8ne5YmvWtHNuvs5+qR
vXDlADn3Hxz6NnKIqkp2Oh8xcF4YFOGqiX7cFvQw9kFJONJ0GBQZdVBS5TlVAEjI
6kftWQrhYdqjWpcEbaDxauzZUV9EyETq/AtlfxXXIB4eYmTvk7vyYbVCenmhX07o
vnMinXw7PzUpycW+0Kl9ct74ZWDjN0Xx/aAwshzDQspWlCdfa+Q2r2ChpspZnmcy
DCPoOBwAszG/E7xTwLp7rTNDiYapo+I1ycu3jhocfzv+F6RLr1UPQsHPGaxjozUG
oxt7d3aHM+CXlSnMFnFma7XUnHRl/Px/GyoCY13B08xTlY67C3T7ICYblzOpYkoC
ZySqLSl6ctCoqlK9iMvWiS4oQI/vS0u5ArLl0rr2N1m+JETpoTpKgGiFKRf29Usr
+zRO1ULIx9bHbtDvGgaIlEatEUtT7htf5z7Nst+TjZxAmPaBg4mVzuWR9crQeDbJ
ZuBanSeKZJq8MVbNNonaar81w6NGyXBUwrrj5aRmI4vuKs6Fr5I97ppyulhHCFrp
Pi490cIQGcZH6JwB4nLuPv1MpaugdSD4iUSi7x9QEVf04eLjRJzcYMm/z/eSMON0
YL+tOGdJJ/rohg6KyfCZMe8w77fzVuyZLzDb86zCA/ecb4UWA+dG/BlhMwDRnEry
TfdkuXSa9uX6xCzrlZT8LXB+OtojWJWsM71/e0bYa78ACKZSjdsdYRgbIolgQJKS
/uNseRkqOfof5gLMZLonLjEpOeuFybyHBzcDhfzDFa5ngN5Bihu3UuBzkgiS60NP
dL/XobmAxw6E11MujA30N26iSODCTGIUzSVT5Yg3+JAxxfrQ18tnvm6dS3mdBidS
oyol6+hil6JXzyLSrW7WOeTYNXGkT3Qwah/cV9w4C9Frv3aOlROWWaBbg9eD0SQZ
KFmIcQr1r1TC2NjCSZg6pfovPEKqW0l2Rk9cYUX/FH8B/ELF1Ttd4wQchp9smokK
JqYFrcP1YTR5E2RvazD8Zxg2/NlCQ1bto/uwF7S2uL7HNdw84AT8ZC5yIwGtRv2Z
QaCA5YGRHFgt1C0Ba0lUzyc6A1ezATKJavYwwtNwEx+mu1tZGNESKez2xYTFDfpl
wTSSqk9HFngN4dBna+joFLnmM3chZIWSLvdvaS8PAYzk6x3vsyNJe8q4pfsK+g2m
bnkogfNK7QE4nPmDhL6LczYQz5gQo0cf0hkvaa2YcmikOasC8udgkMBHIjiQBZ/W
ADGgnJ3kuErHoqrBwZZ6phO+g/55tmYXEacxCR8VBL88ivQm+hl0UhGBSaulclsY
AGd2M1bSXTOPukMajcCjsMxQsZxuw/CepOZKTAT4xm2A6gLJsN3qGDif6Dy0Gqkw
9Wsa4ct/qPiHdzmkmOYNzca5F1yo5M4vGeawS6WwQtGBCkySP1XJ9dkf0zLW/d4L
sGyUjj8mi1IEEz+aXdsQgHAiR/kEBZu25tZjpbK1QWORYEDf6uvdhwSgxjrJzpGO
5UALwDcHjV31EAhJBdj3FDmZ1PfzoVOZgKHlPrZBByuoZ0yNgnMEFuL66q1xVay3
o1toA3M7vM0KyB1ss6HFt2uSClIRdnXkUGzZ9+WGhphCma6BCf2kFU/z+eZ5vwOy
Snn3TvQAhv5GZEJ0r6uCgKLe+DE+5Iq77SADGQaZei4wxXFVIABCuVbrvyE9cR5M
AuYQJp1Mu+14M93TsWtH4iRE1o2rNAoEEwMEeWf9mYjgFEriIOwr7HAGdjgriVKn
XDEQGR9D4auuEAqJPVDZCdJRXYc07I5glVWu3m35NxWOelC8LZFJ6ZjpbrFBUQDO
+cU5gaThrAavkdko5Hz0+NtNL2wLpcDr3Dr5rU6UF6mSAY5ZOm0t2RQ9rcygi7Yg
8ARPPdIcOnUXPmf8x6XFiK0jRTF7a+WgnQ60o/Ooy4deLA9wUvW7+b8F3JpuFDKd
0JYzTPmpi9XtqezosNLTvT7sRHn15x6ts8WXkjep/tnL/idWlS67ac2fOo5Gfddq
rx199LZJCxRCt76HQADk8HyNBpykOOCamBh+m37lyJ/sDFjLYBke/aRqb39t9vzJ
rJv2+YurMTAUjb578Do3L3L9BPpq4qiqDS9zLHx/R5dNy2yQXuVmwbNCg95RoPzs
9xFgxZa/3z6bV3MeKZsLb27HbiDe8p4t7wD53g69khQiBt1v0jGs93hiNI7HSK9L
J29xAe6idlQq4kZj4aXsbdq+g92fG77eDJMXiGFmvYfcZdHHGa4uWJpucWCRSDz1
5+Pb257J1homT+PIRyEu45zs0dqAIO/U3f2DB5aR1hcvuFkZMmB3xgSsKBYmMvI5
akv3rvHipLjy8d1HH2b833TKHS3yFfdU6OKfa18Vlw/qLXoVB6/IxrLmw7JuIDHe
79iYvcUMDxGQ8aMLirtWQJW7X6aeFHDTdlHm+G5TGRRCkESUykGDofa8QKbfNELf
DW7KB0X0Y/zhjsJeWgNqcEAR8jwFGhf4Vn8P7w04Jc/73tUOuGrlidAQ2VSq42qs
/mRPrnwtpGho2ZBzHCStHD1JQPfSNn/3daov0A6+qHG2WXbRb2gfg/94B0ELtBof
sIXLmQXMKObcg1pLkdiUQQcJLpPM8XQ7Y4CvAY0Tq1qV8gZiipt8XUfWYQhkZ7xx
0M22Yk5HDoNGh6Gn56tsL6woSKpwV+Aj/zzJp80uSwBDgMiSkyno/yuvnBlPB347
D0LNvZas+I2SXU6pBZ+jzENs4P4T8ClMCeCiEvM+hhdbUXJ6qMhJwBVt1vxHcRHm
od8DC+ug/NJmDZIA9FqI5nMBWCG04QaCbm3sORlzvIFQrKXd/aJzUT3PL6HWe+Kc
wGDw+bUhmdTNUWiPFtXQNGfurXvhWxlzGRctHTIoS4EjKWlrOnrNn9DrcvGfbMM9
WOiN2SIsx+2cNscwzjN8InitkzWVsyekP7qOf61N25Qr+pzsOBWCXAdFxAO/NF7X
c/tHkYB/GTIvAFf8Nl/fgTZUi4hj0m26PjDmCO8EQHgj/lIaZe67DSEMnXJSYlvQ
CCDEkj0Nv4wffsz+JOBeJcFrvdFWXPDcWxAWwCsXPtjsIKvMwx9B+HiWWKlvjKpQ
N6WGteO1LbxBSQ2ogYzwxCHlYJgxVSXmbrxRwEgb5cfSbvbJPI4OXXABGzBmgAXC
O3qlmgV7ai7T/ucq2dcjxPxSukXtqN7Je0dWMq243MuOeTA0lzpw6TmcfuCpp7TS
zpbhVknh98lDQBStVhHQwW323mipYzOhVEqrBYn/gwd/C/sh4zfNWF9CUR50yEBd
yOyw+GwlMmq88hlaBrbHkCL0ncKEwZxyaUE9JS8ociuwalG3ORQqnWnEfObx2t7u
kSnT0ej/4O9xWs5X607ZNwuoBlMbiHoHV3l+Y7zWB6k09DPb1vihjrx0KCKq11Rs
tgy8PinIaPRwaVW4/nAhSSU84hGygx+yJNY45m6KzbfRNi0fOEnhrIsXE718WjCm
XTEqkCIRCEzbBts1HQ9uV0VFJynqddL77/3mAtwIpSdGOVmsiOzMLJpSa/gRiazW
PpkJpYdM2WbX85Q2tkqPFPswwrkVvs1Z5dTFk3N4VEG/Yd/TMoQ5DZGAvQZ068/b
UF9b/hZR0L2+PyV/ynIpe3zSy5rVzpEiPxHBi2cPur+na74M1WSRSylGk03yhklw
JE62KnziW4rTh02g+tshXiOFfgFTNp1TZjT2U363h4GMrms2Oe0VuekZyvv0r4+5
FfHGKAalOyQ/YjwBuHdga/pazdIH80pZUQsWSYQ7KfeZ4q2c5NMv+X9S2dd6BPhC
800gmT3tHKKFiXRsZsInsOCWiF5bzf41Smpv/bsfHbLGWbfwDKpNMGodzuKIHY4f
QcNzL5QBokCyiTBM4mO2tucajZBLdciMjICC5EsoLoJdLWlRLpJgoFfeNO0CO5oz
dWzBr+IkEpSJ0Hu1fPgrmHWSS1fWpD8n7FJNzqdquFL1xxvBpuKMAK5oSrxpBLlx
Ds/9mgVyr66sjRPwv4MyhLAIUd2ilPhBcm0lS3iNtWpjnEhVXe/6wsdLF3EJP9Fc
bB9VE5cJpE8PS2B+qWSgEzYRAYS+7/2iG1OmnDPfv7nb3hKJxGGl8HmtE0IedzXH
Hew/RuMNPdDRxCvXxuc4FqekaMUlgan1HHDD9Us6H3BzoHtF0EM9ha9MJJr/qeUh
IuH3lMJvTjIqZXaKvySfO7u8vR4JR0jAVp9bGuYSFB1LGGJUYBOWbYOQRh3hGace
z4ZGqB39eSpytAn8DyQPJTn6I99fHDDLrl+EgY9eluDsl77wz3v0sHcQ1RY1u+F5
c3AZ+EctJYXJbOMaxbIuIb9np2iz/bmuEH0M2yrejaJy/hxOmmZBFMNEjxX5JLn4
zZhrB2vO0bpoi0Ctdv99FOUo1hP10nmV4A/12vEiD24yAqKI9RxcfxgJP7EiL7Ie
COQWzTltNy0lHH7mTQ7PURL9v62v8qhsOPKXXdLFnvgQ+PjuH4CcCgUgpsN71qFC
suLHNnM7Jrrt5SBkvLL8GVQ1cTwRBgcpMvOUw+HjuW6bIXAPXhm7kaHUXxsz57Rh
Awp7ytDXaqNbvvj6vsJVqsdPUsIUtvv5L/vyeU39Hg+PHGmfI8rAljhfAfGK0r8Q
cJHuUwAMUH1fWGtAGj7QTVnbtqaBFlJCMKBUHVYEpdX4NeGm/gvp3HwIWK1bvUl1
zf0iNhZc9JACRbB+FjtuPif+lD0oCnFmH/nost4Ioe0aLxYv53phWttcIpltTnqp
hN1Us66gYP2/8jzr+pcfA0OSvumdWfLBtHDPAgpADVMwgfTRCnVLX0ukcgfrgoiL
hNxyUkdH5Kv4X1Y7AtLFDqIhreqM5m2Y9JZisQdkG41wjmoV+n7saC1Q7jnfq5mx
1+/vvaanJ3Nx6JTUuiz6m2p8pA2MMa8EM/y3MRdmKloFFHMXR0B5c+KlICl91jB5
Ph4Ws6gHgUz4d+lMEYx0w8y3n/4yfG/ccycq06Dp/Wb+mqf9qPZ5e6YcqnyelhoW
hoYwwlN+9Qe/0cJIfx0k8+xifpTZT+jy8fYuZJLO1M2u7xpMkNkDdwHFFoUXOojL
aSfx5rePqLubp5bnnZ/MKuKc3K360Ctf6YvOpVzkIzlTb3rRZm5nwju9f+s++PSc
dnzcD82x55QVrbUBnxA3/1FFkIdnxthV01Q4SFTdvEdcD6efI5KpPjgRP1NksIIC
tYdNQ2gFmkwcMJGhNq1Y1GMsF45FTQ1wWa6xW99zxnwd8HoZyiJt/W1Qt3mL6ruE
WK9GiAUPq8kkAkFyT9qX3e+l3Ve7xT+cAefmSvHVv6C4cnIAS4n7tCdIflo+039u
T67c0LxSNS/yS66EyIcmBYMO+RyngHcYRiYvqTIb+sIVNit91MI/IZJEFVBpQq3i
Eit+EELMn7TAMY2CDaRzbvC3o7hX2JoCnarQCsDYfSS7qj9XryQIefodF4VhPWIS
xiQQvAxfWdcITz9mXDUwR/X5yVh2xIqV+w2gDs/rV2ED9l3QXvo4F2rAmevEtMH7
ZKbsFzLcdWbe45pMri444Nn4DPZs3Ks66P9E+1O3S/sReIp+oN6mPhNG0Ea/vT2O
7QRD5Fuu0+riWgo0a3ZVh8aJVkk3wpb4SusO+XFxlNYZHyZJArTNskW5KsBUbzh8
qdvEtBa6kXEEOWPEh6y+18COW1BvXKczx2UOlseKXBHMuduS4zTsmxNl2GB55qyc
QQTm+A+75uD2OaNReq5J9yF7b4KDz1Dg6CQsTmPomwMar0IEb1GBuJPTfAiAk4A9
sDAYrHvJRJ+6Q6IXRuZV5QyKBU3gUfr0vcnO+hcI4Exm/slX1a90830vGvXOxIko
snVc9MketkycONwRMMiFE7Jzxu5Ky2pW803FRhvRywgf3T/JuQCd+bhA1MAVjCw1
DvV7tENvpkrpaL24ig6W7HwE7FX8wGVkAYtGkvEsUHkMPlLFTa9MILp9lrOPCrLQ
kB/TUaMNFiZPv3Jns4tn3U0NO6x5T8C5HVhCo1Yyq+E5A16a2WW7OO+1ZXI2p+gK
tsoN1JvTO3TgUpJRO8IPBBmVBeHCFurNvKjFwER3jrUMrLmEoI7iI8TuBX9A6p+T
jrxlERxWkcGntJEA++53k6DpUnFYhrG45HROKp/JTghX93UgImE+MaY1Encmr1ZO
WVnmTls3h9zHFHWJ/a0xAwWs6DCcMqBlBp6G8T6HmGwzKofEPxELt0yjIwyuNoTI
Gcbz8p9Y/g8UEhe+2oXwpoBnvVBkdCGwB1gOUZrCp/wotaVJtmc2+dkiDhVgX5tk
ajy8t+BvQB4fc3jV8LeBAiKM597j/v2UJiljvdYaAYJWvMxAY/bMPXt2LSTQaIOM
w9N6W2rm25mWAg0+Mx3wF5dSkCvq/NWrCdIU1uIT3JjvalrIAn4po/JKuEQfY7Wg
0CFYMdfdp0VFTQ6JEw2ruP/FGGJte63CF//8+oCfkWiqZDlb4O/MGyQ4/xp4hrub
kITfPjT1yxu05Qk8Y3MMzIrRJ66Yj1FKNKLNGQPiTB/qOZUCDA1qPOJLTs/zCUfX
rao7Yl0PQoJIdohMHaUcQUlsvtwvn0Nuz/4zIRtLNJzeC284v6GClqbb67cP7s19
RjlacyLVL8S7wT4i9Y7xNVSTUFUeLFLCu9DqnuXlnft3pktMHbmqvxiVyLJEKLDs
lD09y4QIfTwU5DdAbpaPwTrtaQJX02r3HZZ2deNuZXlCpvN9hw/j+gm74OMg8qfp
FvPoPhNZzqWEI2qD5oJRr+NXy9P9006WHMXieIYYHk3yRtzoZAkTDlSbtJW9BmWe
D9SQ45d1o/E+0SF4QaBFV/9soR9LF8X9AgiMscXkxKJoxyplhW+MZ2qJiEfNc/Ab
U14yRpXzwUax55gMp6Wrt/cZYAllD/2tfM+2xdCQQHoseFjZqeS8l/2uttEq3Pyg
VqhPhVSb1BImU8RVqYlXEizsR6+AN3jbPqftlr3ZBjw+HbzM3qpgXFWmOncN+b9M
ZUoc3P5mso/f9HDXVK6LUeQwCLlGWY19gJ4F4qTlAHqZ8nkmVzpIbSamIEHNVeg/
02SXPakm3Fd2+74aAMcRreg5XA5n3K3Q7V0lYgHoEqSg2PKGs05kHY5Zos+fb37r
RgYQ0gW+QinHUObU9a1DdgZ3PuqO/2fEbizK4bpT5A8494tBqLj66VwBScs/aAx5
3K0yilp39y8wRZTHeFewv64OpL6r0Q1KQe8PvLhdDmjbpaz0ib3bDPNCVHh/aTBC
cK0Duk1AMUE+4Z9jhZ2feMlR8nbDeeiQWtzCe03Enexyr7enPru5JzREGcQ5ks/6
cW037AUwnjeW3eml8STLHIRgKSU+TqyfAoxFDyvkXu0YPy+5dyXZzRiMz/gXvq+L
H9wJej9mXbpOO94axDLAPu2iLpoMxfk1fka6+smqgBZmmZ6gQjgH+3TztvhKCleL
hAzuR6itVe3RSUKTKrSL9G5ZAdTmE7Cxzaey5uKz3jy5UB34JucKeYrmo+e/linx
jZzUqIyy8aG5WDOPcaufwk5iuD1R81w3n/uhUba++dE4MfbJP0gSXdeNsLzth/GH
30IcO6HK9JqZRpRRraw/2q21853/zm/9Q2K+dpPH/Ny7JpjYmEYSPW6Wd0n7SH64
Ijvs6nXhTopMRbzbcNYlzrY1gMGsdVrOJHWATeayP/ikxn2HG8IA5haQafwWJfxG
9qMbyNkZOoIFycq01DDKI3fZ/HsF61LYd/ayQqKH0KydmCkk0LNHxlL0GrqjN3/P
2Lfm9p9Mq6oy1RjyOUDsl1PKYKRWgjdGbvAC2nTjs4eHjh1dX+1fRJVuSWGshQyW
U63h+bSOJbSk0YClcFQI3gtqQ6igGyGcvUH0e2HQep7ZCuhgfa2alKKN+SdsvxXS
DG9GFpVSmj61+3aWADrvXRlbWNhVqElqmAQ4ELnH2I57Jd+53a90JJSZBjciSf/B
lDwAffwmiZ1PITSk//I2ecwFEW/ZcFJp3+GntMSF20UxEXviiQWGCZVC56qwxbN1
4s08Fyb2Eqg8e+WINpyQ6gLSOKesYuxX33ozINy9pwNc9RlFg93ss/iB9ZJqZGkT
uBl2CEEedhiR6FBnktNTFR4fbVaV8Ib6w3eLzK/cN6h4sbBaCrRyAtLKxqhNluRv
p/LpAK4p6ysbPMGNohWPtTJ4+65wFmMAvyIt5Un6GHsr99FwdA+gv9/j0EhrgmrZ
qjsq1CzdB3DkooV2/jgjGn0p1X0PSFqeCPSUcSgj6kT25TVoDap0lZPZJm5LRe/e
+qL3gR7kazt6xHpztiKzwcfLpLVRfRZcBk28HZPv+wGfxb9Pt/0Z9jQQN2wKszQR
JnPF7xDrnCrumqssP6zmTz7wy9X6mk30CO83OFFULVAdLds9r5uWmk2pVXarJ+ge
S1HTuyv1Hs056PsS2XLXBB24L/vcDUbyMF9jHCUYUj0EwFOXPigRXQQ/q91zceyF
ihqPot+RD+UrlNdeb1cNdJ7dK32Ezl08Xi9O+H0N7TU5oV0EX9Pj613OIFq+tSgM
eh3OBvrINVWee6Rv/XuVsa3ye52Y2FEf5a96ZpLSCdvVpBx4d/XUpybuNnhDjtWV
Uhziz9Q8vBr/rRffsvPXEVOBqGjSqbgFayJWVcLSxYQFYM/AcGF6cch1nhEOIlIV
h2TDZZuthMvDFViZYotfxPwwiceDs9rCvRi8KkwmRuHhDc0eoyGeSRNyHk5SFU8q
cYog7VogRvLsyRpxTksg+bWCI7yv9s53YLLdFns71Nj4DrAk3VJcrldxXCha6MWi
9xolQPIGOHQ2PSCyxQ37Lt+ztrYSeDGnttjIjSAq/GcJyAjbZ+9dS9u0NBMANwLS
spyqi6AAsX95tYa3leLvNrYudkVWh7OBz77rpMStKxPQCjFiPxEnLFGBaB6/y5gd
tswyjACEujZtllZO5WwSAo0I+gI7WJaBJhep5Im6wwrwmHWSkZ/NxV6NdBlMOsxh
nQTWrkpxkTeZr2WgXZllfXDIr1H8jotgTU40DNjU4CpIxdJ4Ph5+00ZemE4pWLD+
jquhJfeKDuE0IESqs/F7+QlqducRdsWopGO0MZF7heji8yEv1X/S9hoxw9e15IS8
KL4GzHJwUOF9B3CJwoAcjj1GBpw3HeXRBzPcm4UoV8UYwIbhp48hQmr2tUSrzYDJ
QdY8czoF1nLs6AYvECnNgyFhqOSNVEk/vVG3aPNa971YB80uBvjRbg5CgKxEplaJ
3X/tSe/lC0IOrpFO+jwOEhvuBrnNbTvPT3JCGtKtZrlCQjzXu5lU8yrKqqttRsIZ
Tw4D6k2EEUWkJd53A0RCbwiSAFF0wS3BdGkb+WS9703DXfMjaSBtFtPSyus5MZLx
VV4Sep3pMGmMwiYZUirqBgFzv+m76B5R4QuOz7pd7MyEQMTBuQwbCC1Jy0v5BhL+
sP/YCs7b4wumJ3g2Rcs4k70EpxLr+hwuBeTYfDL5hqYWBD1pi5k6r+p10lFnHEH2
cHJ3HPdusAy9YdjdQW+sSvcbt/yYc8ldqIE2MjGt9D9o4J29cOpXszZgljs7eLYm
7M/jUfuWdEsd+5PS28w7mc/4fYwijRIe63CJMJ4qy1+URQQbs2z4i6CZyVIlCfa/
dnGlnxJAhvK3eJ+HX3XDRZRtnGl+InDcEF1F18bwH5OGvFp3KYluY0KPLVnakiyn
v6unigjq+01d93BFlq1hERHLaeSIHfmcQYMZ+GaDDOoW2mEd4bb1y/AL4DzIHQVm
LisKIg0QuC97mMClqa4ACCsWD/LVlE8KvXFtCdsG8SAn8qf7pw5dBnxQWbA+0tG5
I+ZSbWkOngN54O7apbB+SSuRuHrutTX/bCGo8mPHYKdO7Dra1wD91c/q5XhRJMK6
sDnKpsBGfRDbxNIauXkNe9y+2d8C3MT9RB45GPVnUQ+XAF6S0b7xZNHVowsM9z5d
cBFg5lCYNb4RGfWargnOW+s0x9b1SGiPWhbHupE40LKsJX5BxoQDhGTgBWFlQH2X
F7gSDLGmU4WzyfYVRhi93R5GpBcT3vHQcelBFz41wcgA5aA5wV+H6Q2v+m3xYhZj
tCsVRlUhz5f5Y+s+ece0yWP90JcZZ+CwiRrFjRvUfk1Svc4pN7Z7jexej7RFP4Db
N3UzWnM8J11EstRcUeXjp5YndohLejZvEJVZnSG44tGxe1evEfTE+aLNcuzVpIMQ
Ytkk4Dr5QPuUHURjj1ddVvX6O8DUirlERt11j1tebJEUGiw2M33kVYU5IaiqHvFi
nBjXNiGItRdCc3Mn4DuHU+wqzRINkrCq+FrIYTrAfX38QiI+7riAYt64BKbIG6QG
u902jU4CrbOd6b4/b46Vt5nPmatq2C9/dcY5SDeUTSQIOZ9vlf0F6f67JRQ+dlnE
E6Z4M+21n7aAtd0aEW4d/XA1MRmwxm2tI7zWMTtg8pn5ZZj41YK1YOwvNUAVaph2
16uWqtWD4bQ1HZlsb+VYUksQ1MIP7ET28stJtNyqcTxsW/gHSjUe/2IzB+NTLbN9
GnRzJcCaGlCQGmwYSM0090lcBNsokJ98xJHCY1NyveTNuT04QIqjLAT/PR9HuJ5e
sJHdivcpoyNs5yqhn3bf87GBkGTmlduiuAXAIZ2aPdklDyL0DU+VnxiPzu4jva9m
/xxDk74D1UZ0lCFgI+fzEsl0j0CdpfTVl7hAciM9ylQCQmWZ2gNMpUlbWhmn4tqK
wBEa9wwZOmvEfGLamO+qhiefrF3NgJ/XK6m/UKuSbZjZ0UjmJR0DypHtPErTdfhP
7KUpsiK8QLRwzH5rX+9ZU1XQAbrBTm0g8ONEhzurB94qJQ4BeMdPdylWJ8KTmU0G
tGU9F9z+MMTQYwPFaVV+mhCklXLpFM4K1leSRjOO4Q9Z/vZQ+F6gskuhqPb5+NWt
LDmtOPvYA8sw1XYl2qUWb4ELWC7qWyBYgdETlLefkgXdFddHAgkFFoKnpz2t4cSm
ad0Exr35IHNZPoH4L4XBeBI8OL89LbiQnASZ714OEsFl+UKTlZxeur3gX1O8SwDJ
qCYc0DjTcGAJbAsSea5SSkt0us6/J+VJVdubIB5oFXGUn+uqZK+mEvsbdzkVA1JX
zb9czpWqLIMf9gbj1aSCh8oOcOrOnZN3sZQKOyXfHwQyQGQDVUsjNrLwoXpWPpCR
ksgJ1OfrEjo6C6OoouVtmTMdZPc+6XWVnBmzXzyoj+76mDMFjmUT4KeIZjs8gKpi
MYfeKz2WLijdI8Dt5NNPislDjjxqV2Si3eYMNIqkWlGcGIMXfQ5NKpn4fIpaco3F
ya1F5rLFEwQ5HIzkj76jzj4fIWeZx/LyIXMgROyf+qlV6KW6oAzydNJnEqBqDPj5
d7qsqNUhTzETHNpRMCc0NQM137LloOr0OQca7TRzmvrgYwoKq6p8Zg5qG8y4KGMi
mrWOTLMzr43fgon8vYO32dJ7Hig19fgmgMhkql1E1S8y8GW/MUaeQwlwZ5i+c+gh
SIKDJm+Y+GBZG4H1jejNbfKMJEWigRd4FS5LkB+5bEWl6SpadBi+p1QRADprOPJ5
g/9q6eRTTXaDzSrtgcXbsXrjsJTrLnjPrBEw0lxlrxnm0LwdpF/Ica/2r18MRlTm
aIutZ6bKD57ijrPHefrlHYHDgemtxEe5YFSPvnDsrrhuuZNMcxBWPrQDEpA5pRR6
cIsI+eMD4uWCyazB+BRa+N7l4DTbFDM3o6h/FQS+x8/uyp4EKQrx71fM1/c2qTkR
yOs7j9R0kqZ1jNwnlOER10Mit/0Vh7r7yYpQAu0YE51pG4+BZv6f52ephCya1QKI
aesJW5WaEmogftRL5fzgC71u8hmQiphO52bnaXEuQdf0CDyFsVtnODCJ14YRnroK
idNulLhlbu03sZSR62GnSwz3gNh9irCmcT9jiN+qbf6oUcOhR+H/JJlq6Khz1cE2
xA7Gl/6rDLZUk52nSMQ6mKPfYv/1o3VH0qfSxOoH9qw8v3mgQPBbX7uZA4z2wjCz
X3WgZW/3kyEoc2IVeEjW3YLhGQr/AwXCzUuIsIfv06DyHquutT7YDb1fjB2LaW77
dTZadGQbeEeOMesvukY9214il6I/vb9qPs+BOaYw7Pn4FhFvuCMO0XUuimtvscxK
SGcJocpQJqXNs+biX8TRJALhUoVfxBUAgiy7kOYkw0+SRNi+LYUAoRE5CoksN83f
OrSBveLZ+5D1T7HemKsMS/Es9T169GjnihNNOYlHpAv9m0i+z0CVHqsoLtidqn9I
bCdTroa6syMZKu8nGku+OglEPhJ3M2IqEHwfl6EMvFMS+PJuj5r1ZvzHsmdh4oY+
tshqTg1GU9MzqDpPalYFsjGq2qi30IdcwM/BDVlTepkuSM8qdZNqwYh8SuSnXUI8
1WDFrbJ9C8yGK7j/WJHGLoHWNSHJoI6MdQTG4u2kd+nxhZdyKi8nIZY2L6EywUTf
JVdsZyBM/Qhi1/MncOdi5JKKAiWRvH1na2BE+JRqbaJh2EV4kRgARp+9XfXfowp3
MHI+6fzQ4EzmQzqup2SDUpncIv6VPj3PUJFITOwUIz2iRnM3rvGlgXR1pq7Beqno
60eLSJYJhWuerxEyN9H8doYpMTz81zcHAMo3Uvq8HYeZe3Fkx1tYPCFKOE8UzVBT
Vl1ppJmE6pSWx7RhiaELulYAlOiYfBz7VLgqw+YZ2hCm5vf5Hq3+UWe2ZfluDXWn
HG86Av2Z74Mj456tn3bdlL2AUA0tJCYlWcGNzDd0rrTVwKZDkRvcuOAxJa7IQ2c7
f9XS9HxNUqRONBMkCX1eeyNMcl1a++v3Kw6IhvH3ZE9pyPxMjxO6HrwoElSLYosE
ZSVuW0NLnldxn9vphJ0LHq7mhaYwhufWRv7Ty+Oz/L7Q1ab+6I3WJSVqH+4PSyD5
AawIif7paPXRKBVGSLxIARCbIxFgs8TkG/Cg+6nBiAF4yCIthhXRemksN0UzpcVV
bOSqajml6oMvIO9myxXhwbYM/H3l6r5ISwAtfhhBrKHNr5WHr+T8lZ7ppWtKKXvh
R32qwTcGqi85k8pXOnw5cwXDyeQjs6sE1YDLfZsDvJWxJonOqTsqY9RBxdI61Al8
PV+HZGmNnMvQvdf4tM/eriJms7KuX2OW/wsxfwf0LGiMP100cvySwmMG501cCrNj
d5ZMHVQmJhXjc/s73pPRVLG7wxOzNAovmmGUbI1dLQGhVmTSA244GLv4eAhXm48O
w52K7H+GZe5vCLq+sigyZS4LhS/SzlHd8uATRO8yCYyBN49i3XUKoqHSTKbtybTs
y3uq8kUkZVm5Ujq6cXLVuZRT6T8RkY82dmVA0TEQA/6dr8vhEkaCKVd00ArmDi7l
DhLwTZlbEUzPuP0fnIX+iqdb8C2SwoUzreIn1kEDeh/qCd005UHicuTpP3fN4iBi
6b80rDlgSS4VxQlZh4GB+l/qdYXOXU5E5FxVnEB2TNYNwZ+gPYRqhnLn0n0kHHCC
rBLY/tmvUv+6NtJOq+GOOtRG4797XtdcM5Y0+T/EgD/KGf9nwx6PppUDNNCRJc6k
rItbuJZSgepDu+RgYL0DQlSJ19Z3Y/+YxgeTpQby4PVjcyebfQbpfc5UvhLFtWTz
Dn2De13Jj+T0uSt/QLD2W3YRnCvyj4JhTJIAevpWKzcfEiz6L/gQaFZJysiXvuYZ
sY4Ccq54u0ZxvMXyTCqKWFKYQIX+Za8ktKpVvhxVb2xoVl1jFDvnDOl3WsetAtfa
0A46w7zEcR5hWT90lN8hIfxtcdCMBxWbE5CJ91aenEvIoY7UILcPdX3XpXH8Yop+
aBx5ZBF8j3P/MV/nR7JhMMExAyoP7pE8KXl3j8nrwbnsYu8xvd4ndRTKBBPbz3rt
AuZiztwufBCxr+boQcqr2pFymSJWCUSllUB/fU1rxxYbjZbAi8SKQKk2wQCqId/Y
ST4UvfjwjTLydlmID9To4XAcdCIj5WKQzAz4kpxkD4Lrx59EfS9SDS6mInNhhACq
J+jMcEe5dVKSy+zr/Y6kK2KEoEwF91OlKGVaC3Y8ihl+3wpNPs0jawJ0U6ED6rd+
srkBX1vsATf+fVtApOyqRdHtTR9aC4YcHOjlZ+F7t7gGaQdKJN704L8jUdGSJ1i0
xySa34HIhKaEHqdQsHx8GKMV5I7SvtcCJ6n+U66GED73APgtx8wcQUHQpY/8rDOl
n3vcolQD0Ni0Vk8b8kpOEviQBoJK5Z2hk2+Fpk1xv6pfV1n8KD/vcY7VhySsMVfQ
1sxO+b25Rt35T/K2xI7LlWx1OimpKaZkSXSuhiYkyEB0c00YQaquJNXijhO71/Nh
wlgtfnuXZUsrpZYuUCiow5bSK3kJTOs9gRs0ot7rkxwoIoKMaVgQRvNtm7SnNMws
MH2l0zBWXk0XNNBWb0Se75NtBuml0hByyvkC+ur4OuL7yF3zvx34LWLVL4zZ9NXJ
2rxikAjLQ34My6mvpA3vyDRBK1T4j5wQPR9v+bDVdcvHueDZ+l2Ws+xJR8aP+WMG
jRbpva6ZgPcaVA3ecZ8xdmN1Zey+VcLKumcV4OTgwZfDfNfRHOt6wNEoAwrM/DX9
GhHeZ0dqZejsrDVv3078A1Uk7L6rcg5pZUsXot3nZp4OQpzOC0IKyvDuxprO1tl5
wlTmdYIs0QC26ciCbRazpiuPOw9U285LeRxwt8tPKFePFJaK2OqYqkx3EBX0zng1
+pHXwtoUeuj8lVBCgkGlpppB3k34jhgokqp3PlBiga1+RfIK4x+00QAiqiioACyN
vpHu1fsTb2LThPu8PTVaX7bgfw0/P4RH7hElz+sQcjWrZTaniUI1UxkGP+41YIfh
CA2U2EKWm0wVZ1zWhA48VEdE7yyJpfFH/oa3fd4Dfr14G9od9lGlbKHdFF/GwDcw
H/gADpsay37j3qtuU1TLf+3yb5IRihfeAf8CP7tMwKv//ANYFsOjgNOMOgKwaTb4
SQkHI0rxbEFOzCh/ANmnUoGkTz9Qr7rqcf+QEid4ejevPNuOQTl9My2aCLSpdRlx
uWB4p+YuD5DU6pWnaocUj2a70WMdiUwFyOqqyQJKzQXDXJ+aySpIOX7Rvr0zoX9j
l17ek5WKFDlmoiPX+u4bF8Osiuh3ytipL1TnN5wFJtsiJRQz3LyDrAexd8WBU2R+
kCD/NzM5I4k+r7FyC1sEcQIXaNuEpg2coESIRaZM6HRxbPNGfSD85wXOa+g7ISy0
3lg5LVGGpK1tfDreroPjXyChohSrcpJ1TJ8iVSDiPFs5eLx86wt1Jt0SV+5Bfktr
eu/t6D2DfL6NHYZlWrV+pJejDXDEb8r2FEPNEZISmLYs7WgnfiAVMcwseyz08c7k
K4A1jcCmWVbKNtGcMMMdtZ+lefk8oce4u/YomEHZAqj29gf0ME3/KA9Ez2IHeK3F
UKgSnPdzgnHCAtrtno2OtaG5usEd0y3nbSw8kBz8m4UKPEW1Wi95uJtU72D8HrAv
u30nR0Jz/SB26g1GM781HIjRd/GMUaZ8Yw4PBR4Lczg7RLhCIstu/+vQJBb9YIo/
cvc1+vZWe8kmJdxI2lQfzkYE3bx4gnQWvani7mwt377VM+9xKmyScFtWT/MeP5GI
DP6o+Bss4lXWLGwqVgAxXy4o3LhhjaaxKe3MkxL3cqtJ1fF57J1f3NgYdVg0FJKq
JK0CD7GboUOOdEcgCBU/uGGBw5mg+FoYu0+K2bQjXgZqpRFESLPfqToiqhFuMx0Q
mdLlDc90q2h85h4I0n9KQwUK/d1NoU7rcq4iZVIPu0zd4vyo6sGOZQKa+tA48ip8
3G/J6/VIsFZrAzu9nyeFhe/gc8G5fASARlzsRQO6dQmCUTC0yVoK+cMYD+K91z+y
mHkpajsUnITwQYT1zbxNMQ==
`protect end_protected