`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
ESp8jRyPtsiY+Gb1bQiTII2Q/A2TYHPRTGJoFFqyQM7XLnDwPbBrylQWbGUsrPBA
muBITz5G+6VxhpksMRPxEOLg6dlg4i1mEtmbSodR32sUhMDfgq0u1H9+o1mWLW8f
AbKEiBNy6A6pImqqMU3ankWFyVCSDE84MlOqUn1rhzFH5zagc9NZiE3Boax83Pnt
PIR+mST7FdMzl0yDzXfG4dmNOrNL7gAUUKKYEgRRdcyZLjkNeQ0dAmL036k9pwp8
jiEZb8z0piRluJCMdhGKQsoKpOO4qzgHqS6nNjmuut1cXDuO74dh+4cMFG1IcFQO
6ogffBewW4dZBqvgCIEQHLqZbZIlJxQt7lM1+/SJbHVzPi2TqQ1IzCHU/3vg7f/Y
p3tnLucmprIBiiDkkpqkOG7f3m3/bl6Q1TIUNGX6CoTXQAiYn8AGPKrqyY4vXP7u
U3u2/B0r0KWhi0KKwVtrbZwUGk24hl7rhLE0gAmiS8CwnJMAjUGqmEDFSM2D/CFb
oR4SHNjiy44AN02BxLdn3TUr31DA2foQIveHqOl/JkULR4OMI6UWKoIEpX8fLSTW
jOcPqvO9thKn0bJuk6tM0Wiq30MD/SFN3x95iFcox2/ntNkV2G1XzzM8vI/vqo/g
ExnK799ykUO40n9U4HJKPZ4P3Atc0cMz4g49hH9JwOlUnTsoNqbyoZ8iu9J+M6W2
XbYn07vIilMhgJWsGkGwGUJTzzc7O3Q3qCiXwZRQSWtLb0UyyJUy+QWvAGsfVyR5
ELHK4rqeUfo01zdtm6WXvSfkFPN+NLtEWnmQBhIVi13Cd0Lk7aF1vKDEEHo4HY9G
6/akH98h+QXQNDCbjhR80Nz3mXWsf28amh0VcrRz5YFTu6Dt6Li7hHaD1ASu5jNs
/uVPkQPLY1qF3CSTis2gTfZsTCyWIIlUGKUHtSQ8j619yrRv2m8HdQVy5XPsnuBb
oG0JLjjGv27QNwgqqnn0mepJjWwzkBjL+7whhwsvDKf8/ws5BAxAoBwounjPuztd
/ga6SqJDJhEZg/ArN36Ae9fiuuWNpshxh+pRVUT2U6mnLFmriJ4kewDbbYfetDzJ
N8qTkJZ8ntJcxs//vGT10bMueGg4EksPrc+Qf91oCY4upv5Y6LLtXAAWjyaueBln
3JvyK8Tkp1FkmiwauVeCU5WTt3fgJWpjKldbv6HN6gw9gYDO1Jz4ggcCNUya7F4t
h+wkY5kZjPaB4nfMW863k6asbFrBiAZBqhk8Pa/V6BAaiJP9++Na01YzmOQJefIQ
edsMRU8mkxPy9vh8Vy0ZrUG+D/j7cmQ5nEmJowyNmgHqkGJSdDVvA7ric+YgSrkP
7w4gmTikWismSoZmS3mWRA1AdiscvICgZ9Yc9sfT1vfuKGImsQBTKGmUd45h4jB9
wuVOPsZuL531IECiTNEjfRunQss9br1Z/gBTDfy9TsWEhx7/fsH7l+NxrkFj7D7x
CPAZzeGLDDSAo9NcHHEJbNvLkvBRJqZfBP2lWrpnTh6CaSdw3NlEmmpLySMkYLbD
rl9yB21cqkAtyKYe+63+KbjJV0cU0Aybw1i4VVOLduDVGNP95gUx20gFvrV6BYB3
/BZhcx/gTuX+YjY33eY6Cmywa9jT2aS0nxU4vzVvAXk1kVfih3+VRQMae+QMFnf/
v3MatS0DypuLUfUd/URv2ueFhYgCADGLwOq/sI4nzZd3Zjq8PJjlhGshtDdaQSfP
053D2kEmrn9pCZbknXzQC1SWf+V4+BX8yidwlkYIFuEpmgurVXApbM2z4waNKgca
7to+0ubHL1hhh1H3qAWB9yuQhcez79M8i7e6xKQylGp/uyLMmPNsmfuVvyF6/1O7
34OCn6qpf6kqjGuct+pM+BQMcYSWKK98nQ7fwUe3bSVPJmuAoL2P+pB/YLKA+RwO
cu5uOlhOgwjvZKo+Lm5dMGCrqCK6KVckERPMIjhu5HiPzrMJAZxhnP4rPugpJKfp
MtLhP4IDQ9PdD5D37WswvHKvzdO3dbXHPiEVkOEwA0edoC1w9z1ry7g0WObfM+sN
38evmoujQ3ipVqqIfod18tWkOxddsVBzpjy19VNPgQQkHV9TSP9GaKeW19nwrUXB
chCbU5SSyIkg4r8zRqegBhJ/vzZfKqRmRQMWYL0TTJh3StAGDVJrK3qLbildCfUl
0xI3bJUa0/UsdQfed52inhQ+cVTF5cvuQLKYTQlDRcMZLIQpUOgKv5qZMKIn+TpP
Dlkoan1y2kXKNTYYpcAWV4wPp9k62I4MHuYpaLd4M/5WsdJoYOzQ7P6e3f8lMqji
aQqoUIGH7BWHzhpV2PfDsHQt6oTf+laLcxijozfwdxqVaaZTqeeoYzAuIbBU8I4m
OEvQniYJ4j5oss5LZPc9XQ3jWrfOjVUSw/nfdih1YMsOtaHHXG6wZD1AZIvL5lu8
kqfVpMtNh/M3fL3QGZqHikotc4PQy2TkyTMU+M7Mv09hQCLF7Taima8c/8Soq3zF
WxeLjXa3AJry73CnmEpS0RljD7j8fsCHd19lFGmyT027Em1PjiBAbwv39oZ9LLtV
9SL8bQDsDeC9+rz/7LEdLIMcFJ35VYZbZUwjG5hogcCE/M3qJTSxHIPIpa5/+0a0
gZOeDERmUTrFAoyq4DormmcBKvxnKzrRPceE7EYxv8xVyqFXlNqSa41nMU0cqrvu
5WPvM/lryccoBjApipSCDRjXGyt4YIQw+GUSNXZeUh9aEowYtiWaNbSSmyau6hjq
i08oMYDF4UWTfUtexABNoUWYbtu3YidYT7WYbRlQgQEXlfl1mYDM+FYevcoLksbU
IJBu5ZBgRGhT45Onj2c5ZmeqD1AflNsKzAlIXto1HOY85RODiEMXK/0Q18SZU+xM
99dSKDPDNJqVDxypQFU8P4tMl8F/ESJ6BojXYO56d3qoc2f2Biy1O1//lSz59WgG
4vBSoedDEwR3gEeSK7nPqwuc3n9chdTAdxJpGqjg9zz6dQgxwMt3C8V15xTEyXNV
SDvhIz1UAZ11TYNzSfidEOJGjTJREUSbSjcai2Ke82KXEz/H0vtToExLzk5M2B2g
Wn85cw75dveCXgFtENIR4EHLBJvR7BeqpjQ9Eu/S0Py/K5iLiWf5juGaUGstLF9b
QBE843drJRgBumCh96075nshEdAKsThLN23fKxokOkZ6XmDPEsnQ0DmeLH4818pf
/ysWAKH76swDjsyNNyNWUFwKupmfRbKb1xvjx/2rsnvBmJkC56WpLJq67DddSZQu
I1TjjS2HCslenrM3yaTaxhoa/ACfOlMh3ICpiTY+JbYj/arcmma0/PsnbXKNQbhf
ctVXRL1v/97G7I3DvDohq4rChd58KV8In8KHlZjGPTmAvgO84+KYW1oxXrBI6BGh
AQaW+SWX5lUF1hHXSesEigGXiW9uMMktO1yjr57+OQL6GBLvEf++AcCYMjzFIOMW
aV/ykoB/xUxA2Z9IgbVu6xmoQJQniZsTe7RLDXzYnZre58gvcSfLilll0R07zRGv
Oec4BgbBestURU65f1yABmLtl93VeoT+HwLB2OHR6boc/Cxc4T4iDbR3Sv9m0cV2
LGywSDEoDE9TSrvegvCBl1K0IFej9ou3uZGaRz9cCkYpOeI7GB6XcLLBHz5y3dGF
UcbtsOL1wOy+X5GFDkg7gE+IQXDpe3D4ggQ7O7PwoBhXmqBAexfTQXOdPMcHRtGb
OGBHeu6hpf0PmVYErQjUqpuzhIll+lK88WJQ0NHI9GyqhuWoDig6V3WEqNhzpfcE
wukO5b+tOKCNdsmwnHsTlrbDqrmfVpdxUzydokZpIIKH35UoF21RQBH0aJDu7dyC
RAYJLV/WuSvj69TnhjjiTRovmEdE5oxGZXbNdWZj/59HMzJTbi3FZ3WJhg03g2ls
kjxch43FUUZfH8lhmSQ5Y9tUIafPFKFOlhH+yPZe3Q+OmiXxNNqndTJ1jdSH3OLH
VwopX4OfWKgH3MHcSRrJT6Ufm6DEq8KsAjWNUvsMCWjkN2PE4yVqxq2bXhH98/WV
Bj/oIIaakDw/kBNEQ52AIfi8FffnHfjkIwDE2Bb9El35q8mMVIBprHXiVuVm4j3P
WNHQUmKf9oCJgL8GlbyP3EkqYXqQVyeA1rSAiwfJmIarWZVKOFJhtjjdENb4PyPy
6FCiu9qeyFHf4dlgAOWfzvuslG3reFf2EdTwtisgJAaUdgGGytvZukVzWVLxiPEq
DmGfloebLvJ4TF+QaIm6b5sESpH4NwlEhxDlaMyc4c7cXU7I5ZzdXhtUkesXi/sv
Tcgwg1jAYsNW3kSnkiRRaLT6krG08wll9/YVqNvtqGP/atGlEyyFHrYKUEqUuwpS
6c0O+5VjGcAy9P2nmG4fUY1wlXhBS27d0Ws+mrUHmpOd5U31x5XL0vCo1fYjesEW
9vpLyWjkpz5c1jbN8eHm50HEIyckC65HHwCbjf+H+X46l8hz6bNZwE6+9Lqs5+U2
2tglvoIpO/ZNHluhDBqnPYVpJsVXlGaRDfCGD76ubk7ugQDCKI7/TTVbtMBLcwd7
ykvgvaP7yZO1oL69v9j8AzLimLlLUQN2+t9xjit5byjR7ax+orqceggHD94/7k0w
xuOZzI3MiSLRspFOe3YZGp/VQ6Gn22rtkcXdnkA/hONUJHExWa2H8XejjDzokBzV
1CgLG6j7UnfnIofYVKuT7/bL7NCIU2s4CuRxXPxHykA+RZ+XaPyDezg88Wd0Wr0o
awfu+fXDJ7so9Kcn9oBAfjIQuCvmgCgLKrXK4HcDfkYsecwJc/xScnLQsCcjqrje
6+5N6oyrfZAx2nfUvL8Zf89Wn3nka3RwH668W4UY7JuwJSQChjrl461OwZ2qr+rX
zbD8d9hn3gVUcYCum+nilkJoBZxjXCMTRfwO+dHGzNcnpOFGeooXan5fOKMdZzn5
hJ6nsNUAB2gdZSJFHpvuFEZ4LM+yyaoMGNJWv4x+5c8b8/147hIkkvV3kXAeuTUd
y+AdcZGJ//XsFltNUttGgVU83DV09vrSkCgMM4Yg2KAMyuFp4WYxezh4GPAsf5B6
EzeJP2q0w/kUSQ5i3L/UQhWNEfWBi0wJVqrda2mC7m02r/iWpTwNzEHHA68cwe2E
M8GZMqBbNz1r5lx87JVbjk8VugsqJm3+fV9Y1OaxgJWy7l3WnpcSSWYqkmLsb9xz
244ohHlRCGEgeNTvtzE51WEgSgpIFuWFi4+veZ+bH5DpVZ2tlZFnGqRH9oVPDrw1
7FP/PpoW3wbEmsyU1POgy6W8KNtfLJANTNeRz1lFmZpth7xQPkOCPl11nE0pA1sG
g4Y1yS36rtuz23D91T7lZUJVq3S46KbWOlOC7dLZWK1PT++txxHxNnWtr+Kf7zSo
UHsSMMqwR0qYQKzQ9khs5h4ribIzkP/J0r/c2Y/IJ0io90wID2lb/E2eI+I9AFuM
I+gBOa0+ZOhWPz0O6KiJWS2JTJGLmNrx9GLYujXnhcsW6fnWgWaSzIbkb6rr146u
XIJd0q5wokX5kCGj74/ayQ6ZJVCeS/ahsz+Wd5zap4qBzar+ynK9M6fJDOifs92x
agH0w7duRuVFh57CF7ZkWs/7RjeW7no1QtpN1NYSx8HU6AKEEfNVLoRccQnPUm5u
ttF8l+biy/7DCPyeLeutXSAS9EjYY5spqKAkTyypWQLL/P5kgeb5c41QkkL9Zfar
jmoRI4bnkcGrDYBYLbINhqeUP7y6sAB2sXnU75VzjEbkg0kJPj3DuqjRovloLyUR
5jyv5KcWzYzUS6s5MYks0mLt7TIJDBX8FUy7dlbzimU73rA/e0WeVw3fa+2X0LBV
0Ww9S6a3tGoe4ubO0ag3rLmnOKxz6tXfbnOUcvptpFz4MpMQd54ZiBminRQp7VL1
2KsV2UdkXeRjfDMSRKppfSflqmZ6WTLuzFFfbU788XjKwLUmJyVIHjdwhvgPu6KK
GwsBp60EvAOihTagJKlZ3azJvqv8Je6GVM9rj8hTAETpG6DKe3Eo0v6GsFyuLwH3
/FpD99b/Y8U7Xrp/8RkuEdVbtOn3StSUqzmD9VsIwthyEWYyVXmM3iDXOtOC70Q+
w3M/+DuFkGKJnOiAMPvKZ12aMn/xoqlQH/0zBTIOd2NMTiu1Zzy1zzMV2ok1a4as
A5rOONZ7DfkktwvwM76HVP/I8x263taNFaxqgWepiEaf7ZkWekKXm7O3oh/VuiVq
lxElHvsTUlfwBbuznoWhucnrQYsMEZK1mC8vIBXTl5znV2Fg2n0vpI0nOeJBHHmk
Riyzfamido48C+iAA9JeSEswbAzgp+zmOMOzNHjp/suQOaJwlAem8Ui2gSTpj/Ry
nqNOURYr1kH7t4Gm3mkZFlsv3NsXAUIT3ej7DeMWA21CdwH1pUCsYjxBaMM15rYW
xKMJUpnL4hdaAfTnUluj8O4druUdiztyGRG1+R2Q8OqRizbueXxs+SjnrmAvgJma
Xlxp6Lc4s57aOtQi/3SWEOf/mqyCLtc58DMZMEPVophQFMTVRdVxUffpkMMJgs/R
huReBKOGh9VgGJWxj5K19sG3D58vkKR2UP5VD+efi7ITqWdQAubC2lSy9sPIJ7H6
N9pTnxDsYSNivPJQdpnQ+SljMQfeWR+NiUYJl+0t/+FkhcRacMHrxk3LsDAh9T4l
Bt8HtRae3ihgJjGcfJ0lm1qtNOqEPuUrY5wFBStACa3f4D2jWf3WrDttFU8LtVxV
TNWwDLr9W3jJofa6EX9wiC7MQNuMsJbSigPqXbH5Zoo0QqEcepljeO4BHY+uUPm9
gqV6YkOsDHRotXzOhDMeqFR9dhBpFtkDivmTnfoGfLLiy4wHLpnTS5fhdubh7xPC
uTJ2wPgOVlAp52q4Bt1fdHIVlc5r9WuQO+70PNx2KmpTbl1nBixVpq9ygtsrALcQ
+69pIOy1REpOGL7gntNS3XW8LUL0SvEA/q/6Pa4ggtnuHE0YDZNZpnqCODeP9YgX
3zKFzN6Y9a7MKb4Uv6hg31d3g3OazJWfvifKwHwH05WZrX12ohpl3hFZ+ZBwm/7N
eHiHrMyl/5OpkOFYcRWY/Pp9qzdkIzaaMk9J1+Udy2AoBivQs1Z8QYBTGIvmJ5Tu
OFIqPPlzL9SuSPJhqalaekNNGYaYQTsPGvSz3kYRcmJ4Ynz7n/8CQg3dNCmFZ9r7
Id8uocpCxFJU5YGJiNGfuPJ9GForwofSvNB0/b0cZEVCiwGId7ciJwomt278tdsC
cgmWshcpCVIgg939LJ/A/rtccde9LFkhm6LoXjIPqPdp6Nu5jbQzXwuD3Q65yjl3
IOIMbv8BUJPbxs9h3km/nnWyE3bGgF+cxA2WFC5v3ZROKmIx5i1+do3YOhVc4ciO
cFy5ndJgiycMC+ZM1DZm78j6tpoB0SWcxOg46XT8Wqlx5IYaYnDsqBt9RQzBA/4G
S4Wixnz4aFMEOg3KNrVUheTqzP/25RY6x4AS0VLfyeYoaZUsGNY5YiPlfqS9TjxA
v8sDN3gLjcdCZBjOcOUGuJl14p6FWvl9s6BqLn/O1FARE72zbijsGxmzesnSiYBK
Q7uSQEIcgT9YkA9u3Y556m2Jb73L0LN4R98VKAaQi5l06p9BfmJT5khWgu+S8mTo
abzodTJnen/nWipkAL5rM6xrYyS+/LAG5+58tqrxoZffu49U3POtcIKlC71PA+J8
2X5/geGGZfnicIzlOL0rD4v1841Q31Wlof3QW94FR2Ku0sH/eY2QUvLmDef54ex/
b2ZAsw8xZ0tXCKe51czci7dGKIzZGrA0i6/L5b7hyw/63PQgKDcf9wb3FVoJM6sW
VVZN3qmtdHLufRWIYakgxuRuapk4cGQ5b2hu9Yhmwk+v/SsAl8/x3cST+dxgxtme
Kxq7p+Al6tZ05LUAqRLrJ5Vuc12F0jPdsalOVpCAM41rqr523Uc16N0lwkJmh6Ao
U9PsVni7zfarnvkpv5M5Ggn6jts2dcGuRtCPDgrzK8gCyQgtlwMPcRjB6zn7aBvX
lpvzjHQS5RYQxhD6yQ19VfukungJe8X8BQWrA87o8FxiLSPREdddnCQxwiEISm0E
909oZbx3kwVsXAsEOGiZq3Q0gfkaNEW/zg69ItgK9DujNq3+fkxELTNANT4NibkZ
2qEJ6cbczPAFcIY+C40nixVC4sCpiaDfmWoCilfOI71saJzAgXOtlFEsLLs7xhh8
FC+kbkYugx62nhbA8+kAyeqJsOiZRmFYOHL8wT2vlLLJ6/uZHgfw/iRza4API9O9
A5SaToJE6R2hUPXHldK5muHq8LjTXhvnTulBHdfJ6pAuvYY63QBEhC6luVfJmXyC
aBcHryhDSu288fbFAqQBTZiH0+EybugvwIa0nh965hSn/FQ8VIj+aG0DPh0kTr72
qqAXn0+ZyncGZZAq0fepJPeZJKmfZM1nXf8pI+Zw+0iFdq2SuZXonMWPQK7o/Kma
7KEq2fokmYyRUiVa/StlLtEMtg61O55uR6e99FzeydHmkpSmYQ/eHseKRm3zprmW
y8YCHIQSnI2O/hVvEc6SQQdSaaUc/HhE5hh7SKbJjStrPKlOo9rT8xy4jb8AZM/i
VGf4rUKWG2mx/ssJZveI6XuHCdh9Pr/aMiA5YrS9PkFhLUxUHUUBo+Tj3VRRbK6u
2kTEdGNMQ6yLtjYJ3Cey6q4iIQ1IIWvzISNLut9CN+CMuk+W47iwWiWSHeMB+XoQ
Jfa0jwruaN7cemT+ZZosF3LwnKATB4aIbykuaoyDcAxeX1DWnp6olc4M7yRFRzPs
HeXSqL4wfMsEtwHFL1ZXqv7PwsWMyPTYJpCN8bHvlZ7wCN4+Ow39wyj63Cn50+yp
kutyq+1MqB+PYohKeyd6XLXJiWJCXSMKSucNsxjRWeIDaRAxWY8AmAmbKBkE3xp5
1AUUXz2mdGS9aIvHVTnmcHSFGK1F7BiZyw2MDjt/mHiqdFwzFJJdMFFEE020VgDr
30qNaSn6GRWqoK/4SBL+1qiqyYWq8TY/GCW2OIoyrCGa13B6g/fLRgKyghA+E3n4
N+aLn4VyM1WTV71uHupByWr2MLNjhodfVuC7kAKVMFCL61xvWWga8AjtCLOpZBbh
LJMbBe2uYjjLZ2oqlHBZ0Rs8dhx45ltA/dN9cM7KMFRgEMy2g/j362/xouDBZjtS
PZyFp3rC+q5TG2zxLqckokjeqyjKyBadSjoYffUfb2eWjsC1SG6neoyEw/zBs74R
YGHYCkX1VaB8rgYfWiYP3Jd9N0JKWdysBu/xVbdS+4Ds+gQsct7vQ/oDJYnp44Wf
Q/wOgacp4Ncy7zk7y5uQYctJ/4caAuXVRVT7K9g4DEP47OZVrOGhQUAIimzQ9fkT
fFxBe/BNOQ7FcZ3jT1IoBHprYVG5GkgTKs9sMiwm9B6LCvYzcCDJuLi1G5/hIHgn
1hToaXkYV0p+8xZlxeeL2oNKR4IgUdchXUhCk3JsJidlcPpeHo2f+XgPFpwlQgk7
iNJ4mnOrqPRxXrSjf99cjTFZ5IzqdF9prj5WeriUadmJfk1mp0+be5soaJBaICTE
7Me4bvuH5Rz8QhyiSJAaqRB2jviNdxX7YdonJ6QoePompBwm6Tj8ouExKLW5emnZ
NDLe6cLlwizBas0Aw9p+caD9Z1yJmfe7UlFPeo5pVOlJA1XmUZSi9eNQ21fo2jBA
Gpmj99bN+PiH5xkYUYF9zMzW15kPJIA3Tc/hM1H0qLZdejgkdXz5VA1LyK0iIwyR
2QDe+AETRMuA3NbJ0gcWJSCqaFIk+1UBvA7vKHS2YKyUdkZw5mJqqgx/EkMvH0VM
ouM+ajdDUYp9UquwDUxCu2qU+BJMp/Sq4nCjSXunIfFGGTpcxyt0z6ML0qOTJNa0
b4TPSaDALYqVXzLJHkBRY/BIGDpgrPF/LCjddLFOpe6Lxildm6pu3Z8+zs/j3izy
rSpseFqoa+FNf3++iHmzmwVfCw/q54pK0xPUM6WvIx5OJazEhAYNbZUfSHMq6B72
u5FRqKyyl3TwwOeq57NMMbmUSkRuv8s5dhFeXj5jQZV5pqsEMFeJh1pJlj8HQy/t
OALx2x0EF/XC7InuIEEkuXF51S8nrKlQLvo8aovYYLbYqhXEwwXdLNpqqEF8ouzf
nDC5hyTlHrbt/MXkepq4Gi2N3BtWNsRTTMgjjUqjFDJc55v/tZfsuukNe3BnrGpg
UA6PCLwK9hkkU3DV6JjJ8KPtyfLr8+FUsQ9bWYLnTd8zbtkMnkhB7+dWOBkI2X+a
lNWdXI1fVbu0Oa90DBZcggvGa7lEgpR84WgzFi4ain09uBYkoYWuWA+IGafzdGM/
03lAyqJSMMR06XI9OFVyo5wPGn0VSiHgJ2huOuzxvBlK/dnWrB6szEbthEZgsqaM
kk7WmhFa7ANZol4BRi4UlOeE6YOT+zV4eIzMcB9wW2OqprdwstKSful12qqv2M0n
yvvMXYmbx02moU1xWFnloYiRt8k2r6aYMVdcbYnJYXsGPJPl8w12C8k5bOHxlGtZ
0cLCaCjp0IcfGjc06X8SLVKH82tKwrs7xvfXgkIYMWDpUYsA4DbTRiupNklqPMiP
kdw7kxe8Ol2QGNfpYVnbS7CmNFrUlWtsjqjl39nFaX2aCs16ZYh5MhTvGuKr2Gcb
CSQzNU957Oqp2xWFQKpKqJNdYP3LaPW7RnSXTmNpGxy751gWh84NOoDnXNhxIfR4
m2uiT8V+sS777W+gimD3J5srrgN6WLJFkaaMqMZmJzov/lCc9nGqRv7n31lxLIwy
1WCWpIEM0RRokqudoNDOW10Ow2+PndIk/JUazc6dVBsY9OsLU6Jrj1YeIdJk61Gb
SqBJ28DT0M9uPx6U+OIxR8dNBmHNBfzv4xOASsfmXSWxDmO6SEMHXVicodfIaaP/
EVig39QG3q+keIIwHqscl15pBYO26DTGIYVJNMm9FULlMDL+kUKySosKwfP8j+vt
IbqkGxpceHTeBk5jDVLYX1yCjD/6A6goEcI5ZSmg36jr+BBYD5V+6SxyoW2N9Ogo
hKY+d7JDnmNtStcQH6zTmbN1v9tDP7Ai0C+Qy22KWxbD+gqBqNYd/stCYNTEHfPv
HWNXwthEY3GsQ/WGnDsQNEi+mZJKvPudpf6ZKCWlgh7io6bWInOVAdXXebi/sb9b
0MHE6xgZX5WGf1FvRE/JAQc/DNkUuPbDZ8+G/WyvOVsnnSO7EZFts0M2PIhyhl3K
SJZfYh/kvVPiBD4V77BSf4gsGvqN7rfRDJuuB3uXKBJzRsSvxshSVXjc3Gvk4B41
912JASq5KrGFPqQYfXKEJNbKc+Shzx0qh9gXFVrGZY/hMr7pUj98RTUIVTNArciz
0S7Yzz4kyblsinCy/AAkpFD+xtHkv91oxoECBnorrCqwx+4Cbv7ACvqgERx87OFe
5Z9G6tqVUs1ExPfbCPBhRsREZpcg89vbUsJSLhGzQyc9HJgO3z/Q4dRbe6v9sfyW
UsuwJ2jRxGZcV/HklT9icowzez46yqdiT9hky4SVILTfNLOlloJk90xhhzQzh1D+
kjzfhclOsxHYT2Wk8ps10lN1nEUmL+b/MFfGcDPANcPrfuEPB6Ua3ftrovYmEtIO
T/vvapdt9a+Ogxq/aDF6XHY9ZfmjnOW6nRtisO7ZB0c3iaj8kfXA95OksXFdyGTS
fAfsjVMfNs6FDqe5ZRhAhxIVjlnO0N2fI9WH2VC6yCHemnXcTAi/rTu1YPxShwoo
P5lke8P0sIH4z9octsk1cTMHdkl9c88UoUBz4s3bYiWzUfw4E/exn55BuBvi/jek
2/bMg2QQMBf21EJgnYYwjeMxINYQD0l4AaDr9gTkAc82Z5bAWMUSGFp6gr3wcBdO
V8cbu7AQ8uH8VQku0dxH2camA24aPKVtZWVRPmSneq0dZx2YtZTp3InsdgFiNgYf
0Ar710lfkjSkAhbLR6AAaWfjEpIoJeOEaoCevknNgP8=
`protect end_protected