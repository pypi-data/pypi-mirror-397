`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQDOviZGMOVRKHCOdT+eX3zppN9pA94qbd1FX1aLsDwW+
Mp/NmYaiIf6+Ew2YezR19GWRwvAZKQqzsArYk141bcvJMto3vYh9BKqHxPl3D8zL
DEDwjKHLlUtLrfAGczyItcJhRDDBZq6tQeKBCTyM/e/Ruomqzm51Gppwhbi3h28x
EiVeWJsOqbwuvsB/e6MdydqTq/7fv/EEhHy/K9mGDJFZfqnuIcvfNcELjd1cWfyD
M/skM3VXl6J5pOxo+95lDdPBWauYL/QsRK9jmVH+sbbhkDs71LuTXnKIv96zEXl6
FzA3hYbbX3uU8P3CYH0DoK1jUuiuZWjK1fRbxb3zHjUZlnByuGjbdkq+nUhQcUg3
jnfrTHHEOH1M5RbEySt/cBCShqxfV99FrfwHjy82yixhGNS6TJbeJbFybev40pj0
+mwHNHKTjzIa4+qFaq4GNF/99mxxioUN9DJ3sWHhBQamhby/E7H9Dz/9jjMklFOp
hJhZFalbqZQx3S+ozszmm+OhYayCgbSwwyw80rOmRF0Ljl1/zf4OlQgFZZmnTi5O
jnIbwkE+wPuyf1ZSNki2v47j8gfy/3KrIDTnqgYu8oK93TuNrwUMQYuxDwq3lMmS
pvOmwGUAPpPBrb5/WFcNPyDmieos4Gh3CKGj8nFKXyxV6w147a01umcu0FP3eLZR
Z5QAwZHB7G0eWjnH2UJCctN0keoaoOD1RiWEV+sVPgvrH7OabSkA0yBqcEQ9HG01
9VOYEk9P/K1SXLOV8dLfQXz0WCymA2IiCyhjpGbO7xQpRx8JxzNLDlmU6Q91VQ3c
r5ULy+xl01RTs7aiRhijw0CHH5+pKMEzPp5rM5ZXaDRJviK+pcuQLtGhPrikSo4N
8Oov6p5CsgS/nkSd9xZTboZi2R8oMynTwOwwJdrz3iYM5JNo/Eb+z+mdsd+zxEzp
8DCEJm3pRGYhIR7oA4lGhOr10iuYcG6Po8qWsJys32b9vkPwu7Ntkc7/1XYi2564
h4Fv4116dhhSSQNkQd9DaHV6C1edXTR70KmXMzCXQ5c9VAmpff1ELfqbw3b6XhOz
fJZXtp9ulJKwhrKi5ulp1G5C6D8Ufkoh+huhmnpgFtAXSNLO74Nb3xdYSg3AtAO1
bR7OLPyADX6YNyjZSXlaU1K49hIhN7Oq4BgHOg8OHm61CPdJ5+OlZfhCQL2fdx96
OL9SQHN2mprqOmLKSCxUCHVUgV8pTsGKd6cFnJtYA6L5oO3ZJ993FxrsEjolQdQw
S1UJvbSVWt2sj2meJaNf7VNzkxrYCSHrM0rhFTPKqcppd5x7RvA3B8P7SeBYPsFb
mwqOEqUr6BiYZyT8T+mxcEMmDRmPFuk9PVpIDxVG09Y4twwtD8m6sxxG+o7kQBqu
ajB367dpsjyx9Xz8fDgivG4OQsBkzO81uGzw/DbHCw/mg7l0UbDmehfLbPhpJJf+
zzVi1RVLly0OZegOg6DDHC7iXFNc/Pc5hu+nlfwe7MvOlDalPQp78wb52pHOQQD5
a1Px8/1sZF7aDixfd2x9toSVYl/Ml791cz7l5CSVSsOupIB+H87IBYrsQ2sJhClJ
ZI7STwXSvYhHS4QU0AK9NCQwkXhe26/MTYE0QL8Lg8QBT5FlAV+QVMueZ+sJmaR7
anw1DDpWaj1yhotZqZatIISxpKief55H9NDGkHT7jtJi9PfqEM5ESJwrJq/zYys0
CKx27r+dJJqauzCLSc58qDXPREIXeF0k1HgTBwnLoM6RCSdPO1PjfSwvfpyObmuL
AKXbPNoO+PWdfMYYobkGCsh9YVuocrUs3gp5O1KTosCiU8ixVXQriuvTwOfNBR2u
mI6SOeN7JH19EsTrp0+Sklb52Nx1hTkoWUb2fUCZaKW9KbJMHZeWD8YiL8FxcwQ4
dTGSJ4s2llQ59kdFh++pwIMXpfphZXA7RxLkyfP/BWpxAswHVYYtJJty4M/8lNiE
uxzUv68uMKd199yZZNnQpGknpdg5R+nea0OMcyE74dOSY1DEW96G6zD7UkNRFknT
fDVZpCwaAaOFG1X411ULFK34oHf/k/AB54T0qGp1QQ+RLOKh3hHmt9vm88znaa+u
k+4Id5kTFvBB4i4Cq68eAdhxeDcLd+SakWJoRZlDih8u3Sx2qdFk8D8DteSwjJjJ
sLJ1/tjge5fP7fVal1ys+W2oDtNMmlTSMzBY1a5OqsGx3n+Cp2W95d4YNNPdOKQJ
Hp2wuH5PpXxzCS/DjyrZOuZjW/bXunXoaCoB0JWy5Sb7aS39IMYtczV2a9+ekvhQ
dM9QgsjrB7in1yqp5t2pe0mWjAYe0Mg2u3cNE8jP+VaZvCj04jIs5lUYMwvmYSJE
J4WitDD1LD/QQpwEPnCYTkxsn4sajeeod19D3QqhNQuqtUj5QTjGJ3WCNjri4WLk
r2ieoL19M+cUEdO2xGq6709kdXY++qaiucrNQ8yB2TUmSQRVnXp7mme7Zp4fTjNU
qyVLEFXbpRP3Us4dkd8C8jTG8AVuEgO+fLS7F+urGc5PWunBOhQMrcZ5cBxDad7y
bZsjGO99iGOb57C6tFT115UD3OII65d6Agki38lZ44FjnviWalSToQLMYK6MSOQW
eBRUQKUUPsCdlYwm/CkNaxoS7P9y0s3+Tp88w6SU2LhL8IeMn3duUhNJNJaYRz4r
Q9A1Byne7ewJvipDK3IRT3J6iumEEtJMJLirTsN1qjhW+stwc9yoFRXPKwHXjq3D
MkLQEUBS3tPA0Odm28axcuhhxQUIOCFI3o6InIl/SDDSGmF8u6MOWbKv0uF4tSJr
J9+qdMLwyIjG9FQt8FI+WdfV6fGPvw2d5kHLcaW9rdS5eSP4PAwJoptUX8bFFEn6
ZEB5+fhbYGcP9+aKN+Tc1XWH5ZJ+Vm6gzIEgIHNBGg/bJo+APhv2/YG9xVDU/9U3
A0LoMz3fU1O6Uq5v4U3QrXil66kbQbFGJKxHLG6FTCeV+DfftLq/43517goYZmig
x8HlMQ4DHcdXIRN5dWlyei3OnhzK2LgZGMPZNAwPClfAo2xSyE/H9VCCcXvFM+BQ
1pojlGpMheVAp2INy6rjHVtYMWOSmqEHzahX42K2Td4UKnlS5nXSyHlrwZkSLe1o
y3KKYN6eF2f3LKK6zvNL52rQIPnnfy8X6LL8mw0ZOkVebnrmVFNY6YzZG4v725fp
GX14WX9tqmOjA+dmcovTcLgcvVIcNvT+XhchgWvKmYKIbNiy6VXrNXFwv44x1CaU
pUR1u4fEw7H2xNy3vGq8sG42s19LeLTT8LgnAbufvy8hOiGw7fvQ63LhfBdDKUlc
1fKP7toVGDfoNeSpXlQSuvuXwOlD0PlHduapfKIKGTXEIL9wopI0oU5SztEWHjnr
G2UcDr1Y2Za/LVzGffbDvIAq+IETyCyWD9O8OMj+6tZILieyOtcw5L0S/u1rC8Hj
oAP6xgNsIGCv/phSscAuK/zPRMU5hfUv8gghj1MBcGHSB3vgNFBenzFdyNx7LCRf
AqOBLhFo3W+muYOKoyn9ZAItLCwykGRDU2RE6U8cCTi0GMHFA61nbw4/FTaxjz5l
bCv4fx8g/7rJ48ejjrb1SmBZ6exdVhDEOrAkJBMFn/YFNRjH8o4v5ageFTVyt5FJ
aZGiC4wZbI9/Q2+cRshUii0sF8DLuK9k1WpKbYwDZveA4mBju+kzpx6JS8EvK7Dl
gPB74I/radt5klNgjLRtAbXbe7ubqc545epEK4KaR1AEZD070Ey9nAnv7ZHZd6+q
rBQdDyLm5aDj/tLMbOf61CGRxF4G1mzk179iaKEOT+RqEo4+0U5ur2T6BFwW1TqX
OFTmVjB2UfenXSUz3aEQmdZhuVEDlcjFJ6aFwL/Y4+zf9za8MaROKaVkvDEFVZNg
hu2KZIHSjrm8MSBzLhcJuTbj5oK6AO1rcvHl3CSWLk/Q3VO5vTDLxYgm0YyBuvyB
FWnnZRzEbBlSIdJ+P6hV3/ERedTo3d/d4qd3m/ssv3MEmRv7kBD/b7VfrH1jUfEL
y1T/7lodRbGhVCJh2EBiSdnZ1aqynW0tWlnjn2MumZdlW33aIgn/GQ7AxSl0LcoS
u1BCpZt1GmXqS8gAkVQAyjEplhTxEi68jziu1O0WaNyTk+g9WAFl9+I8ijUY2zyD
RPdUHp1+NaMYN9cW9Y4GqE0Lc2d8MCupyBlGuDDPEtmBgaaAKq15Lw6uHvpe180Y
+v5xZpROJvmazaplM0ntK5d1DGw8nydQGPhWvJiwmYq32vwKYekKrsQhiYdqQsKG
qobN4vpVYOSLlTXeK7sgH5p/u0NK43cHEgp9CX0EeaZt4AxgyZGTBbUhWkWEUfw4
5+SeRc6s/6Pl8nFAiIOMzUgBYz1ECrhZDJ7xVVihVWOZhrEelZHfWwIjndFvavEx
dpbsZlcMhMCEeMETIN3qrOpPh89aXtw40Qd8RgXazizDibd9/uV/liDV6QoEZJhz
9i+m+IrRzLhy4dN2tFH8QkA2OkJkkVMW9qTmmTo2CNXctrTD0T9zZDqYeRA3F+Zr
96wAgcrMKr4ZMxbVp+eIOt8gaPaZVXt/+XPgd1zZLryDKwA5ILag+aQZOvBPp7Uf
tQDkolJClpaozwhcoc/YX7sn8GueJr9g6b+CKDRBsrgQSV/y6SSYY5Tnj44BGefW
XsIrda1ISmwkNPcsKPHUHpvG9qc59tBBUGLer4GhMpP9oT1aMgdyzRC66v1s0q4j
rC5TKqj7ear4odmTTOdrrc9dmMWBocV+d6hOA1obgQFxt3aON9i4i9q3QjWVfp2K
jTN4UmDDZV3yuDHYqnv3I113Vcohmh9+CxIvGsliCw/ZjxFqAE0ZF5xe3KTlnmAV
+5cZMGkp3Wl83vqiECDBQwnI0YPDJe1GnrDoSM5jp7zA1aSCEBbgJzca9qFD0gvv
UDk6yV3C3iiQlDIuXVI0AahJwX/FLgsqyH7MzEWCOrHeAW3ybr+0DSxnrbXvFRl+
YVzL6zBE3DiOs1t13uhVN9kOcGaDsp3ed+qh44F32UJ7WlU4DnrSrBkQaJDL0hI0
/HVB/4C67A0OocBlusdqIIFjtiY+EFdosfN+1iRvWrgTFMerN3KvU8rkf/RWR1dc
M4ZcRbzJD4DHPuPyqhUnJg0aleVem1jkIK7H1hWB/mpqSt1k9yrj39qEWs0jtMMw
gi9gJWnHl4vzvfojWHOD0j7iysQwAPNJ9RgPd77/I6S0SNgTmOGcWpnqIsgAK3yA
RBswJPkk/LJm1PSoqchvzcZjDGHIvG9uvKG2mIHcvokdKn3A3d/g2RfVaXGAn8i8
g8f9WcGQTu6iOcUAc+RU6BNI/7ouEal753h9EkO+wcFSexy6Xuy0hwWXOMWxQQsE
f6oQdq/gq9QTySf8NNozjGNQ7sMduwBf9J/VCYDairSALbuZwa0hfH7MosA3I12V
nvbxJTIufVN5H83J1mH57ezWA4XqX/RWubE7ZEyLgwCx06zLLPY3ziqi2cyt5KkO
tTXYMBP/t02gr7bg3t6kIk9znITtn/fKAkLkpb84rKGoRmYIbginWePw5gRQ6Sj9
3ueyIyk2SearoC3L0RN9HUA7ICjgN1UFL5Td8/NmOAyJ1PXyUYqSvVUZrzC3SBIG
53PB8xfgZKwXNU/1FIq+SdcmzmcH/lxRFdjWPbM04GDWGBhMZYWb7U/ynV47UrUJ
PW1oRQcEqZtAEreSDOjKAbNcM2p/ExqfIsRHoxkyRnKrXVxMM2fYAARK/QlCZWTB
b5hN3yBlG8YZ5Ot7/9D7cwBjbtNcsZNn6PL6JEHwAjC9jGD8+iMOK9bZVNsfh+ux
vrEWXzQgegsgUFxl4ILjnN4Nl+ReNX5jVlkVRIbalvHpRbTKlXZvk2YxJv75a/tc
ccO8vNF8PfLDWQOzsQROApkHdXRJ2H4lQUJDZrskTetgpGputIA5cFMTC8A1V6K9
zUsIGFCyNbnXhI28L9ubOKT/t0Lzihd1+12L2QNNjHToGaQiTQ7DZi4B1WcU05Mj
VZ/kU7I16ooPyyO5X7HU5Et5+H8E77TlLB4P6VkpzLbheb644TdeKmKNSr8P/1BU
9RCCpoWEfdY6/e23ZNhzVQPmUppp/m2CDlWx97RRnV7eT6J8k1J/6f5JB+F+uI7U
ruc2k/R+k1NBVjAeA3EqgHjuPwS+WeesO9bQWyo3tcmAXLJMM5gq5N6THDvE5oRx
WwxTjP6yg3jQ8OAmXQlg6FQc/XMFMuiKhDt+b6y7QUaWw9aj6FfvI3UDvUbQjLk8
M/EikjTXrJSxzcoERrCTjK5oBTfwiL5A/7Bn9qltiPYWpN068cIolhSPscUV4iTD
Ew4skNHpe+voTipMeaze+ReXypqeyITeu9UrkohF9foVXCTpuOV5zknrZ9Vs/d1e
DhwPUZ3RccVQyq7hx5AXpwFDO8KC2/5wBTXn/V5143b63sGG30pujGQLFQipqtv+
J/WvQnUeEPsdlyQ2j3keSvFyLkG4Bk0M/Rx+l3+pCCM2bgMBnUY5C4r4u5WiR1NQ
xAcXU57ICo6ou34X73/kUCTvMyVJX2HK4MEdozevM2crK7jR2fUhea5R1Qd0YM8v
Wm+KnCDgI23N7KSBSJokEVQLjhhfThhfeFJUYsbVFWU5JYQ7QBh+Tn7/fx0afA0p
lrs3kpl2ma7EupF9mcA6AB2B2cuKP3fvx/GCRacv9hilITEG5nmu++3nNvZHpKvn
Sm/fq537MDnlLS3kKiEBdhOxvZu75NEam8CJqqUEr+muL4rTNuvU1h/5lWHjtAq5
lhAnnVcSXvqv0WJVpA0qaDlE3/Xnw59RXR6akUTW4jB5NJS1FrdQy8rFpARujmjE
4jbMUXCC82fUP1lg0Fx0mjQ26hE5JkFhmhTuuRauVYy4/Tj6MS5aLpycBCFZghEB
gzrSfQu7Q7DN+Ys37xrF/jLjs5NRlkLpj+p1ojACJBWSdUsRrtVtlvwp8UiSdPG4
Uo78+aB6AVuU35d68eXSjTtlG6WGz2siOmqDR6/EdsTu4+nf4h1ib2ymLu1Mt3Hk
P6+mLJEvWcjqCJ/FWYTqUSAgFcJT1Yu4Ag9ry127TQHAeMzkhiC60Vsh8wYvF5bt
dLTI76SCTpTUHqF0pZU8P5qoii//bfAy5zRkGHZogycg9wfO91oOCTltnycqhEqR
T2JLR7y5gn48PFoQrAsiMotcwtnAmHhAlzPIB+vcf7iATklUyn2/Zq0Up2uNVaKP
S774eI3Y5ov3WIaMfAp+3mxzEAYydBeAdaB71wb+WVlG2v4uzjiwMXgLfBQK8qsU
AbumcCz+f/NrLOVwnxF1IiPPUoaqQ+XyumEJXRRjnwA7uu3hIDiHiRNBhfgys4Yi
VwK5rybj1ZMMa2UBMMU589Ae3fAL74Q7wK9rB/MATbSCd1qd3hT7v782N/6SypZO
ASd4M77Citzi0s3UKfCobSNH6dTAmOjckqdShKUGZ0tPZl5vF/Ar82cJNZE5xF1W
LoSOWd6S72v5gLmNi6JplhWvBWhUdwph9qzBxg4/gvzS64SJn4CRM2u+wxlHnsCF
+vraqFYj3/EXEty6pCEc9zg4PWC57b7nK7LZoe9eAUoQlRQS7ULJ5NUrixvZ7EgS
xggVdPlzVe+AhXjxn5x6WA0KK04GLLb1AVWup7Yn9RXRMQWNAgcOiolFOgCIOtQh
L6EpcSUCqfFQ1Mnd4wNXcf20EIvJTQZY25MGnti26gQiOskWe8A1pLvoOGUhzF64
5CQA6FiU6rHzsIKi4L6VlUktLiSDcuzo6o0oZD/Fo84E4awAtuOLyW85cX3/N5OQ
TpcHUV/LgY7ywEzQDp6HORnagrr2U4erHpEr6Okj1fd7eAFwW7zP1l836YT151bs
qfkVLeSew7adxwu9+UqxFErYu5WHHqyNb4c8fXEwIL/osSWvGgnJIv5QFIc78Jd/
dBfxLEAej2/XhpRa9pc0bYZVSpZeShxqLE+L0BZXqK59nFEK+86wh7HDsQka4puh
M+yNMlfWfD1GfZ6MrY/dQxO6JfAcGiml7DwYDVIH/90heLIxiZBnUl4ceJA9ByMb
t4+yypZFZmQSZSojHL43iRkRa6V5sN/DzzG82iDxQ58HmYGtmlyJ4JA67KaZ7ipM
eAqHYw+balAm5h751wItlBbCMEMjWrXiqhA6AgOLxV+WVAcLDeF3H9DDJ7ATrdci
7Szbp/1R70IgNOa3gC+FkvVtwS1CrvoYHUwIzjdwnH/v9792bA8sA5wMi9YclZ6h
0EhA81H65KPt+7Ai3/kzfAveB7jLtvCdrLB6pbhVJDJY0gTasqWKOY/sAoTGfIEI
3ZKdj0KblxF2sHKzYWgugYd5hPMRAmzfbZLsBbtN/3Lt1P2EeInjMFYOu6mzQgZz
eqaku8yFlQKYIfJD4020OCFAAP9yr2wdkhIWIFi08fWVH6SYExwYtw6LgnDtWVCL
lShBIFxe9KwAQgYiYUb6NlXd4FkB6ARL5R7TwNBeJPg5GPvldNFLT8f5Ml80CwyT
7xnig8JkjU/DycTM5fQz6nwJ6puXK3d5eKm3KzBtH4cS27qVbp+wSkWibIM6GdZ1
9QD95caeO2/D6wt/sa+lisUy9PwoGZyPJ4Xdv7WRsbM0JCMv+f4HbwKTu8tXWxlL
2mUqN1f85anwLlB1bIwXCWV3+GXNuX0uZxPTL5h+djE1Y72RhRU0p4+ISTSfuami
pYOsLKEcOhr1t//EK/PiDnnyBjJCc/DeMgszD+SxR9G3OBME0gh8zAc7sL1VVzq8
kd/KufW4oZ5KKFBbl8QZ3rKvcdBs4mDdCk/elzMi9faTnOfy830OliLTMWLA3414
vMcscaBh1xmEX6OJkgetx2+/OmVotwCXC/p6WpiLGhZrkr7VFH9SaB4GMEEpVxZv
FFUi/49IiRvz4r4iJRmQTpXNJb8i2CoyoZBbRKHVWvLFw6p+akux/ASNAPwghG4n
qv0mJD3hsUhPKaS1DWw4zNXFUiRCSkQa9Glzzlu7jDKoKgjrT5CztXzQ8kM+7P/9
p18Z+50LV6gSS52WEKxhXSz8NQDTGcgMJ+mFcaZOAePFn2Xlc5hiKXRQaJYFm3kA
oI/1x4rZuLrUYwc2CtnZH3u9D04tE/32U/6YVKPBFBF6qvM+EUd6dQWroSajBsik
tBOa7C5E960KCSLFl3YHgENKBlWcKLN/NiCbaR+7WHRtYYMD0cqbIxf/G0lYkpK+
8/OlsZSHHRVaUB7RfBGnDemMjwKSVqIpvuAasxETe+T23uzt9SF2ijn9hhbqE7r3
slFWhvlO6DPrJT3w1NbCTsAFnO95yzRU0cVgsMkcNIfF0DxYrl37DuEpY81qMQcy
a5rJyyvYCVgVWldioZ7hhAX/KpCzmDdpYj1fJGZkeHro6qdrxt+4bv8Oy20qvHUT
bPOq+s9l/zYJ+aeq75IQmSHTqnXcGkNfrYNHpq0gFQkyuP+gDVxdF+6h5PHFGSrw
TizLwwBE37HvGtYlGm5T+geReyLCerjVbs4xxLF2sKTXBxpMs2KrTnCe+b4vls8G
HJgIxNhLgDPewICmZPpqt/k7NoWdfMqKpgPu8ZkkV7bjJjFdV8kLQW3/Cj9JJCXK
LHFt2lParJ1j1Qcd6p9joJxD09QiqgaQYRAymMVH73MXdFw7Yvftg4zlt15D4yPi
6hlBIRGOCt5xSYUYI2OhoaU9ngkVcH44lB+OfvP08Gkp/Sn3eq1KJufXF6kLh+KR
lKOYHMzXLFWN8ZvQXZ371mLFHGLnKSZGjaviJAI03IpniLCE8BUK7QmjHKCNZ4zG
dujzElyJqTU/Y3JCWKRWyl71CkI4QGhlAq0rZBzUYZzPV7AfD3XdkpYxEisJyIPZ
fKBlQKP2TxN3ev5vClm71CHAGzhsB0dEX6QKyZ4sma79MzAGejFQz6nxpOj88ilg
kKKM0nkrk0rlnPHhVukAHod0c1cewVb4VnZ+TZIOM4NUMpRxQbqsL8WPlXN5lvk4
hx8ND12tywx/0o/pLk4wnGFQRnjBilhb0JQKrzTUguaLgcibcVd2MmFeyN/jGnCq
gBXSi4XtFMftkSWC1H+V5ha3p+aRDBROEtpOn69+xXAPPpJelkyrqVLOXzw29JnW
bEiqpNZbUpJMDAwUh928svDcPGCBh2S+tGqf4c1Uv54oMhsXKnsnhglcuD5rE/iE
Ijx2Ff9b6xk/wV7Tto5fxAtqIKwyaNO7nlSIl0fJKyYqmmj+dOfeINbhiF5+YXvL
+AF88WxTTjRKIOSgfGuqdnrHudMkyVICbCHEaYGPvWIxbQCf2UkD7RMqQraNm8ru
`protect end_protected