`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH0obzhlsarOKkTfjzL+TLLh968MUQfK0sn+CeaTcBgHx
yLzwuSxGdR0b28U38+CxOlybKvaCfYjetTTJIeh7GwTmZZ0nJjzcAx5nNeY5zkVA
psumB1mAQcKxDkEYw7t6ATziePgSAipMOxMTl5daOPcSLC5/M95HBEp30oO+R31H
/WJcT9EUWzxgBrqrIeJReyYxNaZ7AXvqKuSgzPf9+kd+uclGvyk3uKRsq84Ts7P5
AOUjwguKK3gmtqlKqtdsMepu24GzpiQR+IQvOURLONDr6VlXnev0gJLh1+SZVK4O
WH+2gQgUAZOCkMzN4ZISS/SxNjfk3+abziPJthwZ+/XPGwJjB5BF9NY5S4mKiFM5
GoqGSgMplfWmBWlO9FNfl8d05NXia3wWAv2dD6Nbw97irIxJFarFx44X5pt0kfD4
vS8XYi29DZdRr6oqwakB5vyyakLF4Ul2aeGpULihS5pcfrn7qxJNIOPNwSJjeEw9
1+wDvOqVgLK+ZcPVuf8Eq1gGkesxD+1k/3Fvy3sKws22VeyFqvH/LYxdLUn5pCk5
1HXEO4ySPwKyLsDvgF2WAba0aIU73ZpO9OneB/ZmWYVmb+j3gDf02b2O2cuxH8sS
Tp/5JBkmJrEVMAx/5hnJOax5gvocgTOXRh/fpX8CoOH+RrvoCwAjqdnbFoMsIVXi
f4gVTOEFdVuvrArgA+WODL91PVRAIh1mkBOhDSnpgFvGWhLuDLsozowki3eYtdWA
wJ66yz/w34RUag5p5dmAyr7u1Fldwo2pz8+fURQ742npTESGf+ZNypvt1uCUrzvD
0FobY5VMpoeWUUqow5cZiwVkgImlbB79PDlznBDgBBSfOBTW7/+u/use9iZ1PTkg
00v0PKIvK69Zp6/0ZdzMX7+uGUtQxXq4Eg4CuvHUHadLSJGKPMfGrGKt+BzPYhdS
4N+LEamtF6N0yJ99JGOg24JscOS+qvF/DWedCGtAAbKI0cEEyoFUUjz/96q7i95e
vjIR56/ssxhHB8/XPb3hSsjIW8hhYAYU0SqlW1GUfBUWR+EbLFBscRqgp2QWHLxa
P4WORgkWmgBPXoJ6SZUozvZp92MpDyTx+I9+VMtfZrrIV+GjrafHQFEUfkCeM4SF
VZWu1hGxVGXSR4bjB/f2+odG9fxwVGAb+geV2oL/XRmMouNlgxR+Wztk5Au1DIfR
0ju9z11LKzN4Y6jRqqI1FhaoaDPWFEFli0TJbMIB2A9bJDxmxm9JmrJK+jMqvaxe
2bVHXE2y7jz6FTR4MRwrlPNK4UtZ8d6tSXeR2u8wDKO40slFltGQXRJDXaWt0/24
YB8p+oICl+cnKMzBM8ZxOcUM0mNpJqiiVIE37atm5dJjMXyQMJe95iaU8xPwhyfr
RwequeOVctL52s5ut2e9o4HzdxVWJnrWPtFjcfsj9PrdTfgRxKseDhgYWzIm7s5a
ow84qozIufRduszrgRTCXTyt1MKi3sPmQpL3cgGWN6UnB+V62TO5fztrJohM229C
fcWGxvhSlrFg5xLjJ5Iq/fqWYrD9mcjD3Qdvk0jzzmmTjc0BsJadCPEYwS2iIKVN
eGK0c9R2jBwoq6ex8dJt14+69/XoTs69znTyoOMnTAI266EFwFD9Iwa30ahnS88p
6yh7kfTeemImj5PspOYaTTqEg8LXmOF/R3S60tC0TmB+IGuejjhKePAj9fcey3Dv
PuItDQ9VoglVHkk3pVU/NY4nX9D0enrwYGNUezyxdbLA/GLNDNJcD7XpOlFPo1Fa
UZona+3Q6aGUOg1sYv8hwGDM8QjwnpGGpwUOpR3ppuZo6eGI9BIr1ohJ3M9+I9We
RNtjR36ArP0tY7JqBWfoy5Cbg3wK6NZKG6hIEpTiaQFNivCd34yizBlzpEoYcghM
DgV4R795LFH0jJhB0tX0sTFt9IG8jpTxiJ4LycnXfvzIpCcV7l3Wn6J2SkFClnt0
swq8mowquPzMy7M0DlNXUrnLqXHkNKqf4m8DNQewRkStrrfIF1DaC/DnssTOlF/K
qjg4VduPuQ9HzAiDjCWOoY5xCPkvIuRo2EZHSCeyUJQM4N+n3C7sUtnUnRVycuDP
q+Pe5Qbui0zfnSWn+Cg4EZyeRxuYKgCvGbio4eaolRWojzmMqSuu8khrcomV2KlA
0qmG0YXdGSX2pQs17Ef0Z+34EzWVzAVYSuFFRdab8908Z8nc0hAMRPS3mkLZxsXi
Kgq5hU37o4ScKVwDyCe/rtEBD/XPnoylQNHf5xTx8HNG5/GL4790Sh5Armo9lyPm
qkBuEndw4Xt/Dt7YjciHdXCqwxoPoLT/J7fSSyIksvFYJ0YIkBt3B48Qj9X1eod1
/6d4R+tyzDZemoS1uVa1WjCaz/Q4tICQfWliWrm0HoBp8LQvfFI2z+es9j86w8lE
EEt6IM+YxQdimRpZ0cTPbgCuprcARGsg0/XfX506BbIIpBJkvDZYsEXuCb72fP2Y
BHD4e+f3SlCt/Xb1TuhkxhB8JWyNriqN94BJ4BL0erwCGqUifWxXGYxYV02VBL9L
y2vpNYU+sW884a3REIUtHRcisxMI6nHn8vC2KonaAfBky4Nta1lHkjcLkI7Y+mEF
FMDL1sYVyv3nBZBULw3RRpwEMNnTbJGWhC9OICANToXiNBgJuWt8FFmb8bLBbR0l
5jPkuoU89w4EWHTiOuFPSiqZe4YjiBS7i61QMb6tOIEID118UncfDuwcLAG7rgaP
VNGJsAAx8m4jiiOe1djOknQy3RfZlsJn9H3p3jsPFXwEURpFQCuWnvocwdJPPwDV
dE0aSHmPrYfPoL9KbMK15z3hATPJMF26hqRcMaFpgh4FaY/MWXwTE86RwQa4ompR
H+F+j3TFYGNjXyo0qlXArgKb9cWeokZld8ddBqFoLlcd/g0aQL5Y9Kj+nnbk19AY
YBHQp6pelKqLE+pSlg4CbwLpz2+5E7AZUb7vlyAlxWGDgPitN7O7HHM4TCASnlOf
P7S1NLq5Z8PgVrAy1JUIKYgpb9ix3U6AdWupi4DM0DGDZ/M8AkfGbVKh26NXdhHA
1wtT0eQwR1ZQm0uyS4luh9pJQNQ6Ps3eBZZehfxst8m9oHozlrH6SFZdiibz4dQS
M2kfR+r7nsUI5U/Ka3S/JKwYkfDwEs2uj+herMeYD6QBHDdzUMk69wRl7jsFh92/
BoNskfzfOI8fJe0zwFpBcvU4eNpTZXxg4yZJvvagaDS7wGYpK3S7QNKn603kKVdH
RMc0BsU3xSvkEjbkBI4i9/m+7wLOVnzi2uYOhAvIh0sAgqiyeWPcp6Omqef4h4Py
zF9o9hNjh7MsVhqvrGjoC3KXXPHICqn746M2hDVtPOG0uHpno4Bv9neeo9FwpjW1
AJdO0VTvVG/7bF93a/94dq++iNBSZU9UopvdXz5q6aHC1YnmAdL43mikRHQ25sPa
lET7KdUoykYjuqN9xyrqXoktU9LrcyoTT2ZCOOjYQqCkMVonZAN5evRBQMPHlpEB
8q5O31LpbIwh3UBYmInzO+0ZMg59OI3cwQFjpy6yS3Hdo2X4jAjGlc0u05p+m0Jd
aJMSKnZVi/8VIUFyks2prNT692FPvuzWUR7gma78rM3CkCMPQamm+IYAEaOniqyX
yMew7ZFvZIxPhsNJxdwOK61NfRz8xUqR65pdc67ycl0i3iLFvNo/dO13TV2Jw2U1
YDDhEjgABKG5fsh8Wtbh0YslFWOp/66WvKTh0JBQIJyPS9GnQLjcj9ufdC4rJV9+
dr2nXNkXA5r0aV250EwgGHIUReOhw87zT9G8JeyW4IL3yVJcpVvQYwa3Ab26sXGG
4gAdyG0czhDgTRWvGmH6thJFqjMy4wKBCxQHDc8pxlotVY+MObBrDaI7WnHvbqFS
FF70easBrEl7BzBYyMmV2b7IQVSmXhYLB5cUIDFRX0fOeGHgobvdvpLgftSb41ch
7zUW7JbxCxXxwvErjjMgPtY24UkZmZWdIYAzOhKedUHOl6dL6F7/qWa9MrK/Lg82
RsndMQtvN52VrVxXvnQnOA094q5YIPtBuFTeNAaG759DOUBT9uHCLD2W8T9g7gYH
ObwkemO7XwvZzC8IwgcsScTLKNtxZZOHs138obHPK7RvlK0ETtaPUe7cuIgGaS0N
jOsk1NPu0qnhpwVB4Y0E3p0dJjlaOO/L0iyCWoIql3lJxM06Pxq5XPYGxrgMZYxh
yF+ENfN4GI10Ri48QlzNtJLNf+LHLhl+FYYvOpMtbo83Yn3xDEZ2MoruYm4E0GeT
HvsjXiJoudmfwPkGyV15qKXvCWYO2I5eOhp3DPW+2P+jwi2ND7n8GIrNyH6pjLo+
QgpuGBeYdiwIacAdlAONTg7xDY9N1pjId/N1tu8RbVUA/1U71+EUcfNt0i0+bRZ3
D4gNlvqiJVAgDnrCJe2/MkLB0Iu4f0OEIElPg0/pHjPjDwFsc+pxoyKO+V4fbUgc
c/5fVjEGI5C9bN0Lg0kMcuvKTkOjFt9ZM2LG6YG211k/rmSXhKwa9H9ZpDhFvveI
hN4ScXM4JtnBpwliQMX3nuRnkXD8pyw8eytjkvwjshaH4ryrVu1Pk/Vb/Uqt9HBR
MhopbnArtCnkG7JY75Q0uoFnzNMJBSTmi2fsNkPiOjopIKArr46/1nCztjtRjDZU
SU8JrA42PX66FCsAEBsf5Ft/4L5ifXmya0VduXB+0jyfmbkJaso9KzhvoGrJfQsQ
x0cpfBGSNvunYMiXRXxAn0+OmdccG72nA82F9cZ53Hp30KIf7MSx7BY4uXXeMTQS
1St1sB5eWm7kxYCQqGm20RbyqXiHZiU2x8YVkFfjlN6enjfUMzryIQVlwU+duDKI
J5yZdJwF3iWgtsg9uuLgech/aD5tRJwQ7yt0AFUD+ymb8gjl0Q8HrrLJ8TBxkpZO
DB9yjkIB8EvLN/sYsWJ0wegJwp83j5EKLNctn2Fe7TrvyH0OuW4CVlxBKB6BkLR1
Xd41NheFP4lO6DO/8pI72OWVe6d9RPxSM5YIRmFvXtnW/UMTzj72cMFkds6ANqOr
Rcraqpa4Rmr3ihDU/+vi2pGFA8vsVc5exu86F8oTKtkepjbUt3VddiVLWlvtS68U
Brp/rddl7VB+yJ8VaSfcObNftgQ0Pr0JABNcmLxTkZPKcNDveJcH2Of9ZSQjP3ah
4ZkrvJpgvtA5jYT7xiI83j2xWFy4EnS3vMmyzSL7BepBzlmZBJUI0G1IQKH3MF1i
V7aMFU9hKy+Ob2HtOwwk3dThL+1eerMjbcKqOAnKpX0oCWvIX/j+B4FuiUUVjxF8
RJ53bL3nG9YGnE8iMXHK2iVKjCM5iiZReKsK+5ZXPdehQ8Xe/k/MtXLxEz207WPC
rxUZva/5cjkrGsOh5Ju4SZ9epuoXGdJJKyUhakPBPuSK4mEMI6BkXsBnB6Db9U/d
2NYY1PLOASGuuAJ/Rbk9kBNdA9qwjsNcozjaBHpILKNRLjR4PaEMmftLfYWMYhNZ
mR8s4MnGdk7dlY5LqLMJZhYtUt3D7ix1AEVjslmiSRjfl2Y7H26u6bzOfU0lHeZP
1wUU22VNsO6Q/PrmRIklcdkltk/TQ3KlU/lcjI4Du1lP2LjAwmdM45xq5WY/4cZr
DUAYIPPHTOtUV4zTG6Z2OrpOu9xTjAJ9dwS5A8di3F/QVubpoaGPngV72BUGEyTj
f/CHnQX/a0eECjtAIrQSPdo0CUqEywnOkbpraKnZDINh8LEmfqsuUGhKNRIAxqlj
XCd9RhJHeHGftNwvzrH9QemQuMx+Ujlti0LI4DXjcv3s3yS8+gC0r/EVmiiEKvZF
cuzWZAn38AUkrcYi2Qhzav0Si/7+5U1Un0ZjVTqLxV6n+WcUP8DFlMulnjHRz8Ys
2PmPfysXN9s6ofmCxFfbYfCiTWNBSLivX0mhjTAnMkEQOcN1/w8A2uGvOB99OX/d
3R2Wg9pMT4IHRsiAXKRkeFX8ihhRg4OgB1CXDENjOhNUvlFcWWrAU13CWPtLczka
Q1iPQgSUEDX1Do8ZV3+6lVl6zbTG9YJrzbrNPSHP9Qd16MjqBdBTHOgqyXm/blX2
nDOMmN8y5C/A78kVzagq+X6D4j1jSpcZ3ay4pKW/So8XMCJfSgW5WLu67yV38tm8
g9Zj6jYNtgZzXDmVO0v+k1MZh54womnOLdqm7qMknVYod0W33s6RVROeG5hgWHWq
rOB5lc/u1IZc1v33rFob/nYgdVeRI1T0BCSGKayHFV4e5MgHvNTGFiRvXT22QXzF
KJO2HG/fXbqRjV1SNmJSOiyd71HLGWz6dpZwrFWPH4qOYcbaWiHfgKPQ1pDgIQ01
0pFG6MhvRbTIlACw1YZqeopYvVLpm+RPEFcYnsbii/+AO5qsl64YJ2lugtEysxTO
EexWuPpx0qYoeA/lEQlTAr3WG8fqUJCBdk26wSAMEH9A8zdDSje80rY672pZx2lk
ANtMhke8zZVOdPseGMOZWxdVA64Yz0t7vpMDnes9C7w5VgX+qGc2P162sfV1D7Lw
4kLEAgwQXPIoMFnLia6OJaDXDkpgHF3lUPODlemRO32/XDV8p9UTg4BIYfRdzhLe
tScz9PZo6719oAzBoWO+7xNrJr4wcJMzc3NVSVoVHEJJ4rBsZI++6Ct59LP/EXuH
q2iI3/9m3rQDxf9eKgpsgGB5opuFdoEVsR0buwOGuZvnqqDEud0gmE5qo/zk37L9
5Jwcnr8UmLXSFlt+xjxFTkmk1EE6F3M643We4GZ2p1gFmILPoefCuXUmmLpQJOwE
62f7E7VLYKBixU/NDiQyA4TPkctdYLR2I0sdjzIqt9fe8RF/A8nqyP17hfPBnHfs
pGD95Ajjsze4pHeAKFysMF9Gwykm/mRYUiCoNFCsoPAcshvbzlTAojmg3f87SK9p
3NOc6ovk35SVJ6oc/xdeEYL54BGYovMpTcFvfbtKKwXVNnfYWAoGyXO4ICr9Mx/m
//sDTuWsD5YlNM5XIDo8yvh6NPdTmVq+OJ3cHjPSNvVP65SHBMh5WbztlbNnmIXM
LuaSEB2EDC46lAn4v1lgUNQjVduqE5Vu2dW7K+6O6LM1jtRpIUcqfbyXNufkBMiN
HmqepzRBcv2WdfYXQPxzotcmz5M8G4Cv3+FQ3e7fYHlaeQD9Qu/QW0ar82ZDZF0Y
ylDwwUEi/SDFyOp7IQICJ3wGIiqVMhlISeIJDaec79Yo3Evn/asZNyo1XzMeOT+4
bpnfToi5hrQwnIW9cGi2KqfoBUY99rHnSHOP2xDiw8z/urZTL9wc6wWvXzU4Mr7S
Z3ZMTefjieDoxtPp0WeX9mIQQP2omiZVCvqHPhZ+fu/5oq2p65ZlchaKdTDSXbN3
Cy9OXxqBXS91c1+LFq+VvP3xkvagIBLgKAz0JhZDmefsxeMww4DYcSC0PAydQjFv
pSwh90+LBu5g0cGJ3XA0SLkmfMO98mCqHzB+SQj5u72l43u8IBpopKUOw+jcE9OS
yv3RPBEPQA5VR4EiSDz1ta0K4H/TpeAnMKMP/r/pJh0V7m0r8ikSyM1r8Q+ovmLp
PJizU0Mzsh6MHUIuZmL3JDIChQHQ+JYQrOGTcI89367agvnW2N4wbXtT8D7ZDd4D
tG51YTDkvzYi8M4JGwTfifsI9nYM7SHlULu9jyFGtalADF7930b3DuJw7FCicC+S
ZAc9nrcYBwH3MRJQVAEo7JlaM8IlEWSnQGannJXSaaga0g7rZLfch+R/S7gfIrKd
PgbMMmj7+9PvEMjvFEtg4VPIBd5gof08sVftpkwrcnDjuqbmS7QxPv7Wgn+GJzCe
frPH801kios3q7C5H6JnaDijjQg9Pt1eG249kJ9F+k/lFRkZH/GIoq2LsOQfUE3Q
yLSzp/gDMj2rugFJRZfSJuzGhI1EtiLhGQmr0OkQZ16YjDvgibdePMebd7Ig61+f
g2IDlrO7YZS+a/nUojMKVv6Qw3R86uYZ2vDF2E/rfAhYAktWR8fAc/1KweUtuY0u
i1bXKMuNZwH01DhWcFylFBtDay6St6uBQnBSExS+lMapY/IlDhvPcc4i+FXXDw7z
2Yi7GLJcdVgym+YL1hY/FQNKjHbFVqLKFI8rJYEtYTCqQopz+7NVWEc21GwgK47t
EP+scHwKoi+9Xig3Im8lGdytaeq8JFhiSWvkepwhnJXXaI5eSYxdN0NXiRFoLCoa
ZWnJLAe2nLwy6YPN+EVflg38jxVGRDR/p8VSfax37TE4I+NOhO1K8AP2T49xOR+Y
Vw/w9gO9VElKRGdzwC1taDYEOUnHIT8nXrEd70KfhNPz8Lwz8nrVCS7QSygT3aQg
oSW/UnToZpC5/qeDZ3zXxbiqCmnTv2746guq2nSitoYNVE7ZbHuuqFV02U62p/gm
tkIiQxHRZxuA8POtVaoMugDE3GdsajgkEzSzsSNJjd4sitxx+MLWjrCzkZpeKpiU
tlL6bzqXHl9m4lrVgEoZO6BjKT+e7nxBohHPw98v8MC0GVRKqUlEKITKTzq3mu5A
MdH+kndh5cTPIRbhS2ffL/JoCZuDgfmMuufjxoEhwifP01nkh2xCKVXMST4vwq+w
rSe9UC0hdgGu0iHDS/5ydQZBQJz/cAE0084zHJaEVrMOf6dtGFq4F/VszeMkcxLO
Q9VFF3nxwDxtdBEoCYWt3RU8JCRMcfKfNj9zmuxyiUFi3RV8LzHXFPYI0th6tw1h
YfdMVpsqOyWaixUeOJxVtlhefugB1kqbQ7xsFPnbT2e/X5WfK6TmWuUlteN4EFy2
3/MleHKZGyY9iF59lq7ef6PiH7K4AUMKj7oZ9OlEOUtuoEjY2A6rA3j7biqfnEeD
OWJKIVBETaNLQI9rgzIztDY05ojPLyQ7jPKYh6ywaznu/iXF0Wu8KmlXHYKjN8+a
U+UaO0nwA+KT+ZhXh11Lnl/G9gj54Cy++3atkbz/ouAdsDkxevtVZlE+r5ktuHkz
OVmz1qTQRJXBr3ftUtRxrer8K8AAexcV4booWIlIy2ZGCdlVAbNwM2VaYUIppUGv
0uaSQi2PFlZe7twDKHNDRjaISgaxu11sxc6DQuYbCcPEYIW67vL7PnRKThs8tgPf
MOXcWk90PukAsyz+lZlEVOXMZTFBly5jIeU/fnorrx0H1a/zBye289jdsoPT1iP/
PH6t9Waf/xhcvf/EZqwrcSSovHSj4qJChAHQ3NTEAg5MOE0uOCZNlUOOAB5r0UQk
y8kVvsot45zSMDoHqvmtf7IYZU6CNCohpSuX1OnGyzVQxT5SVayGT5GStGqV+6N5
2L3NtE9vx7I0+oEFZ4P1rIMJrA2yhYm6C/hnL+wo2SVXdWaLYEj9EVrdsuU8GGSZ
wIuwzuGakM0N2AxEwU3cl2xvoHO0O49RYHi/21hpG6vN2fjBLfFZzvZFm7jkTxZu
vlRLFetz8qmUYnxn+lGyYGh7qg7FtEqlxrrePNHftBfuF/okfDtQrb1yVJ3yj6HP
8R4WbR8NRzIWR6V3zRBrOWwwS2dkY7fp+d1K2EAt3ULoRKH9ZQyYdk83+xVtw9lG
q4UYIdHpsmiw8DAGRSN6m1NXWpC87iwVC0N8E48I1a5UEZqPmAuL+3Kuk5Z3vzAI
uBCioR8mgE/gHH0KfaaoJypoYD203dsSW59yGiRrO7xfHFkMi+n3uPseIurXMHJC
ZCCRwJLkoiLnZiw7WNIpuxEM78df0is9DFfJgYB5Ya0rnthieOsMNEvJ3ECioVkP
AxwhJhH5Lp92nRFtbixWyaTrYXN92P/wp+8T8KareyNtBlaQe2b5lR+zU95mzh0e
MvoUYvwJgRexnPZRSOxdmRAxV33U+RN++RpvUPJd7mm4k6lIT/hTwwZdvOd+Hj/y
UsGEE6DLfuqFQmvkrh7gf7SxPL7rIzoUGNfpEHLsCAduqb1B4xGjcQTRxFwf+01a
FZcD2YAQ+E7WZIvT+RttHZkSL2kJDXQHFd83vG+aI+/uaaZBtfNbEfLyjNG2vTdU
FhoUk3bpX29eNenJ8tiwCxOq6OYAkVOi3ZI+hnHHmdAnCdY795MXjUxlXQqVTFvr
d/Yl17jXRarJPrCOF9A2xBAi7ZG1GNTL/Ix43LQvn3f/h7C6KGVnnwtUlacTNDwy
vNgcLazeFtwVxYpnnqbpkEW+2AO7904oiYkU08x6sSSZgivUm54wSf3UaE4+ifv6
PkY+3FbUG7ZHWPvyEQ8u8I+CJqqlQDBzlq6jx7YLfoj8tDtTHLiXygxBVXZainVh
OcN8UC7d6iEMUNnfLpUpi1yEccx90UN/+6APMSk58EyN45VL0VirEcXz2ETEaREQ
wvnAePzSsSbdzTkVpVLdKIpf1IVf0MnhM/KIDJyrLQ3A19PDt5K4dPbJXZ0DX2hQ
goYs/DqHCkbgCxKqLpC8FybhqHGVXzmwsl8rEZAsngwO5csQk8mME34Ctfj0NlKF
0aaJr08bhqy7FewXmn5jVJArSCLS4JA0H9s3q9sCi4UsyDKZOQhzoLsaUuWtaC4Q
j3HSoUtAzthtbXsDXIt4PGrO29hXjhZhDL6gdXocClp1/pxfH3arkVpwODfN/e11
E0m+SVks/h78EQnxnrCF9onId+bpad5QzDyvIyY8xRESDElUD5YV4YzPCGStx2Yi
TUf5ukefV+Dp4TPFeVFFis3kcL+4Ssm5r1FK/jfzD1LEqyvixuN9d6UtDXhaV6Go
Z8lL3uRmAMFlqyWz2iD60VjKM1Ln1MxQc558UIhT1uir6P2dZGbFqwYq7njL2CZq
OOcJ9e8bqjyfJCHPhnSHoBG5PFX2173/7skHaiSCYtOyjtukZLBL2Sg7P7+QwXki
SNfjHYak+e8cwu7YGwaCGqDeVZi0X8VMrG2xV+Ue+nTHcU/kH6AmKrIiNQOzsb7w
3R6YDELDr2ZMyrn334wIpgzJvQFQc8yjBDxYof0Mi0eygOLl7lUgpx9+FHAf0Lgi
VqSbp8nMqYlBo8cC34g8pERR1kn+5VZVxqoRAAU98SDpmd9jRr3ZBWl259Ri3KVb
pLd7P4BxNUt9DJocpZEIH6z6MhLiWWSYZsawZF4JgAjBFekWuHRiMgsjJg+os+Fd
RlbxikaairGcSBEkZSeZR54vb7LWAZOSP6Bsk/En8DuElolbHbiCj17sL1TofzZb
hEy8J20fSxbEFrZYcarGGGNp3LKZKNPh/pBmE5sdm7dhXsxJf9GbnLJQc2ADSIiZ
Us5ArdPeJ2GnqKrfSse6HxgERLQ4rXUjl6N2p7yQcu42Nu9wzDXaB7EU7bOVBq94
Ts/pru7Oj8kgsTP5wNo7DXI29o65NmZzFUl8WlJ2vr5wTRivPHXkc7nagvFRf+rB
/nZN7o0bfqjCvNqSD6q0qUlYXTE62ewmvIHlBxPxTHA4hYdrGDDhHSDUTfeDtT1N
Jt1Cz79S/9cqZZoulULCpaegzSEYr5dYYyzqLqeXAWa+ncLpkzuyvMSRIlcjtZxC
aiAKd6Zb8aUmK9N5Y54XGb5qEQwldtD5reoYsNy+YPLOsPFFhpoFIMQSFrp0Op+4
EVKPvj1kW2LSplXoWm7wEmExw/xlMdJYMSR0WXe4HRnQbUBQrXlTBz31G5b2FFje
ZRrdnYB9kp4GHrn5cckLgrLjVfJ5P7JgXeTKQwDXnUduRZyQlFeH/ohZoeZF8RMe
2eiiuoamNYjvMIex4+Q4cm+lnx8B6xYmzb78+QbxFbcjHZzB8xjMdxkSuAfZRb2J
3ggP2l0ydZ02wKr1Zwmfer1PJGmZ7NxbB2QWWdx/yuuzeDQywbdCxiCXMIKCvJeF
C+4/hp5ldfGwoM+ILdrO6RICv3wOOdQUOg+Khac/qeDN5bpv8ea8WU5KGNCq0CSl
0bSIsGbspMfl4NqwfKBhkbRg8R7Wm10sTwp3RqdBm/Iav8M9uS15suN1mgv0GQz4
bxGk8TKm/UZQ3JujUFHk40R9Rlbmlcp77ZlF96E5bf6LWit+YDc5lypNgNiuuYaA
iRZ+i8vot5ZZ3gGxR5lK3xwr3/C9x8xLczK44mD7n0VJQLejt2yJgedr7zF1Qbgx
0CF01uP7UecF4KLn5khJpSNJNSWhKsSwHlP7IjkmSyJ+lC6TldoMy4w6uCtlALYT
8phmnZLDgyj0HAwwmj2D0pn5UR6ckqhZSlM6de5HUo6P/d7s03iOEcipIg+8tjXw
ZLg8cK3XganWr7Ssrhg+Inh1QIQ1CZOO5qNoZuHyhhvDjmg07Msb0GatcUjDtWtI
1KIhXGjM77XI+24DCVZ746VnqF90kiwvXG/sdlYq0hkZ5l/dPuqU/RRfLzm7yHss
4SiCbxMBU2D8q1w9S/K5I05dLpcxBAVXOdtc9yXTnmwyzjAU3cBjmi1wtTgU2JRh
WiBJZykcDJrOqyGl2zqzzxyVpniaEP846ncA60czJFbFJOudySYs0aHf8yDeasnF
1ieFlTjdvi6yasyuvUMT8nqfXwW9sBdAACHBUUTxWs7rVd9FvqQqoJWkIAOwVbbm
vbkwSEU1Mm/6yiKwhNxEywBxuLoTZAv25vSCQCiKyp2ZNv7ayNdnv3ky8unKCLHE
5bBKeCZ/0VBXz2cCRXbBQj3e1ZSoAb+2qy/FFPA8bD06A2OKh6MMsoWi5w7bGCBY
EOrmX7Rl8K2/8VLXVqUkbIH77MjfY3ED7MvGkzgw9SWKNvOxO/pBNmN4oLHL3Bxn
Cl/5mI1QD899JbJ/TpJ704X1HkONpLzDRbnyQNG+zZte6Ni4SJTVxTdzpd6wExG2
V+rsKlLL4WYDOV92Ahnxe+uGeqDvvhAsCZ9zQtBPS6ciBWAD0zjDhrejldbh0dW/
yaOMXgna6s7KfdtWzP7L6xG0xEwxeHvF0Qb1JQE1qki4vI5B+EaanxRmJW6zZloY
wzvEGc9GwblNB6gwir8AKHLy/HagRv6ZuVFbeizhCMb2ScjsjPBraQTFnHnGLyoR
3VGME/Ft0LvF+YMbx7vl0ygEMwOiAGJzIpKbc9L5woUoDigGhbPQhS8JEx+HBoLX
4tSV8R19BaTWJntVnGZbRNiucNgXsudC4DE9IZHB9W1PicYs+Y72twy3uIlblGS4
/BI6zAIe/EXOht/lpr4X96A5m7/ij0TF8yVPXEC5Ku+ayz7R/v6ADPUZ18TzB2eK
fNCwmA73V5SXHVumAubibFu9EJbEnnkH0f/hxNcqJazb/Nmt1U8w61WyuY+EplGS
mzWfF2MSYLWiXLpWyWmdx5u/l0iHeh9YtVTyc7UNbUTSECjry2aMgA+tZz5WVCzW
aUO859oVuAAcwQJjvxRMsDboH1gPJnoJYyhx3ppzm9I7Ov/qzhFC1l5cS7O1nEl+
9h87a5Ezi/KOVDFfLWywh053lG1A7jTFP8SrMHtYfXaB9+c3orERwttGVZh2zN+6
CxLdjf7lwmIfZNLHDs2h/zTMerr6zXgQ1ue0rEod14gD4oTyUZwgWA+ABHDqUXdU
7qnobQCV2bDYXoNW/QGaxFwPOxbsChAGbZbMuBnOrnfMa4Kuq3t1h1qD+dYzwWwA
F8jiEsvVaHfIthTA3edsuEuLTtdeUN+TpLbemI2zdiBs/mspAgbP/xmOKig44HYT
dCuWBCaz+V+VTkpWNO9x3+Dv6HqainAmJAl2Z1Z0ZzOFaB3wEXINP3F33uGj86Iq
VHS7raWUT0xpgLeuYlUxgqw0LX1V3d40GIUYgRJGXJiEfChUM4BYoXCWIBPraUm+
7CFmZvEv/W6Memi2nbmHSdqq7KbASDpGNOpDVxmqipnL3yotf7mcQGj6KyP7IKNk
oUJ4IJGujxt0wWpS9+yarB79pw05Hvgk/RLzyIbrGQYLSMS2PanOQl8m9lelBU99
1AzfLnXeX0ChsTHnd3tBFRJWhjF2oe8EsJDoaZP3B+WbNXIat036LJOcX4uAu/oR
MzY/fjfbEiZhR32CvKtKxj0PhxBWAzzu7c5gKk/Jxsl0Q7u3j2pkwuMppmYOpdDd
TxmwG4kdpk6zReXcHP5JOCEGagCUMwxhoshlzB7i4Ioo5fmv0eq9ZC7CrWqmSSy8
0AmX7lcj28vjOkrMY6FTbIPWJBNaKXz3z4/rR6Csw8Xhe0wytmcJoZIw5u1ZkIhS
CY+gJFlrrxP58ZLsvrXv11QMLgsPDXH1/p7f41nJK5OgOYuGfhnrmjinJtIbyKS8
CExn3vem/qhzpx3sLSHu5SiIlw8Y0cBHW4cFCFlEW+/RLmRkQYLmtJJ/t0vNkcZd
OVk2p6BgQ27aMlhMxhanIdsTsvg+SMszFxfsaqzFazOVBvMNtjH2fWeleBrGV9Zd
S9fmNMcSkEmLV8CzVJUciK1A3y4n9vGzZ+Nbm08u4223t3LF/ZDmK47G+uw+qtXX
tgoyjvUDc7NaQSJXbimh1J2WmkQe5tIrcHlI3ypT1v4ac2Hid1XOBN+zBmqbVqQQ
dM4P7vo0Tui2K6J/S/cEm6juMt8AfIHecjcAs72pxDq+s9Kjd/ikUdDdhRxByjhw
f4kyk1uNQrU71AjEe7m/zmCrdVW34D0JjGUSje969A2gwT/qygUiURT461mlKN2S
Uw+Ny6oHyMZOo8teyVfqEV8EASuT9M3wJMhFf8LmKY0d0SCXtGYvjDcfoKqcgaCj
18PCvKSjkeaItgXPRrGsNVuAQHVOft2u/riYn5jiCqkqHd5SDHlOaWM1kooc2KSC
pxSJswSC5nmngdE++RxSHjJDG6r9KqcXFoQrkaym6KGlkv5+sfbRIKKDQmovipsJ
h0YjWo3cPNyouKY7muFZh8VqvetcWb54e2j5orM2Xe5GeyiatGDfZTG4ihN5W1Dg
Ob0eTYHG3hQb0PELBhgrs0tzPEQhtj0ubxCOV64NuCREWgv8FDj323eSXO/7tMWu
KPE/UQcgiUZ3bm5WTVIGfF2TUulT0Ka0v4LkGb8CQnZVopxfmwvhGKqVE2+1TsUc
2jfbRpVAgC3B7dXQE9UdyId1lvI5J9bsnjcVI7TIE6qNgcSCS1B7jWgrA9FIJHjK
I4ekUEu3mj9oxPGrGa5IpJWIKXZWExwP8Va5yCPftjRJr7txd/LxjxtVzQnVtIMt
f0twQijfztBDpWc7G6b14hqW8+BizdaUv+hLq5fswnop+t5Ju//vEI+TSW3HwVXx
F6IgFFnLBaYdb65xp6M27d32o8UYRdbEby38rIZuGvuJTbYGJXAab2jsYL8PeTo5
lDw8/s8IfT6Wi1LRGry0gMzhwyoTdZduAkINWJQ3EtukdRQGnWmGroNaHwT+m2Y2
hGO71PwkXucfDXLRzHQ3E0HvI+cN9Ysl5MfQrCjFwTG3RmVT72ok6kpUGSZ7O6FM
TyV4tC574wKK9/g/HyqYjOVmv1bPUqHCWm8kE/j9ryty9LQ+kPQARlr+JwOBj2Or
3uzzoNkK5OAfQUHkAo3SdUDhfmgXzXASLkIQp5jogJgjzq7Y8oxPmZzoG39Wizax
81jMWQ9eHoK0sw/jGNj3JOFYwDc2EOOHmZQWiA63XfwXomlx5H4qpIZAGpGc2v8B
L5AtlyYwfnmNMKki2plRrzJpn3mSmjGg+utJxO5rDztl8iGByPRg5Kp3bFTjCnTj
NQ7Uklezc8yx29a98VCw945hsrlo54IMEm2nhpLCe1RZbN+ZEiur7OBNUkCINjQD
76wOUUL9tPY8JnYB/Pk9MdUgwORJUQZwebZ0JFCtx3ybbQTZ+KIoPfXHVuTpHybf
nWWLa/ttb39HkNJeEUv1gnvkrfduTlanUFEMKYAXU3NuUTPraGq7JmykIG8xVV6g
EIZTfXE5zEsd7bjAutR1JInmzcP0T6vlxsMV0TZbRDj96VCE9tvEZ6q2451Tf7P1
9samA6fM5rAHqifvm874gW5UnMYAJognGFBagRNg9TroENljY80nhJVp7Lfecs5E
jFMHP3XkUxeh5L9SkBTGiczfNhMWyU65jiys7ZFcajiW0DhNemR7KXBEmOhJwwn4
hfQvsqJtVkxvH/S4s+A4DBYVxyyEP0GHTVyIJgiWoN7V3AxC+IWuzMx0jj756tr7
00j1CQtTJIDiMPsZ808TI3wozSZRXeHdodntXZb1ZaUCQC3ZATiL09OgkPfpj31y
1Zs/OULIlHRQQWhC5jFHKuD6hUyfgqJpz7wxFjr4a0HMASM3ZfFSbrYfwPmbmxPW
7uxZ4xdSp8YKGltb3WNN24c2SvsQvrQBwxqNs2CaAMXaaxyNzWji1DUhfFte/9Y2
qUyTrFb/MpGanBFro09Zso9hhuQparDdrCC/RtgEiT3iAggSDsjI+1eaZO3ZycDo
DgVACnvgyInO/sbwI+9C8+jvYP/MFmEdkSS1G7Z+Q2XcCzoYcdLLxT3OcdS1BtYv
P3aGBOPsF9pJ3STFMW50mw9AIo0elwZDVnjr+cgOsL3fkf3k0EKEghVQd3oeRsWC
4HB3u+ep+SAa24W7hfWKW5ifTPCkbiZgpTUpTaXLU/xIk4T7C1HWt+Vlom2rYymC
x/hSGu9BJHU+MgtPKvDAkFHbv2wrNxuLrAMGkf4E44NWAFvpM5UB89EkqdmoZak5
U7niIVyLJ9W/YuHoVfipuGfo/W1UlCVE8gTnbEXO7D1YjjqmWTCXi/8X4n3J0qN1
7tfj6sLMCi+D9Dsw6Xtx3YRVmb1DpJcT9BbM+hM4NzT8p9zJo3f4dp62vL9MHg2i
7zA+smpWlNITfvbjhb8vUksc2QuhEIpNbTzVBOyvgGrDW/Bxrk581cGifnX0HMr9
RpiNcKA+5noXFaita8EwfRo/nKUf7DD6SMPDhfvaOfAwnBrQ7nl6n0IWyZnTXrce
gFwrP1NSzE3UIkPhpu8qU9Cy2ERgRcUUqdqLdWDYvKxhwncBWFoiY5jJgI4+U212
dfTDgwhs87Y6wrX+0VJI7utWXNrCnRM91tunYAzoEqfY0SOo3B+hLPmGXVt6MLTs
o9WeoO5AbMupL5FRUxZ8dcsSJluMy69vfbrK3USroLoq8BQgFSR6Q7dhx6PJGKfc
86t1VouudOsjxgDifwfuXILUyks/rdLqyEU+UIkw9C6C8vQMbM8/3SDyu4jaYzKz
mCmcad00tqgebHnyddTNsxOSX72UxgaPhrfFhqt1eh7AGi/T15kcHRyXXTNi5Cq8
ZyKYGPvOTzdOhIayejlZ0St7UAE5sIrxRaTmemYBUaHxQCcMz95IU6lLOsqOMNrB
8CXdp3N58/ZH6xUgP84OB1cJDyfV4/Kxbvw3STfut2+z+hJ4ExKOEYWMiI0oJUXn
LFvf/+D56wFZWie0g+KN2GtgogHNssFvBdF7rsWLlAbhBMgfY6LksorcO2iUUkjk
euiGvWVsvy2mLKkdflJH63Fo4qFaP4tbaPgfpwbkzk7gyuQO+BYfVbsQ8uevNd9R
ks5FRTfipO8UKdGhHTRcjKf/aoTfIa+oGUpS95xqO1rrFL+3fFBAKO9kem0A9VSE
O1U7Sas2M5O8VUPhJpxTThW84RgBDiTikkwrBK4ElHgRBQQL1FtjWz5Wxx2LHSxA
ZiaNa466pYSg5PzHXw+zYlws8aKE+vFyWnJJqTPtQ1F9gLfiD7QsokdUQSLWj+dx
URsOImQ8lwZAye1qqkvhbEppQEVKUvurJubpM33dcWyyVatSazdvnIdOkvri+6XU
MnT/3CDkSFJeSa87zRlIU6gl5+tOIQW6gNp6kMlJEoP43axPaQbT0EIH0bbAtTxn
+PkMBgHxLgi/6meQk8UMEMu/TjI93UyGWTNgldN6OSgkSXqD48VP+Pewn3eeBXQ7
dhkVmZWEKnWZrb7li+LKBDfDXy/WiqDvDmH3/tmJXdpXjvIC5Pp9loMXx6Xg0Qhp
UfQM4zEgp24CYKmbUPvnFPUmSh0RM2DjUZRjyrEFBQiX7h8vpBBUt1UfEZrAkb0t
2pU0J3HHGfjtiscuq6LMzPgRX1Va7z0opfE+wZGWUSNdbegZitxRJpvk6fDDiLL/
vtyzgBruxuH42GR75T44iRQ/eXCfAD0NddWzrmKUIV7VtfbY8EXm11Td0SQ1d/ty
hmqwjXfHI4lyFXlQCkC3TDMSVoqZY4te45etEGCSbrOCFdzvSFhqjpCERglk4wM+
ij2OkOsEYJT54aFW9oh0gbOKQTTQ3rsxa3JpXMGETMPG6OwTmUOLAESz/eFFUmsN
7FzDIF1v8JIyZeujnJyHfdAFXShVuuIh/HhjuDzr1tgIBUnL/p5ov2AAcDExa/pG
ZEpGhG89F1DJ4y72cZawb8Gywhm0rRxEcORD3YZiQBNCw7WGSHitzcLy/P02tZon
CDnR3iq5zVYWiDYr0TztSOXU74iLl8ClLKfIRWVESGFuZTu2Kr8ZBNwChODXhEsj
3v3/dkyUNm7XHW0nlsXgoun7kCVwOmWC2r/iKhb3gD3MUD1n8b0rIyUba1bGmZ3j
zMGpqV8hmSLT9T9/pb5hFBf4gZdygECGZnIME7tRIgaeSi6vPPXopCrdf/8iPuAl
kUB22AjGR9VbK+C2/Ev/oIMLF0NCQvEri8+Ancok/205HEl8gDhB1Fh4Dl5juNYg
oOCTlet6PuEPUN1LUy6RSHMvWL+hg3TkCyuTff2zsV4fdBwkmSXeDnUZuZqoQ1oj
lHuBmIjkZiawwTmQJ8BlKctzZAPu1J5k5zlxMJudHxHi4up8c7D5H5aZvgUgWN4D
/ZnIu6F7+jQA1WmARH2vd1ErNQgAA8zXIwkVf48Y7TOsJ2cuHCwKZulBhAqbqbHV
lGGiYYK2p0sEve29mkXWWDNr5kMUo2ehSbnO1xga/BwuBHW5Gx/uT0+WFV0gf655
BIeSTl0GPf/ZLTceObTycu+JK5U4uGZUJVe48bAmBzNRMZ97N1E9zKeuiPgScTzL
6oBPIFJ+gCM6i9vW1w/6/qIPRIRH8sfwMNjqblZpVL1Ku78+zkZSUChcu+xgafPE
r62Y6TQKlZ+x2ndgDJzDWERkZ+5gjA9yFnYCtlGGRmZrLeBqCvyG+vlOZxQv4FTp
qYixi76jTOaak965Vfiy7n27OWhY9f/vXUAUKSCpCEN90j51p+VkTRR3Y/GH1lng
W32MLCBPoO3RJ2KdRgrN+46Ox8Zp+mfsy0PX5eCy/WsYiXXL5CPA4XNLR91appWh
Q89x2LU9F2hVQphhnsQKsnmakprM5z64UhuYU2/yqj14UwwqmSy33+G2kPMcPfQJ
sN6yPDWbPN8eTbetXFWHhcp63h9qKcW9e4kFgSdgp89AFM99e6ZCg88y3j3SzMW2
exVR3wy+jfyXog4jmSAKwkeppfrNfbNPzyT58MJrNibFYlpeNDkS5fCHOrgSN5Qh
BRkOxeLKMJF8JvRaaoaUzpSbzhtlsCOewmBsDzJ+AI+CB9mG/ZlyhaZYTUNTO9Bq
X/cY9AIM1/ECcwCQJucAHBHDyNRQmY7xnXu/AcPxIZsRw3Lt9errBtuUVb3r3PeI
x2T8CW+W71717/dHGyakl3KJmzDs+ylCuA7a5K6YJLhnAsv8luCSR8pVQ/8posGU
vucLbBj2aPiFkXulIFBGWV/3xgVGbIXt+qKK7emLabGRuUQQgi14FVYF84qsmk9i
Vv/vNOyi1/vCzorifS/3N/G2Mq54Uh0EVgNxOgIxDp57fQ1iCw/+u+JKDx6Igc+8
9RrlWzZTGUJav9t1x1vJPK+thf6CgiVnQUPG9Pk5ubjcpwaJpRVVLP8dWoLV4Rze
9dHDS8sQr+IUO9UtsDK1CnfGThGVtW+ZPwG+2SNKxnVQGIN5k+0Er/CnYH1lbFWR
78QHrLbYNLALkd6Z1axeY8JS3q2ZPWP/fLhGd14058IY71kcn8j1kXv4gI4ofsJO
S9wQW1mSNE4G81DFv2MagqIlwa6XCJ5i/wwWuf6JUetZugppQzC+TpZ9H7oFI5aO
iFT0D6OCRhNZb9vHlOkOElMctqwmsuzTMqg9Q4KWz8grX8hfevnMVpG6/wfpi7Q1
1j1CwX4+4kDXAaMGehdQFyKk6ri+XyfnldFjTb8kidl8tX8/S8cwyTMwcbN5gSOs
cRG/9Gh2cSpD/1n9FVpU7Ej9wD/WVcqDxDQbqIsBHSJFvyAk8WBBOqJ+YugxrEoY
Xy/yrZCEPqvzQjhqRlOqVFNK1gblAaIPNO0j5osXCJTQQXPiQS5uQG8AmibCix88
L++Tg+6opLEBo7ynQnpX1hpJ9xrWrJZPOAhaxljv+mEeADeKm0Y5ct7+KtVRwW88
kZIxluLMWsHnXZ031S7SlFYBRbqa6UDYat9oB48Yeq7Aw0SSSfO4B7KqhILJDkPH
+fY1IOqsu8g8t4Mver5dZXpucZncswwSKb8Y3wF5A6RoM2w2h3YLRXFeo5SmUj/b
9QvSqunlFwVRNAryM0tKeJ2MHSFGQwxp8NfFu1+lJVc+X7RQWG3QZpsWSsOO9lBH
BNIq9RZbt8rAbO1Nt92NXKEYMU6Dg9NaC5sHZk20Yqslw6F5Zg+/q+r4+soyAiT/
9rx+MP0SLftt+LidF7Pgds3qdjvcVto/MhdVxvmj3vvPuKpuk7wqzpl1yrNeMFcT
CMFP3KfgOleXJo8wfnxjeUYMXfxaJgl7Tovjq00bA9YTgneQJ3UTd193n931QYgO
FKPabBAT5z4tJduE2bpwHNgrAIC4k1VgN/D7Y7tfWwiKlSBlsIY4mOGjULu6fBwV
CvdfjmDK+h9jbir1pfoU16MVLDvMBtv8jsbIk5jmp+FdAUhdFza7E31GOxiyUaa+
Fp7HvtBikeKTIRtGZcBMqL380OxVSrPjtIwlGGwZdZSjryJe1QhxRCl+8ryIHkFq
x/f76FFvHmSKiekUVaVdi8LIgJYREIMn+ai1eLWpFAFzsasixo2XovPNvAZXE5ZI
DZA6QgfJ24LRrc7M4gxZi+8bPWLd7ckqHgTzQcAG8Zm8kxpVdKb/5pfp3nx60cDv
KQBX17kRUxe+JGBWV4KuCuyxDgQ7P/EYe+NBJOwgc/4fCb28IIHY9o3Va3mII4WY
EN5pra6dRObiN7QztUa4orIuaXA8lVIw+47Qlgy0lqKnmvfiVXcEPgAiTPVn7Vg9
dIsRN8SEGpjeHGyPO6QfIZ+0PYrQEYFr4PAap3lCPRB+WIc0hxCvRi/Q67/oEHcN
ZIsJcRqTJOFgAO3WiypnOVTxeZiJEVaGUSQH6ybR6HCl0wa+vk3KMsWtJqaK11cz
HK0h/Z0vaoL/d5KwrDAE4IANZKDhwL2mfUs/vUUTfnUZ9uLK7zjIGMNNsKTN0UyQ
Y37Hj4N2w8bsXLQAKTuqu/bbZRSSb1zaQSAvVLBzygmdX9cnTjDmHqnnT0WtIt1D
e/dyEbiP02wcwEitjWYhX9qdWlqNaUnI8zbj3fSo+rZiIjfeVlhKxI94dKvACpVE
9sC85vHCMHWODOo7PbhQ6wEDRSFX3wY2KpKG7jpsVPqiq7rS8KcRdO9JZggRH6rO
yfh7gGK6Wag16PGVaAH2fxwX1y47/0TssbmUGosY2PTBS4NFyu0rbo2R5OKTTv2Z
pMJAYRJVjzHF5AUVyC7Uyxpb7uZChgoHLMP6Yv7yGuSAWW3KZnArXVxUOSKVcnbF
uX47pUC8Ub7pBOf+Pz1bmO4GecgKGTHnF6yXyKcKdQsWM0bX6znx3yeCqgaeI+le
GNmYBhRpLnism5U8wwgGhy/CGR3kPWH/I3yOhblZymIqtlZxehEVkMWy7256u6L4
blmuj9cNDkprb8uLri7tj8dqMbLlgn3sq/LG64g8oG5JehXRx5VI2iY2bfvaCw1G
ir+UzXhhSwwAY71RyvQ0/dGn89t0ZziVsyzaA0T988wBn0qDAnywzeh06xLAexJ/
ks8ERXXfUoFavl09MM+3HjSF0hlAl871XeLZaC5rrT2mELf/jIVxniUfEel8kWhJ
PnWWiJMWfh6eIvNsvV5eUNnpbBrkJR9AvIRB/8J4vnM6KS33jn6c/MPU9kG7YCCN
rivnDhUKLFtje2bpML6+XAYauFEYAafazlcAnH3LRCECkifxADh8gYBBvM2azbGq
6iM6HPbIXWEVvYySSKFKPYT1+kzQJGE3IGwcZ4Eq8p01ItKK5mWEHP5/bja4SvXA
ziVw8cU4M9KOKivcHgvy5dKC3cnRuYFXyCY+o3tLkrN786rESoZxr7nuoYnVBgwe
tDo9oWs3zVaqMFEjIHlJAmxcAyhp8wjnFgBQlnJFC1MsAGJhvUHmGkGLmuUXeuH4
UePFwCF/YVRkvuLrGDgvzvAG8EJZgZ135zk85FujueyW8wDbuqSgWHhLgyysb54g
CkM5t5ORJ5yKVFX9fePrA2ZnOqHfmtevALaTdjtnuAd0D4rTU3fMOYv+lrM1Z0Ln
KW3fK/DJeE3+ybzFOTZGassAqIBliX/IbxSKtpER5ONs4rtVhS8cmVqq+DbevtEu
phW8m88BjFsqx7Q6ETjQ/1KPQG84R4CD/ktMUSjusUdPT73lqpNvM5n+ihfPopw9
4wfVnsuPc+siAHVcipwFS7qzS0wgBMX5G7coqzMWRl1fsfptlAYFNw94m/T9S8gq
bf3MFMsGgvRw38+h+oqWrmQqszE0cj6vB+nd/9IjEHWTILb2tUpUzHUGKIEK54L4
q3m+TRe0UlmA5VBJ77Wk9GLUNV0ig0Xfl8QDGphQBs9+HT7P4RDJcn1vYYxwJHBO
W1bRcXrsR0dUKgenpc1STTlDskRs2LPLIuCOZjSVschUyPxhDSCQ9QmiukvcSN0n
hBd6/zdBCx4sqXcC7/hv9241wd2wczLW6v/knE/8MzaXFJB98ExoVfRuZ3mi+SoU
JNfzmcVi77SCvRVvWoeNg1qvb8SGy7OvI5gWMvn/8cJ0OMjC2RyjztlAIx0QgwsA
z7cpVEN86l5q8eiJB/cISdo6d/8+RaySKxv34Z81S6r1XMK+F4vhBqj3JxHSx8LN
VrbNUYA/GAAhi3SW0EKeMHrIf4fTmUiAUI+CKegWc0Km8Y8obh/cjicDsPFjwNkA
wG9p3/7AXmNWvJubWxzUp5qkdugV0MV1Rxo95e53mVD8dcF/UOXo2kuaTSMHp6cM
sMfjTWCHuvgEcQm3cFdHfwydNILUsRyuQDDJmwmi/mKwaPZzBTANcdqos+wI4Fii
x9IVEB0Qf/FmLyrrC/dZHfLFAjM59tvdDUY/uVep14UvxSp+WT7L92g55VPWKLi5
AS4MZEvaw8UF3cZl6swAGyEF1PkHzyV0QjLK0RYAdlVjmXbNAYpFsI0LptXI+Hd1
gWkBFurStVkr/c842yZ+Xn7553SqHD5mCnhNbVUnxcx/YwLk2NgVazMD2iRpnfF/
REwKO6IFIKN7LMOCkq5aqKJ0WuLduRt5s9PuduyJdqIRhf+6rrifnpBcq4/KOYwr
jzwaCWUYX+Zy8dLqZSlHqPzB66Sgs/fYKs8i+B4d9r/XKHAUBdUgrCJQwsdLNwPe
7sIMzEmCFWKerPwopdLlmfXYb0dPxv0hKEpU1CNsSTgOQ2ePuAGuMxMwkM1EK+rk
B0hSmvPyVslGa4hRzdlD9dMMyKNkh2Kxd7rf4ma8nigxjkngW6RbjinIn0du3U/Y
CQxLNAMXGVkJjWL+l4G6ZDSk1QMhsH56fdijKACG15fUkKNAqQJr6c7S1q4QQJyJ
gNQCFEqKDDbtoBWIeMYxY6Y7v84bWJdBp4hTxIe3MqrpH7sO/Ik8iVFwsWQ3wg9c
XgNWlyv96KWeoN+tUxCUMy+1NK+4wdlaAiT6V9oGq7Oy0e89pWlKszF3yySxvQoM
Ur3SE+gIE1hzeggCuo2Mg8RFAfR4xT9K9MetxnpAd5Ff5vwLKl4cKFt7E5QYmUKw
SnEEBQL0GKXHGsMvXk0RRzvtNCpLcv6Q56gOqHXcBfnav1XnpMWrlEG0Z4qjzwu9
zczG3XaWof4O2iDaweg3ZmZUv8jVc2WN1IZ1g3iZqz2DYkvB8kar2gP7A0B7lPaY
5vNpwqu6t269fMJFw3RviQceK4dtpl0r7WBF768vTgulR6pen7zQ+Ntj+NsewS4T
HE/5n/g210QlM/oNdJMWyfyjALUX7f7fYPI1wwH/PQPbLppUwlBJFzygNtgxToMR
U5tppRsQEUEUNN4Pw51fMPHtdt4c3PolqfdY6ZO/ZII5nXyMV/nEUH1B0eqjIcps
RXy2AG/D2OwE+kEcCvpqPoOOgNSbX2pE/BLcyOF5uu1Le+zADa5YDiRWVS2ELSkQ
CiK6DVJBAHQfKSJ11sizvV7mobPhsuXQo9SYKJH0rtd5+IhsP1VjtlxjDN9hNpyN
9/cPRfJ4EHTugXsuo8rw0qqlhrcXgmHPFdbfDETo68RaKWoPQGZ/hJgCcBccUtg3
YvqwYA9aWdbouLBxXaOE/P0Py6ZB46/ZQj06yXLNgKrJzc8TN8581yvVCQjIjY7j
efP3GDA9jpUu509n51TEZvpr2K+Ij9LUvPU2bhZgKjyZIzomnc3nIeGMS/9W8Bqz
+70VeLYG80/8iYpE/dInIwzl3z7pChxofrqmeapY8pESpmL5/CUe2kXoV9rSxjjc
fezbaERRsSq8/QTVGHb/+vQ0FbQtS6knDsLWgecIeW7cxsG1mcL+KoIr/TxZULpZ
pqa+guqshVLGA6guJN/dWzmnPVaGbKPelJJ/4ZOw5Hw//wub9UaGhzqjNjv8oMbi
k/Wbacvm3IcD+b+dBOqHMtkur8OjhtwHG7l8VLDudiBMGzDbD/fgy8QPIH+RywYf
aH+reLvtNwk/Qy/kFgGEdfVjvy9hnLF91nNKvuRF2N2eYBtDAfksZHSPZayoiS19
Uw4vA18qcX2JW3F/K9931rA3T6EylbPJwiWwMJGBrQ50cYrGb7zf6UcjLHCTTtmg
P4QeHoO8ZAKH5eniGKqNbc3E29x8nov8LgsuIMKM5k2dq1+DItXez7zDBTpCA37z
u4HFwGMD3FG0oVPwzimk47u9s+ZN/YhJLf7ghP7KJznCM6+qWmRht4PSTXaknBRy
+VRVT9PRQ0ipiZVMe+wa5Ly2MKYIRbNxpgGmqfKmpfZz5a25SorMo5qW9jWe5AOq
34RI7yzYVr3U5GMSR4/YWjfzg639kFdnAKbqwHxJEXi3Rni5J/WkXY+r/D2yj5hN
adP64+WYjL+hMt67vvcEjGmS59XxRTTV2QqKFZXdKh/ymGJOQNkDZNk69aQpA3u0
0em3MiGXhVKj2dUI5K1iU9CKDB16K/WLfwhIKiv1FVKa263c/4+K6OUjxoHjNW9y
Jj0Y5DPlcsFXeooNLzTMzPmXeZ7WQ2k2uncBadwU+AunDK3rI6mdoqa8iAtFlQ7T
Tht5B9EX3YaNrymeEtccfjnFKZloGKY77lcHCbH/51+uqYvNpUiCuWIPjvCQv35A
n3L48c0MtmPDvDkmCvVsPtAKcuY/GpPyCKA6eRypasptNqKVFtARTQk3fKi6V7BS
7u3Ph2hVlTyOk8pUYGRtjcDsl772otaZm0iBuOVvEAUKuN4K3hJLNr2U35XIhaEd
6GX7aLnSWnwTeWkBlBvGIJ1agfibyEQFKtAChS4S615ADf4H3QyasKIiI7wef/eE
wAOHpk0kmyFiDn08ftE3IAVvgWF46g0If6lEhNEOm1fmS36I6jkAntHQvZ6/A3/5
smWBEj2XZcWkt0ObYRw20O4uUz++4FNkW1ixnUaCcFiYVwb16fSRqygjTr4qlHny
Xs84GcX2waOGnkyA7rM/U8u5R03HrFzEpBd9cTdn1gnnLK+n3lexejReFgUqwqcM
Py+2BW6zoe7oXDRG/q49alhqq81TfQodiVBq82/pC7qnHFhN8E51H73piibSa46b
xCjcvpzqDw/6C0Rxt4rFRcuUc/JgF9cpRjTw42evgo7A1m+A/oEK4vP+dvX4XYdH
1/ccMAiWwrlybWbuNqtEPRT+SpaeOfSwaRFgU7D40sA5N+Eqcn/lBZb3i4aHzeXX
gMdVe0MPgIlK19qAOgQW1SHcTCHlAjYxVbE+itSwoRsprfxyC1Y0REwmAmV+gyFb
yFsTVvJ3qOyhoLk1Rg4XgJjVWOFq4bncp4YSIg55/sFlE6N7tJPRMMshj6v58wXk
j7GWtvmPtdDsE2Y19oMQTFoX982ZMpskzX9klRzHQK1M18d9y2NDrWhdaHZy6xza
iAd/SdqyN9CFv0npnWQFkZuOQwtovq92asaHJeJt94d2/TBZ6GGlOEYUR7jG0xDQ
SmnFmTAYmJ3mmQbNK6g3SuwhXJ11ffdpwZynmq030ZUmqWzB6ucCQTwNf/e/G1dn
HF49z2swjYBUautb/HuGQB0XnbNeepBWVO+bD/wMtBnCBTfou+0i2QPNIlPQwo0g
fWGJLQW7sFh3L7HBpkvqIp47kQ/N2zUyqZ+b1hsNqVUvxpjFluJLOSR75dmQCodA
fHIqBRAvayDgE+bkJChFxyqn7npy2gMcjSSMsWWgd6TDz8fDEBs5ygmZ+bkZ/gTd
SHLTpgTKZuJ5tZlvzk5F63ULD5PwJnfGXYdeBGGwk+8Sh0/pStGg/+LPI70QpR+E
G06kZmC9u2WwGVcyDOt55qOkIuemdMVducElxRGB8XkrXa5HBfQ0C1pxBfxYCO1T
Ct+HKNvhtV2FyFZqLk2ESTOQeLnxli9oX2orhhjl+hYTXgYwPQHZCgI8tq3KkWT/
P6Ski8vI/BfFMyhlaf/gTq9Qq02emZfxHyz3xN/Zb0FMp0nCkK1CoYoZwvWXKmbc
lX8+6I0Zbc1BGohiZaOlE0dqBJBjdNb6oQKpV6ilNbjupDK5TBSTVEkDoQbsR6W9
J7EwfA1IExF8f3n9TVxnrzEs5WHZst3RDX25zeP8F9oTUlW5EkMomTZgoTaKN86n
L9WH66UkuZwzwn5qyKaxBmree2+mHSchioW4u34veGY8LQwysDTDNtxo7Xv36xKt
JMtnjnrh9wcJQr9cmCYc3WehZns1brIjq6c2wi7lYJb7ol4Y9FSqv0Pf7Ts76uDV
1EaUnyU8tKzYlsuG6S4iztuW0Ye71/QQqFu4Lp1td4NPaiHj5VBvK3+cOxDKw1wf
9FpAkICdmRpj8vHaxVQzYaRmBDg1r8TrjQWUhJgnNEXUoy999ikLFNja5zhhZUdY
+gSijUxHUq6hJLY1Y4x6pZe6fhU35RA3r04PZVkt2hbcbsaoKmurnSumxfFux1Ch
AcyjPwEDQUlB8mozsifVZbNia6vkEyjQHCYyzq7UF9v6nrFU9j4Be/7pr2ESA546
4XUEoxwu152PFVrmvHiIpDLXsTeiWVPpyphVQqk+k3qDgA7GBAmKvJY6/5dvy72A
pBqKjZo5pCYbZYORHOqXw1ON4Pj7+NTxg+M8+mtRk2YIU3TeRAqw6+4uhSByk/NI
kzSForF7x65ochKWJcVzJp18zmhn1c+M6r0U4dzqu/7JCNOHIjW9RDA4SF7U3dPs
OBX/OjnWPVDRltJ20dtSkDazZI7Iykk9TSVctL929NisSmo8x/mx+5Fe7/b+9Z/z
UO+rIzNBukzlMGHgEM/arJOPl+xfmeBlmlRHiwY8lYmbgmJkEiOYYqgoRAxyfso8
s7UIOWf6txNN76aj6F+urKD+U+0/H9DXAsRmJcDPXxfCFVG0DT22KgI8NO3XzQcE
0jM9fBdK9ICKc2crvQsiMx67WYxq20XxXMY5bwAdha/dIKNJHHwisIt5ZRemsBgh
uAnSznThwBvjjDX+v9VPGj1QlYSsZYar+85tpKbmsgj5sVyhgn/fnQT9F4y5ayqN
JgkPx5Qxi2luY2CuEUKWb2qeXIR6fQBHpPMhRTWekGfEFUzDHW2djdv1h/IGa1UG
6DOZT6eEfPCnRZi9/NN3h0qrDjrLsMBfzDiacIiU3nrxJ5+Mpv0zzPxAR4+aDRJS
/MGh9h7hsdW0yRZkcTABy1QbZVBadsNk+Y6LApEgyVuqUno0wfnuHpUVXQ7Ygkpg
u9VOOG5xy5m0FV7PmiPEw6ct2N9SRhXq3latOqSbrGVHyIdYPgXlkr3mlCVm51ol
wuITnJmaW5p1JsXS+u0Zi+JQdOLh4qyOPjFC3qCCeBs7ObsLZvBva6lrqrwORJQl
6C7L8jyh3uz1F99+ycD4sZg0z/knNq8miOBJJ4QEC0Nr04EpOs5p92MibHFIhocx
ZpM/j1xqGj8EE5QVIM+2EyfOYvY8i+w01XjBjuZqg9zSdHpDOzAuejv1VuaMErtO
LQMkNTFQEbLO0HaLNBMJfVarK7aWwVMTNVYZiSnYU9lITeM2NULiAU6JsSuICViI
/Wbs6KKwGxMQdjw7LgIkiIoY6VOkQCwAMEEi9rrnh0R8iIxZicY3eOtV92hFwyus
JUFDAsLurMSljlSZzL/bDlMVBH4ouLxjbJg0QyRJRz2xEbraevrch6Fc9gZtGNdw
CwM1JJXv8uEDa83cw5Ni0R/RvX8ikjCJs0MvCpEKjJmrTscaf/7d6kK/0dXcoBRS
/2LZHKfPfHKFCExp87+CP69/+TGvGcF8LFN0HwhlCqSiJbbkecua1Sjx18RAj/sY
Z42qcsoW+dzX4F9s42VOcOSPIOE87wSxYHsPri5i9PC40nviHD6Dc8ZzrRc3VH9x
8flTlRFQcFWw/U4pcNQEIIIXJU4MQeE4rA+ph2B1Atm8QFM1ua3oe5akqSE7ykxe
IAvqhGWDAGhnDI8u04fYVL3SGUledJ/UEoYzkFqYHvKAw6vRXl/mzWBsTpxZBO+4
mwX6sKPyIbiz5biB2nAuL37QcbfRTdOLO4kn/7mg2EeZ4HeUBvRV7CCqSEm8aUHa
+Sf+8PIlWHu/N6zZF+aHgk/1GxOpwcNHmQUKtl4OnqGn2O+ert0QWYaOG7bzFA4b
Fk7+i0yXg1qYmyytoyjXB3WbKv2c+//zF8WRrGvar+PiNFrxN33htiGibz5O2tAN
UZxqhBJn5VE4mO6766fJqVtEqeopnUyjQHKdDzlIgoYzCE8YCtLYv17FcAKPA/zN
WAzynJXuQ7Hlohn60egSh3K+yqUlTBibJ2FLj5YNcauI7g6njCIywFoIHenuzuqf
Zyi/wcIe70FRMIsKmyVOwOUtdJJJVowb4yzQF6GSnjzFpg05sxAw5bVkULNqU1Aj
rXF01ns4EF0l/Gt0+v2M7aDRhy54LRlutHv7xvzkxIakFoedDYdjTZKLHZrj8JAK
/XfhV6+ErCeIi1sOBoLc1I2rsGs+/t9cv7248upJP5rW4z6/XzEkYcbIBIcBhd3+
KoERl/ASEX4fchpziWKNDxJZ1UFkR+DSE5u5O/K4CONMFWHOzqHSP46kto/JVfLA
fzOE2vJFrqC1/ajrZTV6AubvcfzoCkrQUg3pPsBp4J/zs/mFq9Y0j7cUdPUsnEz2
iI7J7vG8/4jTsWNXl4HDdw9f3NXJFW53dKZTDSED7hAFA877ur8EIYgg8uTDy8qM
oqfep8sJVKia2o86m/o1Byee3MZ1bJeaMvRSuUvFXWpdMEHE9wsvz8DRL/R++OE4
iGQhaTfRlve5d8cW2dfDBHBOl1VXRqPsaLHC376eNO3cr958kyqcd46XNMQ/S4iB
x+Gj0s3e5l3V4cCWbO9Mh9pppojDp4PmMqmAlO8R4mQmwmJ/gNvHmVK3WTBgqZDC
weB9ZJOpQr4blqCZgWI32aHZvfmcxVBxC6LzVpiqePwzBcnf6mlKvu+r6xWswqd8
JdcfRFufhzoPwpCAF3ZhAa8oTUu4A2V03TBcEJPETj8JuZjCGvLdCATO7eOu7jTA
WigeSLYXrawLj7zGZfyUpeRhPcreeLro4mLjO8sje/pg35giT3Pw/9fSplM4HYJw
kwmclacuPSedL2jBjpwEJD2M1TeRqBf6wtQmyGT32rm9sUNgKzxJDHG5p4+cQXqq
CLJRgsJOvOG35+2VOVz4L8nO8E7DXLZToXfbPLzFbKGn0R0ptQ7fc/VTtkcDsG2K
FfbjdfeKrM9XIxwq/EHXj6LLJKzTnZtqiP2zRcSO3oFP0FZHg/i0bsY+UHkHe3/T
mSNYaUEj0EiWuzkIP0ydi5hVuiHvEVzDMkYU4cNWW15cBBy8TWXX+h6V/snDry75
KQ9iFIjBu6Tq257ij+6+g9BygwHE972vliIZ/iGFRpLItUC2AnmP6gbuhOHIgC4R
a+sayvDs70SnTtNEhsnme5999l+FCX4kgdC/7ivTrLGqZ8++iDUgBgzg5iYvFVcw
Mw8HG2OpYcVESkqEbuTLB4/R4rFtj7KyhNCfnsYShrDFBwqXuJsvALQhRgMGoEZi
TO7cSYzmyZ1/I14rNxDXs7rgj3SZHOrVvU0cHwMdwG9EPuQ8SPNKhzmUyoTXX7dD
YBkXV5DwvMKYzYm3XRErgm1DQsPTDGaVejzP23Ky5CGTqlv6/ur3GL2QfaeK+Bne
ePh5zYa2uZLAn5krEzikUPLVxeuHSA/fjTG3pyK3Y8G4Y2tmelDO+0xTT3pTKHAH
Wkz1gA2/o4t53Tb75Hop/0yJaWrAJfubYa4VCyWfdZHUgYzInHoVJZhserRk7Bwh
RyXZzyuUWGhYCDsiyujxB6Cjtu5tWAXRAw7FtNyFZe21bLRNHcjr6u0EjCfGhO4d
KHS11M5qIfBkLSbnEYQK3BeNjhDeDc5q0tO0eMZQE6lmr8UsNfsdDmLG/vr3LvVh
U8cS/IWrK+B1C11bNjEEPTWFt1orZADV4ZDBJrt1S6OrF6PL9zxSsJ/TryZE7YZ4
WFj68vdzoVeQoquu2HNXMI158GHlV3PuMbXEKLwxvaFx1DglBQMeTiYhI4N8OChx
b4J5H+PE5MXWBibXlwG3xKQw/h5CJnw3PRuH5eqA7LSkoiiYOmzp+/qDU2gOcl/s
KwqwOyGy2lqfni1O4yKq9+S1Z9EROKIjbJfeuW8NNqRVbyi2Lgxi75cdccga9JjA
UVelKA7h6ar3VnENc9sJTSvqTovZCm5u8/+DKRVpE3EbChCPC6Rqf+E0/wJh5kF0
HapWr0J9O8PJ7+Sp08m2/9canNJSpeJTL2fPVcUm1qWMj7mrf+0OjuqD57kwddkd
yWh5xmYoSnLrhqHScoPGfxzvgsrsybQB0bqADlUSHOIhnmAURkk6inryVSx9i7UV
inb8t3H9cgcOVgTXNTJKmPZeU9UnSemXFDtFYjvGfB1TTICa0O33qCKQ5ChqFRfi
K9z6iU8AUyZlJCJBL10W9EQu9qvUcos+pJiEZRFkrzGGndaht/7bxaiJs4D695Ma
BAn+ChHtd3HHbi1Z6sFbdfjtHen2Eji5YNatMWXGJwQJmgp8U97YPyPvELw7QmbW
NjyDEXMoTjoUqxFcBZkhpJffsRZ+DOopWNZxJivJ2LnY7fpNnhx3tZOspCpSPuao
XeIH+WyJM9H/HI67JvX1vjeq94TPDy7H/OC6OBvfDkVy/dA6SpZdrwC1knbStBCd
PjAeBpR7+qnkPd2oFahlR6Er8SW65aU7cZ/4efSL1Wa0wG8H1VeQREAO2ogEvnGW
DHHQa9pTdm13XWBcaR1Cl6+7b8SUBoJP3MHTTesenpVJr/DxqtDPibrZwJ4AjxuK
Bh8P1s1sinwpq6662LMDfQuO3yjk2Nmrf9/1dkYV9EbSdg1OkmQh154YgQGdaT9G
sxYaMcsbyhc2nFzIaxJrUgP1htASebw2nSXd0rQWEeV91De0yezquuBr4hvgOWfF
z0GhS1OAhh8dDy0RM7QJGPYEe3Wu3YaGb4hddErOwkgctsTuNPEzWlkmCZXub8yV
rLP0At4GetU3ybTafNRSlS9KgbDLMJjpjteHStOzWoVyg9vd6+XQ28EH8wGViWc5
Sw+U9Py++vPOiDbNwZWTxRJiNX5xjGE3AjJCjkL8kgbxAY7TdvMOx0VZRk9IGG0x
cEWfgrmuHwQhAkMnkSwK+XvlEFHXXWEM6QdR+l2mBAosGOhJvbOLITfo1N2UO6h3
QNLiz0RlytX7ZXF4qCJgQDRES8timB9ji7EGC6umc0qtvNPmbNaHyboaxI1dbnZs
P6j3233GoDJssrGLM8n4Jz9SFasQ4+xdqXxek25Up8QVX4kLnpk5AUaBTQyfZi+q
jsKSQc/RBiiK9HbwPOTOO3BjJZLzXuH7l3gG/xdVO0Y40bRGWK7x6Rrqg3C49JDl
WdX25Em/Hw5pzF/j6qlwp6uLUiH5rcB/c4E9S/tqK8QLVc7yQmGt+23E0c3NbPMi
QrkTqMGvTMNpL/Aggst4lR1iF+J4K/HzA4xPdh1Rs6MmSCYjCqek4pHC3vXCPM6A
z4NuOP/UzMG9tDi+sfIsOHAqN9CLCzSDVqVyVB8lp1zuZigEzWSdUTGHZiuj1RPx
j/i+81PizVwNfbiuhMiMYzZpq24i9H0HyqKwib4MTQi+3a3RdKr+Xpu5EAeGcnXa
FswtwLo0RIm6unuEUTz4mltuIgedWeUSt5aIu2zkZX4jN1MvnmWvf95ZbQxW3AvZ
ql2d10X5hNCG1xSZcm2BzMkChE/2ndoZQksut1W/MbO90sA4kJ/63be1LnAviNJe
q/e7uOnIbDGRcQg8VgPUJ1aNgg5LZGbLOE6Cmni8Qa4re+ZBo1AJAfLQhzEEzNyk
o9O1NDjWlOwCMaBclpbgSu4/6Bd5Q2uD0wdrmHO8CJDKkydLaTQMRHs+d37nBI5B
CMx0alUYNbJFIkY/4Xd4rZs0jOCLchD83+OPC37eedMFCzeU+gOlVoL4lTUPgtEG
sf7FajhnaY/59r4SUnpXpWok2mGxn3wg3jFTKWrVe4liASW8IMmRsm8MiAh370gg
wjNkt6VtaWHEZMNAB6ZCdpLNN1h4pGvDS8p2EfnYOVBu/liOJr9uVAqpdsySwq67
KNl/cjaRGzNPeJZdwMyj2uEqMXY++NEVjkNi7ubsNK9swByB5kZylhXe/a+y96Zi
phsawVIK9J26OG6YLOaSW0sGJzBLRzZU1MExElngn7PIpm7XEqR0/qcbS8Y2uxWO
XGP5IomZW6sgMw/CJXRlg3r0P/cZF5bVWswvz6ER8O1lqgVCQbgBdJmCJNViCKx/
0+oMg+U57rliMq3EgsoL19I+W2tRotXUcT3b1Ws+U8T67blpJ43M79QEsJtMmOq3
mj33qvKnB2L5i0ThF/ZkrYHvuLY9Y8MSuoZGmfRYWaN35VKgG6Bp9ZyWAvVTjQU2
rGJDUjAqj8UUGHGG2hW9Psr+6Qy1pOtWGuEXoC+0fIGl+jmbDF9LmoqoI1hpfy7H
iJkdsx+A8ekU3C5FM5eUUUrRwyj8Axd3JTJJwXKs+gwCjlXjtkyNksJYElKPR34n
68mJk6GM3D87V+npLBSCNfXCJuZFQn8uceN+a9IILQXGZfmEku8+1wiezwEPVZaK
QtW12l4A+Uri9lvRGHlOdNjhqVWzBzMZDe9JVRIvC2Wk4J8CYEi1RdsOIZ0YE5SY
5rswiJpvQvlUyCTDdHNJiqfUqpHiKvikuSjZhEEUjJy8YoeT1aj1E41WId5rw/lk
jT1ROKbRzv2cM0KGcZNpmXkefSxela0cr3EDLrKFtXvy3q+UyYOtZkM1nsTW8Lqx
2EL/vWwI58pTlqzj21CMgZboLjsWIPysOZSpvCzpI+BfYZHGD6MZHmw/0BzoYzYV
BhjuMgn4/N/DIQ9R7WuPjSfNV0HdLIUJtkDzpcr1+URtxa1YNr09jI00oMVeirJC
Yn1mPv3ZXoA0tefuxCtLHtkteQ3xqo8obuNAf1/k39HNc6+q6jlpbTNmiFbliYQz
v/WKcohNWCUN9DMMcnVuWs5b1rDkrNChnlFHMkaITYel9i3b8iuIF4vOScwjBY6P
hDxayDQoKya1XKectfETjFcKcsLsY/w4FE91+YQQNuR+SzNUckCwfQMQFc7JNbLD
1vXzu7tUU1rRkkUVmNbUk+Fz922vXpzrumlKGwgdJkjkKqPc/WEYseVM4QlALYNl
NmV22xZ8UPJAdyNyTEP5DzyK25T6hK3uUy3tqyQTubM7Ql4dVuPwCXWKeeQn3fES
KUU7Uer66DeZ5WCmbDruQOp2lofrIhhmZdZ4h1GDhrQUIcdtuXN6qpRcVEQs+qcG
Vo/pmnlvkfWm1TVWasWiGc/97qMD1SkJ64MUlN4DVETLnQoeHhaiko0j1Kw63meE
alcbuvxmCbYGeWICH8mwjcpqa/y2pzw3P4Dak8LqfpHdBTW+B58YXhBqA18JRSIR
As0xfzdSEOP2gL9SZRd5UNwik1dQM0qy+onrbfX6feNdnsDRstv909MHH9Dq+9ab
2Ci2EY96oxngtBWG0PUl0dZRG7zh9Fp0ZzUT936olIAhQ8vbbXm1R6pQpmk9Pzzr
PKWIHTEKU02h7goeB6zy/wlhwXIgb2fJV6olT9nb+FtZW1ySyl4XcFljw0FoJeVs
VeOrfqKUFpefegC/LP0WW/saLEoJYHC8Ia8/Y8YBEfYgnbwBZFMYvC4ybJxP49iw
QC1DUdfMoqQYyeDg8SqmF0b4oqCWTUAllp2nGtPHxNTN0W+fAHSxfWf/HXMBbnHL
zOQSBIbdeeCUcTILxV3Y505W5Loq3PPxJeYqASoHuARUKWhD7OGrKANF46KqPFNd
PRi2YxC0aiCSZ8rHqTcP+RMXWOqe03bta5QqEm3F67ryVePY1My4c7y46joCLRaw
avTL96YB2Jel4XhLvK7OEhwOl2S+hj3IAgw3W4qNw0AlS+tPYYtcKEe2rqQIJhCH
MwvFt0PbH7ADAFM9l+d9vmMT0t5TlC+bW3aB1NjhcsLvVu65y9eByT8Rjny0Z9ZP
wJkCeyYGCAxYCHYK+zalzBFUq5a4I4Vrk0Q7cFLmBxuCvl1weuAFj56isfkN4Jzx
uGZepY6o6dRH0TJ+01DbpL6XU9AHLc4SnLxlsIeftw7PrI4F0ovOolMegzT6zkTJ
5SSXVXBFSurUn47Y4AXL3oulX82luMh8h+1oZXR4Fym0h2OvJ5XFlEFDa6CJAZdS
ZEonBTajhwePCCM5h2nHPCQQzytYiMGMOrPK7UFzrKAUhS4M7hTe1HWDugkVZ8xO
gaSQQ4d5ZeClmo1KhJzAk7jGyiG6XrDje9FgBt2XzG5CAC606Lem7La4/4UJlsIT
OLuBjvX+rPyAUspMQthL9Q6SS6KqHbImpx96ynquaociky7GOe1KY9yUeHUepFxC
1e19KMQk09/JCJEngLPqCKXNFSd4hLBF/lQVxukDR3ljh9YtLOTuyy4103+GAYXY
TXlh1dAs8eOIWvU6/mQh8VfL0qH5UZsp4wYfhgQL/Vn83SbpCdNUtQBJjmS17h30
obG0ge6C9y/AKWiU2KpmB5dPYzYp6Oq8wdmn0FeCJDLgnllx6e68d3RBzDavOZbV
qZO1Lauh4g2n7bR+tUAEg+9sRVxaz6zmXExRgv834QUE0mqLxmTHw+S+xw/a+ult
m/C/gfmQeBpl/iyBytrMlNnrPhpPmxOFK1fNucSFaPWaCufNJPo+ldXtrCQ4i9om
MiETeg7EnaSaoTSC8fgpSHVCYEr+qmIYDBhn5nFtoI2MtDjk+TPZAeQYT7IdJiUJ
bDcYtYk2n8CmCB3ZWeJTFMoYXbYJ4Chs67kKCwwmrjUoTYx0AedNI8+l8wS+MB1M
013sDZw5E2UeRfigBQ6Zo+ll785CjrxNiR84LBQV2vgcM7hEEoM98fusRqaBUy0n
3qDnWvCggwsoMzFK9qBflUpYCIRIdtnQ+TKDWakpM1XiG1DbG9n3i6+hcwlaMf0d
TKnIMELCD1manSP2eJUMBAUMpS1Inwj4K6z4d2DTFzHRNenVBEcCutf/c5PtvnDO
joFRHlBiRwyw+4BBBr+fdyWsnWcCbj59MYkO29esXlb521snxtRs3l+TNe/rHAHd
FHyNczXr1g3XhqNN7i2HXpFuaFEfSQS7Sbwr5GxLVqkbMKKv0SQnKAlupSeGGXDt
OM6gJgkitBLbgSyUr40wzHwXzTXfOt8CITj7oBG11WJTP9v8eadlcfiHKHqfsFG/
lsQz09VTwGO3CEnVy3MhlFwOzTh+5pXXYgrEwcqklCCNQmCFpRCcRmRfEXnf6O7y
/rupBcHS7YYVIlZCAoN4p4EvjZGFqh0EJetU+RaVslQ0TariYJHIpRi7m2jNKWvE
McUg4HY/IVFuxH66HV3hwDyuUa/Nl2FqG9CX/kOQIpc1n0pXh/hklplGtpkESxl2
HWPSMUczcFPZXhElhNe0sNf/6nlyaY9SlJhG/YI35P3LiFIk7e4xnryObNYT/FcQ
B+ApDbTnCiFUM04tWG+o0JoJ6X+ErZQofwKa22xIlvDEov2SL0gJtl8tPa27tOU5
YDAerwnY6Gli9ACchZ0WkVtvvEKwDgfN3REt0qlrRTtDcTxK5jynajth66w217Np
LeEKFw/9VrDygF8UO/Xa6FrqdrtOICyxHMpzQMDyy/0RWGxT7yBlZB99/bA/gbsf
ELG5cYObGGgirR08W4JTpce0jbagU3FmybwdVMPm0Aax4eI6FzZIrVR17SDp+oEA
xrObwFh9vT7V0OGg1LPuYu5DctMUOXF6EURv1ME6oEbZQ0Z+yDekxzKaTJKe71ld
tFINqI0BxeQwlWFfrSd4ufRG4jxumuVPkofDJY16nQp2a+mUEx3tqy4cIPldCLZJ
+H3lSHAgM0GVKrZ+1fy+KEDpXUfOvpiNoTOQLulVn12KHb9uEBr37z2v/56WpHsj
V5PpGREhPMClj6hHO3aoNCNCYEqQmN6GI6g8aTmemE2TTpBiqDgHtWtaEI+iPGXl
O0JHwhxOXw+DmIBhQuvG/YqBtsF4XoPdX8eCPUhaIJ2jv8bBL9guB8OAks5KJq+N
o3q77fYKmNl2c3t9soWE/tjdmchTEanjXMQM+YfmpnTjMdAauIHZBZLWrA/fZga2
i8aH/8/6YjdoE/2jJclAdSEtCtdqwaTctou+RiVlJ8OkqEpryJAij6RqUxCtJR2H
gp1n3tssL0ZwYd4guPHqk8TrwqDlc+yiDQcdoK/V08XP/ouablFwtdIqf/P7itdA
w6qqg+cFXym+EZTr+1Wz1Iszf6qxW87uULpHhNtidV4Yy2KEinpyrcXLJ4xy4/YV
qlvBMio49mM1H54W5VlKovcomsKHUTE9kZ3K3Ot5p0IJpRPscUZChRKXQg0IBLxy
6CKnQxemXzRevO5vZV1IsK/s1WUG7+YHXaqG05DLytQsYQuOZZ50zDWEvxSHi8Ar
w/zsNveN36qb9i6lnxy1Vo8GxDa8gyMp69liFdfwBBtdnhyt+89D1ae0T4Dlf2Gw
y/h69p+9GmWOZ2aRVgSXlj53EcHWkxipontgiRqvGpoa6A9BjsJm3eInWc/9JxPY
ZV1uqvjJM2Xh8iFODnV/PxHMorzAzd0F2PUq9SfNhjZvf4+QW7zADveRsMAcAHqx
46aheeohjy6FskY+winnnNXPkMrcBcrQkm/tkLJuCqYAqX/xcwNccJ43NawY7uWc
FbLVFiBeEKQz5v8XcuUfBmPAiQw1ron7Upptu8vl8K1q4iZEHPQ+z8wdqNfKoNCR
TnkazTgbHKhYoeNAuOWvuNv5OI7k2jBjztUG82S6mUqExpRy5lciMrwSlCs9oJNc
3Gc2R8bNnVcQVcaVlCcwVecm7mhiY1+3wr3j9XbyYJjqDuQ5tzf17WTHEA/iqm7U
QGFHVLbuCGaDS5LQ3qAzIrBI/pV4EUf5EFWfuWF0r1MRUin5FxkWtPw71NGauj4l
nEPlKRF8hu/a/Tyar7+4huluJlmYSGBeaLJYjnwIpxuTZuo7OPpNsVh+3/6WeI7O
6948SplO4SiWrlhuF5p68yfZxn5ytaU0av5x6r0P4+y/qgdJwB1OBUZZakq9MKZ3
G+gG81LhmDRadYG3AgSt2SER+ufBSZgTr+CiCQhV5SBYdozbSEdtpiHcSbF1meZ/
43/+5itQrsaOi2O8+O0Mv2lC0yUMFnUxAMRwU+voMOfuICLUpqnS5hgHmB/S5AHe
g4nod8HX/dmfOwerG3q4J9+mNMTWjGRYjaVCPg7Ebfoe9r2wFjH+hSNrnP9JMCS1
WCQOKtm0AX8Q/TAG3Qs97v9Bu3FCiRTOO1WxpLFvytRPoZ8yLxp917gbmw8baRUA
LyJsobkxvajjpPjL514IUeABbvB1WvvgTKr6AddqwsTBNRkiUQQh+idVIRUOSrpu
VoG/pP/4VSENZ2fWRpjw9i4dTkAQDG9YQquQFNhUyA3hbPV29FBEQS+vs0y9Vn6y
zFQfRwGJGbhCOqV5OhyuN60B9VpSRaZeKkhtnTgIkQP1on99XcU+6y5lT2V20Qhm
bU6YimKfg+M4RuGaKroKSGRaGFoPCU34lafJvBYdk7klqYEUCdS2nSUvZYgUBSP/
57f1/iEybjKa0AQHwT9ioQYC0cT7DowQzcBcINf8zDtOky9GYxedc1V793+x7yX6
AvNiVnd8Tvr4lW80RCmhTYNMPFxT1BSo6OidPcoNb5eJ7pfrbqTntYnALkpTPHbM
uxpvcrOHcR83GXlCHF86rSmvLkRVVMOC41NSzevB31cI7/PjIBzllhcBK3U1QZ5Z
IzIPoEgMb9ZZPo3gfDfaqGKU+a2/luN1SBrvnb16/Ssc2SNwuGt6Qtv7mO/ps57y
Nn73Pl0q8v9LapzvFOJnmqJS7NyxSaeGktH2OjzC7DeRVKN6JBxscKbIE5ojJIj/
lRB1TElUibq/n1xJQPKsuErBbGWeSFtfy6Fw8lAjjpIqtmt/LM6WmLBvRfj56F0d
CJSikDA311ZOOHUbHetzCABGo3CMc9vmacDmf9X2euPewRnPrToAvRfMyF3bKcOE
qpQGQrCHFDBioOUCN5x60XuUueAzrNoV0cmADchNuMa5U/Y6rZQ73lCQhGF3zOdd
HmB2907DQhpoBgGZ5HUz55JBHT+rn8SRebuczp8kqqr6/CAyO9Qxy14R5SvJIOti
u5C/pzLGtRMLXvaXpJcHxBPKPE5nmQygSV3lcacmmpYUfBL27/Lkh4ZlTZFDxp0b
7AbCUCmCHXX1G3a0xsGd6x3yBeH8DUYu5UAgmpqSokIHM258T+Jh8HLTUbnOHf+I
tLT1slUMm16kjHWNMjsGhlEZOH1rRedvMDowfHMOxwxnkXCKjQgcWpmXTBPgAIWp
9+yqrk4ScV0/8O+a59S5o4x9fXQMKwWrH0yM4806xzKxYPjFgG/B4PWlGRT8fUHk
x+J/3R9U+Xn6WyLNiqgdAhrkUdh9+u7TofqPs0lPxeHg0e7nWQvamldPUQeN0GkU
51ZEWM+e+ofF6HFrGsETb2yh6ruYqiYAlI3RfgxgQ98vOcijMqbSFSi0sDONWM4p
xFmiq0zcbcfLJ6NP4r8xpqV9P6hV18kVigrOUeCBK4SixLsFgYMOK94TUmHtcnGX
CjGmgYem49gkygUurJcNBLW+4pmM0c9fIz/PEuccvDNiGgAsepHH1rSAg5fZWU1T
GBx+2IOTj+wDoSIire6Y+LeKb2uAAaQ3J8BB2sTsvnw8NyguThk31k0m8X+eG6ar
VH5+tZO+xWbNF/qglLYmZue/pDpbgVn7V01P54iro6e/32nxpJXWMPsxfrRyvoWg
xaCjLwLKnOHOvQwszJoDLun8/Y64+t2645yN9eG8un3+RvGXu8EdlT1g+gLISzGV
ptpTFzPsLbjG6sUcdp0+rAejmtYcALRvRXozVVQGOyqzUvW7+Zm6h077MHjLnbAL
zsoXq12UDfa4i2qUiQAdYcwbTCFQ9SP4vXjBI1i9Cx7WTgo6vlyfzc8cxp8XlUl2
aNpX83/ggJxnfbCCfhLCNRpZ38QXdlrkYVO6PcIojiUkbYUP9lM2q99TLmxFCq6m
kuwkHzHAY6TWmKFir6LltS97IgzESbQ0cc1KccWHAxrVZY5JoTWQIswJEQx6m5ZW
5LXWzGwqr4MixjabstQ++1T94H6GJ8M1ikz+E/9V5CvKXcYjucgJU6TTRAWYxdd/
R6LS+N7ty8pxHfZaxqYJcEDLwi5oohfcgQMWLB6a2Rwh7z2xe6sDmt4wjJRPWHlO
J2gWPBjXIRmC7zz3QGhgjZpwCq3OC4+csD16chdOevKBjs4/Sswmy6IAnrl1JIGx
kKMGzjUshbW1Eve1LOygjOxUYdOZa2vCBiN6RXQzJTySufclcWAH+vybR5u7skzC
aJG/dvg2emOIDLumaVUEwC9VCEGkNLGu2lffFDAEUGMULEl3OsTZrh+rj6SiI+7x
R9FBB6N77dJhYZwXWTzz8f+OrN5HObIi0bAqEiGrx739Mizi9qb28d85y8VGB897
0KZL7bMoDoCn9pIPzWkWcvDYblBtCUYa3Xza4yWLoHneK5K9qavo7mtxbsy7ZDTz
imwDRt73zBL/sZBjbo0tjEvJLLMrCWJ1U/1295bBz2NZmarM3jKEo+ASHTxgTtUf
Xg1l3KSqYvG2g20FjIXuw7/I2/UaPcqYQW/zpTpHAqGjzfTRZ0wdHAyjfWv7Sscv
WViNDftkCbgdc/RJAm3+bWNUoquywICeCpUGVBKAjtW1WWrobkPyCUlcrwfcLXnD
PmuxH+aY7sPG8XQxwvofUiH9g6K9e72iXd6MSMK82fQVvxSvlKbsTu0cSr9FuHW0
eVQytFf9Ou0+nKawjHW/R8UgndKIcCSrurDFx84ZMtBiqT5hjIwv1smEeq1Lxszl
GkxBG2q3mCPhl5AzcyBQOezywHKm3oEit4H01r5YzE0bUcDqwZyWLgEigHLLb1kh
abcHdUPlEHnH4kmhqSGgfXkhj3tzhxy2KYvOu0lC1ztDOBKglW3zN2fK1cIrsowz
f6hCyVymY/yolaATF708ofdX6ZJLY0KOUbAMkx2v4yPS2B7ggT49HEEtg5TUZhR7
XWN+FfAMnbr/hlUlT9uGDNJzOLBtIYeyDnXiH3iuqeCEivpQNC1Tl0mvzLh64IcF
S/Aikrm9YAHA2CBxluPUFBdeglnhp+EifOvq2HzOets9SjP/4F5NmsBqZRSeCa20
APmuhj7vk2uo5JqD7Cp/q+rhLJrzm0R2FDt1B/7gzuqCIqqNeIo4ls8Lyk3WYtfA
1DyHwart/GGKjxu6DxtitQ13+pycd2ik3czwu1XBnqDq76uel3s87/xEmxWX9nWV
tuPTrnAINF+oMFuNyQLjPFbT+qQwiScfi9OnOz6CqWamprpydpYtupv1o1+ea2Ta
/1eOHyo+4bccfF/cgboyuPY+J5jvOSEqqC7aHPO63EIyKPdIKAegkEiDfrXzku1h
K+93GuBhmmw8xv586bfYLpgH9gVxVM98DWOEAT4a390Diiudl/sMT3bKgIIsCvvG
dlrI0kwcfP8FY/QODxSJxzpkIxwpR+3iR27GFlpHedBAOgJXgu6IFrtWLXnsQX2Q
BtiUw0yJaVfbKPY3+CDUyHjRHIaHUqya0WNGyBOj2g0c6FzqCTn0WxQ/XMIeWFO3
b/jGJbQdRjKE7QClFM4Ku6flMH+b2H9d98iDRClJ4nvBygxm77qIp/GdN6CiWrwQ
nCl/oiotOCuSCEogXp2OGnRzrgznYUjLCFdxZEWc4glGYXWxDTfbg+pu/xosc4wU
tUhJYZO2I2dV5LCRGeOTW0FYvYB4Qovl5ZLNTpqirlWuC6vhRB2/NAIssnyEnzUc
gxwJ/Eb1aQLkbWdgHY3UiRZ0TJVYpkNlCge6EgKoIimlMFMOTM+6BppnEecZGoQj
zkj1UgeGUBufjiHl7+f6A8fsthlGbQ7otm8QF594SsuUXGYpW5ezkLisl4q2esLQ
trDfhEs9YRNAX/2mi/hMEWJYmpsSawFfNjSeRtF9STz/88z39hZaYkEzLc8JDugx
5ubpP1MdIbN6x+AKwB/tX1KguXWuDrNyRqu4TPQYqD69/bbTRd182elgZzptwBIu
XY0Jny4crbX1+TDdMpgZPJYD0XndmDMfOxA6zvaczAn1NBrMoOTRxjKfWxSIPodT
eQoPWgm94yR7RXJygWlauw62Ws9EF8IpvfMyIyqdqH+hn//BgQN/sSxbzqelIumZ
Ks5KvRRxprijhevQEIrsBlUeZNgklqcZ8gkJaTNSjPbtp+BjqyA4wcXAdFsYLkWH
U+t4mdSlYLyiqiw445TWlSRdJ/TOokMgFoyivwFj5iYIXDV32apEIrVZv2SVnHQ9
CSFFtir8ATY//ja+EbM6eADyqskhvcZ2FT1g3iwySv+PP8YrA6hODKMT+MTNJ7/H
VhcEW3YjraqQBBZpwx4rfMIW6jvXChbGnt7Rg48018qQVDuZuk+DJEzi2OV5ZXnJ
vc6MTP8LSYO+scPQGKRfDT8K9FDLoLVHWi/pwHxMo5JWaPC1r3i3O7dscULRa2++
tYayub6wnmlHjCcu2raELAzlMglVcoH9msUKNc+XSYX56wem5gQJTh6g660cTq+s
Cu+LQGiR+GtSHLWSpnt9gbUTozKdzUjzDhQZTEcrtkOtGrVGiv821BN47UiNO+rM
tND/VWxVaLt3jSLZJY6HbHztfKATTLF2nhcCySOWA6wQMqtb/1O9zip6T2yNz9Rc
qNtCiWJPD7881F3nMJ3Q09gKSeDb27HseopzrlEF/IaCRJSJo0XnkSsT1D5eoVM+
mcHQyakw7Jv8eX91DjpNJ4eygBxREsEU5NfYBnkxfYmDfZdSETyPXmN4Jmvc0Zt1
ITSLbdPtB6YND/ajd3v/37RPDDyj7qQ5NVCJZmniYbbhuB3K7vg+r7zmorY2M42I
z7F6PauWaHz7AFIDpdlX6VT58PSpqxbcKLP9GSVZKC4HSOszvL0HmNbc2OTinCvG
I5NtpTdWBB1AR01VQOHg2OAhVRK7hTEdZj3VruMuJkfJOZPUvh5hYI88cfVtDkab
HbcTSvjYUHZXu9QZg6WxMmkGD/YLqBZCA608RbdlCwFyJUJrPRzY5mLdE8pHjCvE
j51Y9PJV9o+UZogING7W4MWiG4l0ouc/gJ+QZootuoMcv2WGc3kbCLdIjy57Py7z
T81w9OVgDcYG8Ry2C3LVP+En6dxXpr5TNqHR7Dqgw1SCbIIBbDOyT0lBUMhtgw9l
p4NU+f5WhmtagRQxWtd1yvn2wh3vKC6iesK8olMX9LVqD0lRtA6gXjmX524HlOAq
OArkN9FZAHua8V2IVbDPLrntAgoGt4f57RACJ3wxB/BFKF3kmqRK7XfxBQ8tH2NJ
J/MLN6OIXUriH4PUMwCZ8UaCWhGTkpEIZRhkiMDTDd5iSFU+3ES3d4fBXv/GB/nP
+yw4tjOTftyKYHhVMZ3WsMUIRiTWllNTpi8mFG8dfLSAvAKuqHJaHZarQdGmN7Xg
fOkNfxTKJhLuAlyBTwy0WP+3v2WZm8QjrBhRkLYIg+/sIlVrJMMEWdOp+WdeBi8H
n0Y9+OumHpOGcSQIbTSLkl7MAouNLseLd5ZK3p3ZzbB3QhVdA/FEr5cutAw/PG7I
dzHViQdRVwWauUYyekCWE3B3cyEUPYLcIudvVB4HiRChdRHx/CohvgLD/0dpT8ld
Sq8yaKvOH6m9tDrIAGJ9kAnBH24cKGc2HnEi8hoFI6noN8effCJSfFU+Qrg/DoGn
pc2ct3hKd3itxJurMLcLSwxMsmnuJ4cKo9qdjN2c0k+EpXPtE5o1huNs91YQdm7Z
iIx8op6U+zueIKFMtg/dBIk5Q9u9lowvmfKvafhFRiUXel6rN4eEcJFhlcxI4s1F
t+aa0BUNsGtcqpbJ4v6/6qCMEQsHyNHLucC9t9MWV2fTEu3NYCr2tTvJz+XQPBZD
AiL4n+sjN8SwV6CeEjg/8TSMe4cUpkTCUhh4R/JWh3ZMqzsUX2HAS9sv9w57x80a
mGnDOXDCtnE8G5T4/9o6TjFkyA20n6kjFg69rDf6k/Xc8kP2q8p88B64d5/n/BhE
MKa/7AKYEMOm36x/6cwhMms/mlJJ96haNFBhp7tVrR8uDRLuBtMw/xQQkkCu3L7L
RjEBDlIF/2pvoIdgDrk+lr+8VncAmJNHMEYcSClKHPtHQzomqecaAMbQuWFubuyB
9gIm6Y++VnnVC5vyY/L9AQ8sesaS1m5+QMqcmcCdU01fiuINuaI+GXBWng2mOHUE
y1HIIKsRzhDStdUg3bepksnj5ccgYBvX3WUUz+5aHLKCHvMQGseh0Ubf6WSCGpZp
Zkgi2RLcZm9yRSDL8Y5aIslYhJY74f8x/5K2A3UOg4L8yWPnLIdgg5Q+L+P+W7id
v6FprM80kvgPZzJb6eRMRMs9poaiWNvuMLEb58KpoPC+9o9XPIBsLKom1f0HqUG/
AByjrb/bkdxQc4APq8aRwtvKGwygk+GPU5WC0exXDRzd+VRT93TGzUp5Up+wjGyb
A/9qYgGQ5KJiciCgJn4M34QHqPP4X+7jtnqR0Iu+XoTy1MStjvK7y6H4a+mGDR73
sIE72dflafirrRQWlkZvrxUiUPBLYQ61KytbXtvnzNkvgtLw9OpGjQlHy1AzEkiK
rhK2Xkvj2RLEk2yBFrqE7yMu9zXFMY31zzZGS4XCNbGhd4J7bvVBhafn21XEtUDX
mJAYToPWl3B4dB3zOIb2ZrZ57WVUaGFpnPlPrvA78334HBvenpUCk0PAneA3kUfv
9r87laI9EcHsf+MzT8rKtA+xcGm2KprAQspJFZ/R3hwU4j9Gyr5b7/7uF+/J2gB9
hy/6kaDWKi+mcbhoo0xIiyahvGaClHHrtnIWpEcingx2/7H9ngEeLUaTOJ7xd+rR
dF04C9FdbnhWEORqpny4ZH6k0hJKXoK9ipQc1U+nQhTBigBd/wIrx5q2RlcEOC5Z
wjfYT9LkeSHvKFhhjguFkc2R5yC+dxtLPPd1H9bBKQJusVJ4VZ1qY9i4ir3/mpv4
yHBiuvqX67y5wa4R3H9CSibgHX5b3vEpoHG1x67CGHn8cAGMrGIn4vbKBXUWv0RC
Kgtgy151lrpo6+qB5Gs/mdGj5nwoWRLe0rfRQqAr/qNqs5E9jq4R2NeD1OtxSf6V
rE8xEq4OFIASOnWtpu0l8ME01hUcMPCFv35FR84Mp8GvNo6dmG2DKuraTL8ErpMj
jZoDELNkGC1IvTHLQDeyKcTAZdUfscYdHDqyJ7zuvU0vp3dBNikWXi/Bms7A1Yr7
1OcRak54VK6Iapi2zeGyFMBMOi2YxIdA1MA7/fMqzEP+m0SEJ79Tbj4RY9Qztpiz
Y0Dmb3w+iYkGfUto7KGy9Zcs5jC639DsH23dw9g5l9NMPgBB7iPs6syN+EVOshiu
rzkIpdRz3XshyR9UQs8ILT7BSzB4640bRx93OU2styLbSKTagpfGdduhHd0Ij3GL
Gptm+wSx5RPGrrn9AtIG63atsg5cgkZrAfpkvYA9xpEt+jWUqhNgXc1IN6vDAc9j
gIJnW4wqKMOWzj0WCUu0czQ1pLKONYK/4dTB723jEt8hXZW0xO/yU57lT9SZ2S5m
S+/81MXC8Xtu+QiCCsR6LAKE4mtvEUJczBAmvQg7nDGp8YGX5zh5wxJThyzF917+
kc56qI+ivyxsNAKg6Xbj1gOGvYACtQ77zH9zfcb2Jy9OJ036Xfk/CG7jVPn6bTVI
DobJ1Gj+9b3khr7L0IlQtBlt9F1YX/RPc2L5230XdRsIn0cySg9pti3yeE8/ECZB
JsBrYWyeFtQjyD7sugPyP14XDM3BQZi7GPw+fpaLiKNJAYhip3GK+hzxVJUoXoE5
ayzihVqUAhWw8B8OEgVwWz2rd+dmf/cgHxVnF0kJYfEV7uZFlyGgC1R/i/Neo6Hc
QogdQV0csTu8mM8CD1l0QE2Z+LZK5eTvlwDNZLCQB2B5fDAorJWVPE5GqoPJeFhY
pxCAOLEJbI/cNBr2S1rs3wWw94rkfVLa6cKDvtl8snIL16Dx8G0C7Y6zazZddTUs
ExaU3xv1Yt2STu5b9HBqMVOG/1NjLNudy1uKI3QAqOn1Bp6EumepCylyaPGjz8cy
lD9Bwoo3OolJp0zo4ElsBXfRFa0SEwuhCLHLYy4MgcKpSF527dgX5tWp2JX8Y9MT
2l0ueVckjijIV9yP+QHUQx++RIPR6btzOhHezaHSpmjF+zYSAK6xOYM+ZjzH1BJe
QI5Xi9XNQxf3v7jYCkooJWI3Ky6jsKv0Um7DPGMi4OLPUN9FgKSCoxmp6CjxVXaN
M+MX3UgUYNfjgknkYjwFBr7M7aqmUsuRXFANwz+s2OwGPvZnirg85YjirM9RdSh0
REqBdXCE/3BHLr0INZgAa/LJQQeJUiymg4XnpE0BxJ9ZTzYmfpZcVHoqkEcsSt14
i4MHRCNGycegy8tIL3Fkuk8DkIe04HNPzHgV9uSn3KRtH8tgjGMxYlLZbD81ptuR
DYeXULj8Jffwt58CUPelc0TL+fGBcZlIlFb+6ti7nk/Zrk3VyJpuqNJ2+xd45+V2
xlvSqWhpSs1TedMNtMkk7ziZNBTfLJ4j0QWBHTSb/hxMpx9kVzefGDR8XZxt8hqs
/p6L1q9fHqWt0iboQ43OqeUly9XgsgvO8HId3kmhqqZjsTsxlLKZnxZbSZq/Fx3S
YGyw5IKIWSb3d+LGBLieneSQEVP/wVLw8BmySAFl3bs0Xz3QcZ24ui98FkQ4nsHe
g7wVkb2h7fL+dCRjVTdX64jZfVaOWkZx3Wn/5sG/nr399A6dYV8otoOm8C+ny+3U
0BkKTDpTwCxDd16x1YkKpIuoDWNoZJrepNvIXMRHdIfenZOaBEq9vulfdSPP9TGE
Vhq4PweITSeIUDwJZhEgSotj+V5DWrr6qRDT9nBFLoarb5uwr6MFjZQbRgmI/CLv
cmixEiNmejvScecfMy6JTC4S78x8UKcAoOQJJHLPyVYZYuHblWq3J6VpIzfQqAy6
HcHB7vZ2p5RDG2CWeV/3G06Q8vA9DEUm9+MZTc6a9CdmRmZoljiZBn8sCFBeZjEt
9bSnMVkpaPQ+NivsFSTd4jkyGh3mWAYtY8MIWdTSvJGxE953/jXaJjhW6BeCeRW7
RCl7NLNfodKv64jljew+bO/EjTpJb/MdHawkPxCOuoQIWSc64onHthyIyGTRi+2l
Cz3LamJeg61IiO1RvDTPKL3CtD/saP13awUrJnRW6dLMiNF+w8nPmkaVNI5h867A
oqH+o1PzVzN7CmgA8U7X+yvAD4MlWlsWf22wM8wPVLUaYQvPQ9FlYTXEA3fvqBz2
PWNUzsm0wjl32OpdlXUrLkwXOwzkFcJO48jdzQ9sNnnZynjI4Fy7fIWkxD7x+6ca
1v7bv3pNJGixkOo+KWotCgpTajUFRnUYUXceQ2ycQ4kCKNshpIIH9Hpk84HiaO8f
JqezY7T1ou0FKdcL1YvWYGUIcrf6xQiTM5gV2k57fME1ofSCJH6cvuIOUtkqVVqD
xA/Cnu1XqvkHgOYExrf/ba+YFXU9mByVOEJv9kJ9AyysQHEdThmM9Lflwespji5P
jGEg8kkHktMXGN+rwvYuPJiORVP5UhTLighvcuT3fmbgGIzMJ7Q1zYcPVIBKmIFs
+d4n/gQMSVBUuVuWDwmgbLejZFWztDYc8nIl3i6f24XLQXh2yuHmAI3NivMCmv37
K0xNpEM7HsTQT6ZT7VIGdw29QvInNURVLHz0jYWpvQgpm7qr1DWuST/uPsItWJdT
DNKbcRsr11dJf26Q2ebYfFQZs+lBEX9vOsXrXiKfO3I/C+Xty2dCGH7nsHGFoy9q
KkiKrLvFpeOIw3Dx/7D+TmPQnEMszF1bCB0V9Xr6jUszl874M3YjJkB/yqklekwA
k7IdyFcWgBVlOZyHokc4LcQYGDn6seuOzHRxf/EuFICXlXI+Ao8jWQt067nY9YOz
rlfz4eozf9bkxDzMWu3MG22pN73lqwRk9RcX8bSAv6IApm4Cc0PkrSGGRqYPCD8Z
RXyiE7meENXjOLimaLbL1d00iKA5satc2CdU34cFwzvFvB1/wxXpD7JkfnS11+5W
AOOQKBxaktvgoFrJqHLhxiHb+VcefDTIiUhyjtorNXqgDztiaHYGpE66yLGDZ5di
Avu8DZ9PmEEUoy3K8lVFIMYZ0LbKrBESnp5HEFSAesIegwgOb2n53KjCP6JhvVBl
7mjHsrGI2h7eaUtCpatL7sWlrXmCNt4LtPw25ecgjQiDx2b6tgsgUzE4ZohrOUQ0
DDOpm/lHcyRGNVP5lEv3Q1qjBhXfFBmKlzTixwAAqk9noa9G5J6hm3/3pCZsRC1x
GN5Tj9G/DwY4FHrFghByCYJWNnPg2gHE3w3T2biLiCdU3zt7JM2y8Igew9gr0gW7
ctGBVA/T52kuh9nQVHm1dVZAHf5dKAEo7vRgYjX/7jyP0OaeMm6GnsarST2yJOmE
n6pr09mCu6F07O+sHVlOsFm4ohe9gPGCKQyNBxxOEwTisvF3X0ehAx9KfeiqRZml
OcUte+ailAnN6xDxkKGsIzCVHJDTVMuhHOh571DtaCXnGMDhmSlUhKsCApycBFBx
Mw2CM+EnixvZhGa9693KvDsK9WadEeq9f3wWE1IzDsFPAojENtkfO4SN23J7VHEn
DShZNWmLIVYA+VlLlMSkIA8uckAZe2vorf+94kaUZkTOcOwfZS5LFkOIWMaJjSHS
TkU8l4GN8upMYc7n0zkcr+o/iQnktYLLrWAoQhd+lj5fRzjSvArGUziBvNgjJ8/0
hJrx6XTr8O/eN6Apef1pHjdLOKErIm/IN/o3m8wLnzulWbJkwtvpjDaf9cwUTkuI
lL5iFkSUyC93PalSd2OWtJViD4Cw2ALQ7ZIyMByXRH3/tYyonAvnDEnA+YFHY33/
O97m2adAAqZKPD/dLrZmAR3bJ8VUwZJCWvcjDI3YjeP/7ydEttGz0SG1BIRI20dj
mTvZpt/FDfSAGMbyworsHC/U17qqN72z4sYNPCYPVy/10dIxWp1I0lffJBzOfxyG
vjx8kmFr3C7ePGpFtNJFiCe2dqCHe7UNRO/cQMj2bE6SND38PW3MHvq+jSll16So
EUM7d1rN0xSWpvif7xM64T9SX9imZ2aadg8ngHDJU9xZpxhkF2rNpVBaD/CED/m5
i190aRxSeTRvZDISyvEXvYIytMYqKW+CIBHpMnaCcDRcsglJIhzkm0CD4Ac/elTA
po7vNC8Jd4pJ/1xwJ99K+9sF92hRJRX8lXUiILRFW6cS++g8DpF2yj/fzsrABAzQ
DkBSXWTDJ0RYgJeT/3yAAXLFd3RPraI2QF+GFzR6Re2SLQcRbY6N4naqH1TsYK3k
d80M5xDmFp2CDDc2CeZExa5A9RW9U6l9Z/9RxU97cF7A0z6weHRdGuLFm165kaQZ
d58/gw4WR/Sl2KaTZ+2dHXwSOy/yt8dBd+fco1L2w7jSFXcYphUxxoZXtDkDaVX1
QZG/YrGoMsYWtCsDV/gAurhKeANkmzoToyR5RF6sopY+bT02ld8S/SVNUXAL8y18
HFDRJgw3hLrvTzC609qCTBAs64I1BW55Va0xLzoHMWEM5LZfOvFblNkf71gxqooq
GhXjK02Cgwc3sehtGGD8ogOr1mFZczLRJY5fLNKKV+P180MdF5hp9UIibz+rGPR/
i+U/5C5SUv/yWFnxgIFvdAO+bJHpwWQW8RBUBDpExN8kw5X6eTCqGJgljuQyN2xY
+/zYorWecfblSeQieWAsXu+VYUCvCfKWU4ecAI8cNjChgyx+c/TevdmMZ1Wr2pMW
wWZMkDUZnUEviYVHstGA8liihwSqY0+fRhRIEnKoFswaBT6IrD1i/lhukHneGWff
P4L9HV4jqOrC9I72TBuOrX3jvTAdaYSdexaCb/dv9N9/cfAXdSf/3BxetURCrCeO
1HbC2rwvTThijkQQO4sLFMKvduf3tPisPOQJbKsoZ5CxkUKs9bmVwhwC2cHDHOXU
C2sqIUSUqozXmyiwntvuUMjYxFu5Uu6u4waHMEfrqO6byp/oKJV0Rjq2Ks7BCL8+
UHf2HNeIine2YHkK/RiY8bLOu5Nzf5MLOvcJA3T7wYC9rQx+3B1765C8OkC/O+k0
vlVmgpRyM8aedijhbY4OLkKHkrldc5JdGKY3qdzCHa+2rqY6xr7rjUl8yqu+lg3E
6nBx1SiPxBUFJ3xwiiSk2fNYoklQtDlyKZSbhd2A74RXIdEpRmsRIKPIF4+r3L8V
HKPQ3RRHPx1hYtpU8HYoffKsm+dTK2bx2dw9/E1Ht64zZ/aRgia8a7d0z8wlIlyP
kiSi2JptBaWdkgGTE8btz9+P0A1C26OXYu40iLOXWP5UdJfXWpuswU0shAJCWI6g
hxDS0sqv75JQ/7PB58l7KU5tMLaeTk/36JsVJSQMzKnImWBDKbwmEZd+WnhW3Yry
8QI3ZiGTFyffybJBFb4wV7lHAPpq+ke9aTbv9BODyIHXyxMaEFoPFKeT3YgUsa4N
WVaGS1GJF94DY39nCV6aBJXzx1i0CoZ+9xLTLpSSm4dAblg4WiRD7JEnUbwT+ogV
nBnqnNs9dFMqhpR3J0uz6TurnDR7jVWIyEKSHvP11VB9fzRh2YUn57ZZzi/rZNll
i+EWIxsu7QzF3FiOQvXycpSAXLE+q+T/kfSQ66tW+xeClbxiIQ7RxyzPsPp7puku
Z+NvyJ2EVjW0iUU7sRPyH9Bbw85Fs0ljHDub5RoukPYA7QDTgEX48zyDLkoqVPkv
sV1QSXgn0EwilSIQmDfcXYD4uQm4yHlGE4LGin1HbNBmjnyoyd4RvhRoA7snihsF
fmKjD1/d3HJS8a6ySvFzsFS/drckOU5HhpdwWXfLlrLBnS4ukr6SdyM7mcmWkKqr
sDZCaaqu01n4TNQij4hPavzW8lVHqb6bGFJdjTHUxKP38CgtmxxXFUrEx2PGKVha
8xcA1X3iKP6O/ZEZvWVBep2YRbv3EN5pGIubpijpk6z6ZsEfDvPuOUwMXaeX9ATu
wnPuaoUSL+XKdapSggGxJ9cbkkEDNyggWpjmltebEiYwgXyz+tYPw7Gf4XHDwvtD
R1q7MfTfP3bKbX7y7JrYh6t07mX3b2PgwL4CAf6N6h9YcbtX16uswEOdJkx3bXiD
8mTQDcMevzXwD5treMBa4JWfLT4tCs+oSk/5I7CfkXV8sKUh1LIpkWXhGYTl9KHU
13f7dPsNNtJEgxH2WoRre6l40U2z3uLkCP/OiP+UBy1quCFCVbl4mwSHOygyTyhh
6Cvi5VdJs0lfPxl8QkawYmnFLdYoFN1m/am4RX7Y+CTdJlcm2+lTR1bcPki+A5nj
JQcpZ2Pmp7U6S4O9Q223Q5IUopnHy3LUqGblUNZynF4E5UgoxQmcdauxCrR/vqdP
oKhp7kDP2DwV3cfO43GAr65NxKHp9NZUfOZ4SMk9uRNCic9XRXFO/QN+1MmfVfyM
NhsifOdvuQdRyLRtgl/oPgx3T+lENlzY/HIfvWWwfAuJeuwcIwfBQV2siNlMiz2t
ca8jeJAQbw/hj5Ahm342SsafPiCpWZNYeaD0VYe9yKW0TuF7Nj4Wlr4fCTaJD3jX
NIN1U/Mt6hUTiNuNq5rVSipRShka9OtLVV6AExFgS/bZawcQkhNyqUju1N1B5uuY
D9wdM3aeEXUmv2sj5eWOWNhBFzUbsw+4DbnDBmy5GodxLxBnFFMqiVc1zyBlhAIA
egS07SraiIHGTVVrisTTmDgml89wTrjIV3DoHoZ7S/ztJEKN67oo1IX2rXILcb4E
CQgmRhwDOz38UNfA7HtZN085WoQzYc+rCkFMpZxPSDDCjeuo6Re5VWK/s/ftn9pw
OK0fEeUS2DQftFyXy2TdCFjZUkc56i1+H0JRBdx9poU9xI7PNeu/SXtOssUPV5yD
vCBjHzOJA45gqlrnVmutHeGye3C9dEOb94zpI4b2JgyttP2DkOVGnlseYQJ9dNhV
iePMyqWtqEGoXbO4iwRF7SiLjhLLtDVWxhRMx9tHXCun9ZRzOBluqUG8qRXcW11F
4nujKATnKAl1xo+SI2KoYgSIJimBzSuj68XqNr+U0yavfWIVG9YdHbDqhdDodvY2
+iRthCIELqj02je8QBUT4pQFJzbzdGWTwj6zdAb4l3HPV7PrpOmyvl6aSSL4rd+a
QQRlVC6O9DrKxDvEqlzJ0b3z62GJYnzd1V78SI31rA+MECbNjmnc1vS1k30eruL7
l2UrBI6MB7NcjirOykn0V3nBv4Q5bXCdFtbracDiPlh2HNbrz8MlzVNsuL64TK4z
XPG/gtGLmXcMaIxvT85CT6P60Jjo9MYX6A5x2f7A3qnNPJA3O9h5wYvmrGxlJHB3
yK/2WOo6TDF6I4ce3f5wbOZUkGk+ScO1z4ZJq7OOknS3oz6y1lDuLr71ixuzELlw
5uJkf0Q93vXGKcW95dTin/NqxekPhmYgPtx5DsK3mRX9zJ1G1FG8KpqEaUHCaKSc
E1lPsumcUSJ3VQBPp326TYW5wWXlyPayUt7Ie+M6DcwRijRm6cRrt9YoafaaMMsP
ww1xvTEn8/Kf16AX/v7KIVA11JC6lxGbAVsZXoZuED0FjUC0G4baoYytzkLpirKf
IDjVRX8rGfyjpaGALuTKZ/yk4w092FI0XUk4N8O+TgqsnRFetQfHIPRGEeY+c3UP
2Ou4EmbKEDpL3SgTbGKqr8bf8JnUv4jY0lKgcDKPCGP3GZReQDF8lHCrHRNAHN44
XB3EYFPphk6ydzg1YoYVUkQnU0SCzT2VjXIhZ4Ole2VzOpphkzhn3mYEPR1qCRF3
iX5/Aa/oqrZZYsGuQ44lPFo+4JOVTa5+TJCOPH52I+gKQQ1A/S/yGuZBrizukVen
M8k2iltY4klLYPmfJPTqzrHqQrlggDC8cUXBSVDJctxjx7dvnjQ1yuS4oDiTWsg/
uFM93DOcuRiSOKSQkh+3WSfEw2DiLhvFf4DgAHP4moF5aTgXFoRHw/y645KpGbtP
cWYfagUxnhslklZ0XsDYS5cGHlsmKynsxHBqgcelkK+K8F02nEgNLrE8f8PVjeiD
DOTb1n7EtlSw/EzeW0py0E/7BpiJ2S6BaNUu0BJa9KYVotZ+4dz51C6cwmTVW8bA
puQR5mJbaQ5gmHDxYzbk1Ysq0au7ZqJwmYccNqZ7Rv/7Xxf7Svm8w9jIAygzb/sm
hidL4pUJ591Fv8JCHut00ubpfHjJ1XFAegl6AX/lc6l/yd2qZnNCcdcLEbmBvCKw
iTXKkjfYSWq+n0Azdc4Z3j3GOr5pWgVvD4zYJH1UOFxk3xUzfTO+/OwDIBwluvFw
7CHK/2ImuRiKHMzecrYz5JB2EVDNMe0ifEoKxGkWPEAEg2miD8KN1aFQv09Wu/H5
qw1MHbyaEvfpW8H5VGxZJEDmlrN1+4dC5eMw83MgxO/xujcpUFCIqEHrYp6eV4ET
F0NVQvw/Sfz0yaXGlrRdXxGfqcCnmRgM83wH4iad5wTegQGMk+IpI0Qc21Aguwr1
k3LitKkxrrkTvjIqPTATvLzld94BjC+XdzkF/gg3vGEma+cnytxwfpKoBNwCKIWl
HnI27X+iFiYDZWNVodxpo2S3b73W135znjjlqtRKOCGCWGqjyfJgaWFV8ArOOiza
F3iKn7Wxqd4KhaZBLZvbgtmkzs+OTHP8apW9ODuYwrrjAljre03bRkAdcOz7uIn8
hSlaCWsbDuCDNR0TrWAqLd+iBh1iLmEQ9FJaKgc8w3TFtiVpX2hyDHbgfI4AG16K
Nzr0vvO3O5vj3WJP8r/LxXcpLTbGRvOOIFtDQoqpp6dwLhJwazNPN+zNnxHZZu3w
yxbe2xDhfaygYZjlRJvVmWZIw64sOV6VMy07aMPxB604OwA+SZxqOnH2eIU7twfZ
l8OziuwLnJIsJ7yGtaZE2aB+UogsOcDDiAbZvXIWr1Y9JZbaU/VfyavjRV3jF7Bi
AvX8cOD2dwP1AzyW7QWc/VLtbr5D4px8uTiBski1vxWUF5iCGzC7B6VqOO0PTGai
1MSyAzHo3kAHYruzgBR2DMshldZZlcKmpxbcVqhr9E/qjMfVmbX6LWSjhoDfGHyK
tLiyBP+k0KAMN5T0vzeduZSfD/i25C707SAkjDQXYRsXJKG6X50KwtK2Vp8aWy6i
QMxxJ/0sCUCy9AF+pvYRRynwQ3kSHtNYkQzaRv5pvc5XBa7M2eNrS49+2905CQIq
ISsTZYuYnSScEklC4mwK3MadsNkYAppXi+7fcJP1KfwiQM46u2tQkPufYlNgadKA
yayCYSefg6lSsGshNPZWS3SiefPJJHiKC0OCr9VdU4NjnBNfX5UYHT3QnYS9u1s2
6+QtEfRiQiGYqFlrERirTjYuYPu2UvbOWMd9UELcBSk1X6MtBewTs9nRGSF5yCMO
g3ps/7Km2fG7vB+n2UUr1A+nPNV8OsZYd+wHMROpAb369DLTOQZvPLqsHwGBHICh
A3iUpuQ1qCI1NisS5VXoJz/Tbug0323CE6DOJzQhmHYV0IR6Osbz1UQhPsDRz5LI
6pzRwRd9DhsswKOMVzoj/Ey9a+MdXcA9HrMkL9yUdWNmhaI6eNCC4jjGpU1dDNPQ
InJUlmmXrBwIKfFPlD3yWQR+33trgEZOKImgAlgV+KwX5UR1tLsdGRDZG7/agl/8
K8GmvQ8M6l5cvySW/HAb1EegtYeCxJw8UUJcyaKMI60Mgk0Macr0Fl0PK1pf21H0
ySdiSmrIV6BmdZNKrTntf8gCuIgYtUft/6yZdV2UQNZtoTM0Wx4BgKzd8gB3Sgc4
4WP9Pkzd0bVob2EoKsmVoYH8o6+l0rtSbszURs7qzrD+tkKcBnc7XmYJREQfyyzL
66/hnAkKUP9KqWMVFl3s01+7oiH+Z764Y7yWQJOl6ShKIndxev5QuSZefRDG8TFy
6eD2GIx++Ral1itlKNut1mz97o4DnVtVH0XGLQVlCDsIrs9Jhp+J4vro/5ke98U/
DATqClBFO30cMN7iQoE7krDfg51MxjPkJDt1hPSpbvOCPDAYHaDMO1VyogjM9kbS
Q3TlNwQz1i+KUSx3GsjqY+V6Aj8CYRD00+jBCrr4MUEhRp3ifKyDM811rhYrjtoQ
3qY8DI71+o5bj/HX/Fbo3whY+XlTeHX1kaoPzra1/QL6gnzfS9PmJBfHAUfpymmy
Z7K5FzPdt8sgd17oJbIClfUHiCO3tSrVreiyHY2vqr9SP9I2qvuhQ5cWHlG5X55a
Nh64T/g3oed0CMYhrUevGZhrjv2TKVXxiw6qfO5xH/rSJYf9KzubWc35zZROcab3
A+DMMgumNZkwcNJ7QmmjAJaztrR5gTaDZ3fRaoEaQ+rmBkWngbkfh6mRKQaPKBa8
Tt5OClZT7amLkkBvtvWkq6gE+bqU+FHd4pbhEblO6Gfzgi2WY5g7hMwutPmBoGVl
xWbbnKLfWFooTVki97GQNOJwJf6Nm2jW7l2Tcl0Mvml9/NUzpq2Pa4gqtwOI2xnL
SjIGNlEzSUMGU9vAN5uxTHUHeq7YSBtxeQk6RnVTAke5hYQVPde3Xm5RSRZDkIfK
n0p1RakDUmhlKWbGKuqyWH1SPWMVRIbGjmaasmGMJ4MwVSw7B1eBpl/IKsvGAj0V
W7QTp7+fJGejJDyfo2Tjvyjtpv24wmC7Ug+V304dQJeevFMUJvtkdEwBp3tSbdDm
uDKizGGmYlbnZLcNKbiD0FPjsXmSnMTrurIClUJ1THGncixiRwi6Gsw3pevNb3Ab
0+K1e2FxFF7oKAAYRmtA0jjHNuG5kuCfOiCUdb1SK/muY68hyX09cbdAyXaio7Vq
7fLUzcYqi0U/r2bRxo138O2uJukA6YwOgqHhryQR/hcM5ExqyhZYnLU90yb9rMfG
dBHKvftjl/eaFM3JNPlg6eByLkPi2IrZTXHvGFr9XOwpjZVOaLI2vBIfCqOu1vwK
qRYVWciTb9VE0meyfr0KUWkw+LY8EieIxkZ/Fb3ytTCR/6CVxHy3kAyl7SB2mnM9
v25tcSvAnEy6hON/qlbhWoX08DKmcc5e6Fz3IcNtR/oGvPSY8srgxWxfT4upBh9I
TMVkntnen+C+IZp7fdNUGZkawV52BE4wD31S8+cPHm5jHQVcckcjVQAzY/Pmz7DY
1/ttkT2VwXr4zX9PUceryIfEX4iy1Ccjed+aYkZt1PlkaLXUWNziIAQpVdNLbZUl
XsNmhdrD/bQyUgwfbXJwrlO1kV8mJcEknpDElrW5wdNOhBgLI6qXBEJLbeUE1PFH
tYLDo2nPx6kqB/uqDnMymQ9jSV4OANavcVh86Ij6NDgJpB/9GPj2c6Iq/PK6ZJYN
bFTOevvy775EtZgoBIG/jPXk1vRucWoaeCP3GBxnJNUyOUzntj7K9Ne3P9LHmlhd
jTHHzouMZ5h79C+wLJ1Wf86wuun+uOAYVlK1qxP2kn3YgKdwA6h5sj7+1+/mBkV6
hGJgEppWmX1ijOWzKRSiVg/E0Ikal3Ghlfu7p3XJRg4ZNp+olIfYyrpB7uMl+PB0
oWYpPAlDsKYP9ilohsSCqUiCtcyAHH5qTLc7YN0d2ylEmF0T/A3Ypv/fr0J/iTg7
0bW8U20DVAdMZNIvELkVAdd6u+aocOrOhpefcSjQ8ds8Fr2O61sLTOvYh2yb49Rb
UpMkNAki9wGqcCWyalrTqDWEoPpa4XieL8IrBP4HsDunzVHjaL44vEUWmp1i7GBS
poxRGmezz1iVJzOH3Rsl807rTOihSdCwS42sJicio0Wt3XWxlinMePGepKRhG5Lg
XPFEIKa+0/jdgAAZkneUeOO86XUUuP7+4KTj33vQEFDpXak1PN9OFjO/rvIYxOCP
ok9P+z9JyvEqH6pKfbEuE/REGdpp0ymoORJD1nJG8WN0+H+FfCbj9DT2CPNoJISB
KTUEbSSFSWAAwza3OSuug5X0ysT4dkaly5DRWtUd3MkZRHC+AZ1ScS1UCf0kt3zT
KBk6bdnz/U7WA8CbGxNVQQNj+zvIqZ6cviswyxoxhD/bKDH4TthO7ywfX1/Lk/Pa
aNbbFazmYQU1e+qRTvlg2/PrtQql3YF1EXDVV16nFcoIvDgPb5p4f+pRi/pjFBZW
9WxMNK8fMv+NEUgDgTyEXleF4AShy9YW5i1TJid6r6O9VM0D8M7CIMZiPfETSvlA
q1jX0eHahNVvzDR30bkEouiEql24//QuonYpt8iWihMftilHE61rqoBVyS2RTccx
lLIQaIk0cgXlYVIjNYRpO5fCKWKlB+bnAoDeJcm8Tuu7WbYEkpToasJQC6llRvN8
Zt9yV1578gdjebSLcc/dyyTpMupkx4sxOmoJZOWPh407xl0zJXQwlBbe4BZBdRzD
R56UthGYOw8Ijc7e2lm5J5Do/pIDCVVuBquxFByKTIbe8RnRc9pIhgcSpbizH6N/
7YaYSySTkSV9BI2HcmM3irrjORChJmKgr/sfOhsWb01IeM0Ae+AFNoqu6S6iiypA
IoG7Uwo7rpjquQKPR5MgjWeZT3Vdu771xU0Aq/7/WMOHHa9xFdXRJwUTrPfBf44x
8MYlh1KcOeBXvdMY/qVKDLCYFU9X4V2zPdiaZuzzhU5MqJbYWGHZqA9pJuz34ZUJ
4+Tsm05HzBngKe/EssaV6M/WDDWXjaMkp5Me3uqvzwubwwv83GHEpuGpY9uxJTeV
s9LsJHmxuNhVN680dcnSj2pEorzIXTV/uaX/6Nqzv0E0I09+1DPzvobUgERjjyjN
XiWIBlnnBPOGnaJwruUi/dhlfCECb05zu01K336YI0UMQAF0CBPYSmW1TlGUM5T1
zPm2EFmWQl0lzMF5sOCoOaIY9imVVxKWS2nuAa9ytlV7oc4jsMkS5xBUdWgQ4NuV
+BIO9bVeO5AZir51Pnoj72486VM8M/SQ2f/oJ1Z36lzlw4qVHzJZ5UU0ZeIe1Gpp
Aut6/tY3f42NWfleewtDpPtOvAWXkTAauHtP6nRmMANXVL/ONHGqFSmfRYzRqn21
s9cltH7Kl6lAx6ztOc3ZyLS+bAX+5poqEIkDFYZF1AJEl0EdJw5VKc01lXXZkEQ9
RDV0lFjt3aUSAUTpUc8UHQJ81xlEQlvrp3ZmKH21B6JcmW2brIUuJRQEK9/9ekqK
0xOKeVbK9XgDXuxb8vMPRHmBo4qx5TuQBz/C3dkgsOZUy8n+j6dkfHK7z8cOz+e6
MQrAEOX/XCZb1x5JSdKhv+0OdsiymAKCIV3Dc19VoO6Ik5iM3WcnFSi5x1DQdwos
BfuvXqoWGMPDGwBUXlUoNgkjQVF0JquyTGcr9azYjtk1XStgHg/i6+WMiflZlzI6
ZaTOFmeiMSt0le/3bhTi2W43HPC08wOZ8zuV/tiOBwNbdmiEILJFkflC82gvhrJ9
s2DH4sxsUq6j0XoxUtikpiKKu0wxqpvxrFnSDamNBcwLXAcxMTczYxsGUbOYYBS7
HklnNGZ6v4afV0JBBeUW2e7qGQFPt88D+zZJ9rYFqWglw1KnUOEpQ60vzxI+BDse
84fcbvc/LmU55Xrvct4h+nHJPsvkW8XUnyWJH28KjLiNpB8DmOveTC14nZokzleB
FYAn0uk2p/GRv77kQuxePf68Jq3kpDFiIgEY3sKxfSZ1YdK2YeMt9/B4o1oKJaah
8pJEgJlZ9nt6css+6wrQc4Vss31FL6bH82et3VDrhI8JoS2Ozy3TC212Hg1NHgk1
6+UwOf+YiqTVVG2Qn6PcV5LAzGKaqcCA5OM7eIbVNAGm/krs0KrikO8tLoyQS9NS
U26IO9wafYrisnEQwlrih7Un62hZO5fyqQieTaBM9fvcXjGQtamcCu1H3D9LQrgN
32D7/+xZTVw9dpvpSgxGM1W0Tt7rYZ/FINVpzTgFiiRJoykpwenZW0vRfpoJeqxm
yMiBgj8lcmimPaLyw51HsbKYAJydyoeKl0obfSa1YXbdThzlWQ2wz7gC+VrCQoIZ
LSgzfzxPR2gTay2sSt4+JOHpn5WuYy2rPmjT9EsSUoqUmTkePiDmcUxecJEPEtWf
B1IjScvV18g+biv1yw4kw9ri1NBiDMYkiVbpPzXo3CyfO0A8HH2lHI0jfh52fx5K
Da0ZCnD3TZjT28eXHmUoN8QFoWIuJTWKKdAfnXE1eHgOfQseXwFkBSsKpnDAsHI1
7m+svyA0MoGDAVcHnWKdpiZDwJm8JQjNSncJt4nXzxg6vxY00ek2sOm+ukZIDnBC
G+CTlnTNcabGQao4dD7aN0WCYbTCqgjML8yLnTsyO7IuG4YYkgfmf/i5Zn92BGnY
lwZd4gGT3FzERAfX/MESgyZTwTskHwz0V0lP178U/6AHrOLuzYZoGjdeo8n+zkdk
qDG8HVLpUnrE67ViykVdJanEjCaQM5VfxP+4wDn73/8iiTSgPB+laGdxCysWez4z
J/mr8eCZ5wobY2t9qeyk0Ihi4Nnyj+ObHTH2MjOwEYFqYpRrWePLgdhedTY33Xzd
gZ3M8pdX7yNB131srzyMBW5fHWrSnM+kFqsE3jE1u7BVuXVKJaltIhI5pPXrGN85
vdMccF6doBkDTxOwcUFcbB+2gDHum6JesgZEDZUwG/BH52sDRi0JBvwyIGDg0hZu
5VuoFrIgfHPW5Ybv7BtidxNGbJoZuY0NPCFCORQU2nER5GNi2FvrbyF7T0iAcwXh
RsB5c64csiveC9H72rQxnbFIF/xJ35CVK2KdxrAXWjtzJneoui6wUJuFMIP1l/GU
qvDJOzHVtZDecLUdgiFh/ipRGs3V6fMc4wARWNJ9ChzZ4SRq0gFHKlZ+4HFh13Pv
12KZxXMwjwmkXggll0nHZQf7EDAeHW/nOnjUxYrYBV7li7J1kHckmAOVhoTEzx7t
ikY9U5Vb3pXGyS1jVtTgO5YbUf1M/0B/2w2NQTvFpn6VpAkQ3xMoT61smKBQ6Dt4
5cI95RZtdFGNVCfzQhr8mhZrdeuplHfyhFSoik4xN7tFh5EqQu9Y8bZuy0DFMecg
0u913OuS/b6kJjjbmaDHrmEuXZNUvLrG1KgAfM1CJGTaor6Q6/oFJrUlvYQvViNb
Wx4WLaRmTkYF3yxrb2tkSgZ7wX2ir4bEvuODivkjIDMb7JVHjimpJsRjIvgD4sBr
eEU+GxGwoFsWhIIHs18vqaL7eGSu6mQhuNni21EbY+zefgsKgGzmrne+WaR5YW2E
PuISrn4T+uyJTJ9cfQFdO02WryPGsIhiNVYCiAGjo9DAW5iEAX/UA2FfwtENcdAZ
MbE80DJhQd+ZZEVWUsMhuVfJbAVksWj1cOPrRbfkuqI8Knbh4ml58wrIlWo9VdQ+
YpGSDEpZutS+dzkkCM4cVRPTl+Yt/zEZjXXFOqUqADzf9QVZ6k+VQdFdYZJc68Vr
C0MRKWxtt8wUCE5TSlx5fuD6+PQ1oY4PjJ0pxJ6gP+Dz3q7345I1QQjA8lc4Hg1S
cU+JH+fhtg6Tj3IAOo7kO22ZdQhYJz9EmYy9OWNHok6IrCPulcZSA16YS1RIHxsY
5V/Omlfkbq13XxAwJ/W3KQ+E3CAMX6f3ip6deibGdl9rkAxGMj+ihz/o/PelIobl
DWW4zI4BGB6f7ZxMiIjESDRGnV3q9urkxzAIIdhPY9BL3j7nzNsT3YuN6mDowzC+
9Gx4SbALPXwkID5Lw9j3zt4gaEyZpvNkksKKi4k6A7354SUIrAAvU8iMnSDaFfi6
oM+WCF3O9zWKFaJNWPAcO5TVoPavhY4NLnuq7kFSYvZ1BoEb9G4qX9N2ZS6NQNHE
DZMzLJtnQ2mkXcLMxCxcdWYqBN8izUQobChNU1GP9YxZwhIaLxQ9x6BjW0LLDHsX
YfMN5z5Um1li1+aKObQAznQYxuMSAMxgZNyMoxpIATXELisCGuwdWa8CzaGuSYzA
PWYPAPBzrNOrKYxSCnYHyw2bJlmYH/TUE6G+UDJVQfoGutSx6YuwwpmeccY2M2jD
lRwhhBsf1vSc9L54JeOP2o9Qo5HyImg9Vvs34aUl7rat9xwRoNTN7vi2wWY5L5Jr
JLy1DSSlO7vQh66gTjgxCd8sEsxLa9hf+t7+bM7m81P6RbqlkIGzp4ivW7HfpSoU
xrmOEz1ev2eTGs52I2UScNUjfuqhgNG2FgUJ/Ldwl3F72EwCFirpkyw9pF3Qz2rA
y7+Xp9pVF8Pm1dvpi7sCIeLpc8QjupCirI670UVV0ulLE/17jZ5wp0bFFW804IsD
2Q73WRD54bvrQgrsrkX41xygrg6xUIg4KRN+tzzvEwkEajasGdZ4t2/0mxiH7Npw
DYK8pXDE12chQfJyadluIGmb5qK9SWOrDWSxdM7gtJTBXSmR9G2fatziXUMgr2P5
DrpKF14v/Ee3zF+PhbzoJmxqlm5Ophi3hj47sH9Je/YnU9bnfwrPpXVfhfazot7p
FXDewGyKSceL78DBpcduqZf6IoiuqqzFnhod6dltvzizN/jZjtKiF72E3LYL4q2J
Dgl9PYKWOYtK9iZHOL1Aky57dmKW1ZIKxidFMDd9kA2+z1ZxHMfL6j2k16TDXx3W
mqXIfb8MrlOW2aeLVb7swE8oDdQCFZOK0s3FXaG/83M15Q8a9hDu9M46PYNVi1Xx
JLzvuT2WcK1vwCZwEuH9pfInRCsV9zefPaJuEhtzMg5yzPT/5MjuD49zcCxPpHKL
tWzY6VfqBr9cp60wY6tltSwFrkoN89dcr29l0eICF8qvq0ZIsBlsy1HnaUsyE5ZI
7PZQZsshnIPdQkF41ENOyqpzhy82sOvNvEf4eec4GC2Nghw9sLv0n8p5zN9qdJ+f
SYThuFrvPRKpULhcMNGD4Ej7uDwVwC8IzzkTy+HLhjbuI6JaQDRZ4JtXDYnfW1QZ
J5howh2dQv10kKa3ZDRIQhFaaT38FEKCAklM3JY6D2AD/eUDnDwoipGP6OACCiaq
kZsPUAYQwgxv8/J9fENRnvUQNEVeG3/3K5w+LhnV/4tRl8SkV/R0twKCnzQcLMfn
QMxdrMkq4BMOPpy8bSJ+lkoSViyY9C0DB0EVEXE0PQMAU4zj/epCmrNuTs8VetUF
QWyDbF8fRETGVQaHApSN6+cvAJIQ+FxyOgSiVBaJEIP4qplTrQzVPJy/FjuIn5pZ
NjDiKRjHHA7kvyNeTec8nqqEO2+dIitcVjEiXhJ+7b5/khNmewEvWJJqUg357ylb
uzIIFF3Sp4fiKb1yFtiKeuVlQgQEpmlHuDfNcG0Mhvqoqq1wHBYTtC365JG3NMPM
dDn1Ucc8O+ehwIUTdjWEGA2684HGOjBr2N9NS9QnuglP/9nVvdbRiWCW0YASx/YG
osACPrLYPHheqh9daLCRKf9FczlBFL1TfVa5vBkH8/6SXTpuIA2DN80rNfice+SU
FsocwGthdBiQyHWc2PJzF7ptJsUXHlymnalhHXMqtrWY47DDrNc9WbarnZn3Iid4
SiCURmc/F8dW7DtZqP/elKNINRiKpqprtyhTz1YTT6G4YNsJujKuzqH24q0SfcZl
M4O5GRq774YTybsDPQUAerZvG6jxfy/7oG49kFFijq90wgXfTiArdt+JC/OFUQxS
+PwyhVjazlxx783Jr2PTjtvgcNnlaVw+Fk6eaSH6kp5M1jJzPt46pmZQEPVrF1fs
4OkrlSfd0Jxfmjwz0se98KzFjQbCxGUiT89qDkOdAdOpWSXJvWOoH1Phdma8Xp/w
zSd14P9gq80uErBExnYvnsOCj6hNLtt2xERyDA0j4zjrqDUcN9OaPrSlb8PdlEO5
HtDP9Eytqr5B2k/OoAEpl3LBB2Eb//b5CdGkQxFjTGjNeXKejF7DrfIZOZkJceox
8F16EZJzIAl6XetpfwY++54mPFhWFEKE/FQIJKviewkKpdLsi/EIZCjG6UB/P3Wc
l64mxlhk7DsJl3YiIPFrTYQeL8/CfmTWg+dE2z8nsNVePbOyVeeJ9W7qLAcsvPVK
fWPIAmzdu9Ojm7F9wrGAjP4DNF7hy2ocgjiuPNhaOxwEuGN3WMWHM94DgxlN54eT
Gm9bKPaLwrcTKTE0uYB3yd3xQPpikhbyduVZ3+yg71GHiVU9Xt5de+tCDyWvT+72
MnEGbKFcdXbrIkO+olyPVNM/wTN+cXPKWYFq1wQmnXZC1OVMHAjy098z0weLfkv/
FERbiIt+ZmWj3h8TvU3/JIFYocMDjYg/asFxt/D/kb+K8zrqpqznJc/iN83lUq+d
7g4tTKYsFU0N/pmwlJwChoGp1Ux4gF4t2Klkm48Ug2mEsjoAwCTD3v/ElO5sz/pK
A4tkpxqMxTjHB2iRGxGk+CIL9uXji+tCf2CaoRAUPAXBFWtYgk1Y2xI3gqZFb1vk
6FpZH2MKrcpAblviZyRIyG3bmCWUih/EWy+GF0UOaPYg+1EAZfdbWM5NGyPpXwgQ
noUWoBBzQU9G73zLh3/SsPLT4l9EouwIC7BKfhsek2SvoNX0+8m71Dms4s8gKTgz
ALPdoXV7nCRKUbXDfKH5qBQOEVH6MMiy8pc2fpqQrpbq1OIAuS7SXMB5HApzCdzz
GKedVQx8ZYfup2SZ0Dug9JkWkvoEstP/W5fEDQzQgKy41SA1JwPjsUX5DKRQw8B5
od2OOXy4Ma3TwBDeNrQCcERbFkuRhVT8B71hZhV7l4NyVeOhOYqxcxw0kA5NlK4m
2ue761klYLwZt+I5oW2aUB+je0OomrxjEk2lBu79y19ED8LUx/sUfbxUvcj/NvwE
tFat9UHIYLFnB2CxCWCqfIHm8XxC8HR7RY11ObmDcSBn5QIJ+uGVSp/ZQ1k7HS+V
OypelSRLjZ3rygUE+Km/CGNAkBBSwVp4funQENeWsiOwKxnsqESLzatgPp06h3wV
3K3GeQni/AiVa0Byqc/QBz81wEJwWZNUd+EYLl/M5YihPz9npMPsyeMm77FvVzHN
ue0Zf41M9Z4KZ/YS/DVyaIjFNTlIdkeOExwDJpBpR8+OhX1W+zYp4GnzmEDorKdc
QuCRIuapJ0Z6x7HvC7tunf6XvdD8EdV5SJFGpmO3bqIR4x5oVIwmO4syhwiEtg0E
H3CLi/2J/EPx70bRsRm7ELkXYeTV6fcV0V8iujOU0Z6FOoZ7Sml/wKpM69KFK+ur
qNFxASBzS4++2WsamGjMmSI5vZO4soyCQc0Ft/gSJxqz2uXMquE6iGFmRC3rQmtn
63xBsSpP3wbyR9CVZYDLXRN2bPQL1GhBm9VTdxckJ9ikuWRuKspX34K5bnqDajMN
fEwpDc4Qnv3XunSDn3A/KUkTSxrcqBEve2ayhU7C+lxzzb+g1JlhRdAKXPVjT+SY
m3SVIji5I8rn8n8ZRscgtKI/OX1ztiGT8Y/wUT1PgmWXua0R+T6EbdYZHKCiwApY
BeLPXbP9FLINVCM9ztmlxK3vhkONuij9H/pVZG4VOrI5CcljBHu1WO4yAf0irqT4
XLtViqZB43SMLvmwf5KfSmWG13XWW7AvCtg0IX6ivLkgTTqMY7lXoGYt1j6fJUJI
hcI8IMVW1qOOB2kArRCypvuvtJxug136211zK4K5BMyaozwfIO57sMYLs/XlbBsM
fk3pfr1ffpX4bTe05ILswH1lpWJosE2tpFLMeRaI116UAQCs5pQIPWZG9ClITpfV
hDHazHpXSryITftnvfJiUplWUqc8Giis77o0U2Yl9zAtSlyjDmVkx+F21OMuaWtv
pqUqis9YR09ujTqw1T1HnstSTCsFGNDPA3trNForsn5lUox5cluiFRgf7RY7Vehl
slSSwwnayR6+4DJI3kaGhqFyX9zOt2AC6skxPq+9egVXP7x4dvq5botSQCJuFkTG
Q/EoqPFnV71e0IKyqyw/ye01W7IK1S7Cg1+Ru9fBcTwJ2Od3sY+H/3iXazoknJi5
m6yGmAEGriSLMxkWBZWNFV7UwPGc79ybs0IkcwgthK5dFefUJLAQGQVMVFPJHviZ
J4x9Heuv1YY1XGPGVBvWwGN84verLXb5tqps2wsKupSS7I+SXLmr/+ceBbGkrCkY
V/LJwd6MNHTtjRjihL6PWKHIXmWw5DHwlOQN55tHXWCoHwj0KyYt+WCtMVu1LI4R
qQ8J5GWVqS1p4dChHbvHPPSEED+Oc/4mkxL+3AS0Ifc4gZsMcUkZ2UfrGZGwC52E
X5IJJ/s0vSNLijOtQzzwSU1AW+WZFu06VmhqGbnnoCpNc3oY/0/AVtYIut0riDRm
H2o1RKmr2BF5CgLzaY7ssANM6Bn4UQg+ijSmcuySHp4xh5I0wlsKh4mbWcToMrjq
YSN9E3xV+Z4f4Hz3IakdHFuRwA1gpxN74yOKG8mVhQQ67Kx+xY94soDwjr3e1hDi
AuSFMkgH3sgnHXhrs9F+a32sM9t+itaDk5fzE5DqgUxMc//HgjVsGjrM7/HxqZxf
QvwpwzSxhIwytkE54mon9SDboj/POOLIf+KMlC/zo+Yz2T+wyYX/cNwLZ5TCn18N
gY20Xb8qqZtSeVZAWZaM6v5aVdATs1OGLM904tUkIqBf/N92LbdGTneaN7tq3oh1
GPb1IBNhFru+d32d7mDG283+JKDltisxxR4Tc62KSGjlwZxsIY0VXehGKHvApy6y
R8fU6bWvA7beg5iHo9WP4mgIscVoW/X1xtUgucAmIXOvn0tlhd0gIEEjCS7frXze
j7YaXSvHgx5JQ20POlqVXhkuCw+v7vyBCk80erB8GE8CikjKQ/A0Jk+K2hrAxlfx
foUesoItQixM7f7cNKQKZ6ZLcDO4UJwIx08AUrvWYlZ7kxvAlaNdexOd0P1YJu0x
icHJkYCMdbSCPDOT8eVv8aBMeNcLddmF8+w72SZ7wW0GBtyQDfh5Mj7zWRkdAflK
FAO2IsWx90ZlHndIgZ6HXfQkjCj3ve5Sc58CVSrPD29RFY6cKq1XDliF1mCTbVuA
GB1+0AkH5p+l/6aloCRUdHhHKsz3GfFd4apwUqFBJ3T54fsF8YU5hawBZVNsPoZt
2DfvKzPtOWqCPcn5dGkLeJMoRxgIj2nhQLjZk5J6afoFFBMyUK3xCQh8syKODTFj
5GDR16jHHYqtSThnUx0dn0+rpR5eUcTFxDE2zMTxAIB1KMiPM07M5fYH3nNZIJoG
I3mfS5/CiMYYHw/HmONPkOmXa51e9baSpGfgmOLg/Vbf5IkAGCqMKsdifQd1lQPA
IdT1u6KCQaGbyoHnTxWsC0XdTkBc2MmBit7ZfxCkGpszvMlsem4BOBU+zA/k7ZNn
BqSUgqTIz0NpH3jIXQSTuUcjd4/VOzSYoWcwEyk92ixN49I2u/wW5zFTEpc9m7aG
q1eeh9u/W4tkYIJPuTrk9AopPxCWAnPHoSY3/bzwASIaSu1SMtx6zaBfuoXs4gq0
EZzD7q0HR6jyT3CwZv7ij0P1jFYncIX6SMgjFwtWVfo52h6INw66qLE1GKw6oWf1
cXBPSkb8hgmqxeP1wMx32qXRp9Yq+OwV+ty7ThdYZQ7jri0xA3vymRjwGY6m9/dz
GU2FqrpNns0mfiPzN69ow3+7/5jb56+v3+Bhk300YskhCT92XnzYFjbdmwv9Ywl7
bQyD2hXDG6POH3OnezLYAFctAzBxliveoTiy0kNga3T06AxMAMX/xApfk7LJFuj5
5UIQK53eQSlpJ7M2mqN2IgzKoyZFIlv40BSIk+qIETyhX7NSn0mef33PxznyHXqG
yhyd1sY9/sU+vlk2m8O7N13hGCIfczjutkPtpTJoFepGYfyWyeCg6HbGmuYJHszW
CVrL2fVVwlZvvNT5Ow8VpyR4aUNCJ3wA8tsCQ2RAUdhObP2e7RpDzDMPr9GwzmBv
94X3GTPWqusCrZg1uTbx3xx1tbze7ztOXwOa1uQmFknibRCCwldFMkBuiIoRLu3w
OSM+WHotjmVdrN/kYpeMVd0LwqssYeWlE8Gwu5wWFKWXqXoaEgMH78nUU+ip8a2N
ybW/4c/k5eWdkXIc0hpA2Y1RVEZNMZkdZW5nIoE99+FJmVhpwWhHgGGzT0jG8G76
A7MNK7Ygr+FUAjcNAx3PJUSUa28E7VQaxl5ITB8oaJEMb9B1d6FQPIvSneiE74cU
zcbFRtZ+4ECMfk7+4SwcJPoJ4ZHv3JAui0v0ceogfAINGr7A1XWXEXc0JBXqAJgE
bEfaxflViu3C3LAUpoW7xrEj3tcFItzsUYaMZ+RBBCSRATb+nt9HareYP7/M5fsX
VNJ8jkIBZvvKat+ruH/hoPPA1Ue7I+dTN0i4JuTrSSPMGfmsAmz0sWyl0kzrjKcE
VfLaEmZCFjknRz0ketk7Cxo9kFaqDbRKKcTN6a75ejHiMZDDDgKw3rGymsiObWiO
748Cxv6SorQ6QsKjM5dip2K0yCH2yI+CIYzuJzSobxelWPcAkFpbavCPXQ6TED7d
jmUWr1iWWAG1e//H41kkaFrFjozjvDhW2g6F3YrwXYBjwb5abxx29CJO38/BpN9P
FFTAPmEBzebJKZVf/V24wGQvQAxGxbdTqxvGbigaLjjSrkl4VFRSB+hysB0ekwyl
/x8W89+zmgZbI1iO8+vq8f6B6gLwB2mSw0Jg+QAM8O+0heGVmdBUteA5AmoMQPIp
lTalUQ0cGriIXLbpcQJgSUD98ATwmRVFdft5XaGAA8nEYPAAOXLi4ZsWcR1ugMYr
rtL6N4mzsQmDDJoeRskuvQ==
`protect end_protected