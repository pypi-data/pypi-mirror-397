`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
cBJAP4KtBCbUVpRv9njlfgOghDSO0hTdFE6OFAWbNDnr/BzhLUX61NcNS1nmJChq
J8mHf4i3gQkqPfo3u3NAtFcMjcJMPmtgaAD0vTUE/YM5OVPQTEbAU9b4tS/QrUjI
TBIuF9REHC3KMz5AEXuZgMbpSrtOPTPj1GZjpwA4rAkat53NNlIM33WIkNX21Voh
f39+RkOiGj3zwWaFHaT2FCGQHYtXzEhGT12xmeer3pd+on2B+KSlszA7BVo4HrbT
/zpMynfcvS7Wyb6AZI3BRgROlpaANRvQ6zMF/UbGv/g2L76Zb960qKDDGuSq+m0d
yRtqBEIT02vLQeIziL0SM3GksczBVYpbIfz+djXoDDcYxl+SXMGhzltM70lZsWVI
hHpoXNZi37S6DhqvMGR4wIQZO4rI7tPmKRDDZB8JtfwwB4ktBWI53OxTrgsnAJP2
vsuJFzx5PfBujrmW8vTEzk8GCoFSTsdbMLWr4+X1dqztJ+DZE42lnpICmraM4/Ky
zNzy3bmelh2Qr6FA0Ry6NKxVSIIRf8Q6hBGiaWo8tj8ULvGaRlM65Emp5zrolcaQ
8ABEcw4SKoj66wz8mgYEQpIlN6J7eYqq6je6JZxmNTyB6eSCurTVa81uTJGN0ddW
7X9eomZwpkF9ui+QmTpmeO6C89czjpC4RmXIVfkPg+q05CyTpzwI1Fg3hXKTe0FO
J45lYaQ0VDqnm8PG3lC0Pd6CVmb92bZ5EiySHR2hQ9kWje2DsVjlcb1vwLQY35Zi
ku/W+GUwjT8KfxW9Ebr8fUv7+lqOynqVH6hoeGtbg25nFwfHqdHj8Me4IE0U0o1w
LnifkJrYuHrmgwWt2OsdfVmtGEIIdjDOenzlnQQyqbiP4ACY3jBtoTJykbrkZN9I
zcCkfYe6qSeAH23kBBhM1ku2K2O6usUwh9cACAi302C7t/WdJj6ZjjRGRnbJr3Yv
v9p/B6Lx3ZxpskkgqsBCx4YWGXuqypY3bKMCRdBgAxdKgG0y8CP3ErYOCtZH+rd5
ec0wU3d3C/eTRFMw44ah+eiP8z6ULvGTxxOaEFIt0MAVKRCAqv06OI9r9cYDG62E
fcXVc6jzladHt5oemYF4nDwYHIFGxsmMklXVyiw4d4YZWVlSSq/ypUepBvOJd3sY
azidJn9w5hm+SQsr26ZfZgm9Jx3ngkNtRke65i/n6oCNQ0cxQuz84cy4HB5AxlFR
PA/bDBq8e1uDWqFtOxy4MJIHQ0JUvNRkN6H9apWZLoitXUwUpqCL3HXk6nRtktt3
RUIYkdW9bTT0Nm8Uy9teOZziAcj0T37gq4xWCgcOJJMuObZxkdeFTiIjNHk0X0Uu
nyd8I1Tz8sOMiq2WM4XFr60csUzMVkWDc76da6j3kKMufmHFSkFidw4KU2kQpUxk
g3rymecpia7sFYGq+FeHxAIQQuika1ahJhwlg39CHpKtE/kzDCWNy5rmQqkmzYUW
YZrtQsjlgNNAdzL9sijSItwmg3D5PLRtvcyZ389fQe73N+zPosa+7nBqYLtfm6hZ
EuPnSgnXDVlZ6OhHZQbjJMBomsLWBfxyWJnF79u7tjZlO8uUeBLXwVrOlgsLCGSb
AKaP0tVSElp/s1v+bta0um9RodoBkmyvtn/RRVRXxIizwgjB4+v77CvrrDcFwhFR
gmA8cpuJ47Mwl2geIJ+zp66lHuSShlO73S6JE03R8sfxTekmJY9lM9RgY7VSCnXU
KZsgp20fiv7En5TOsAuG9IBkc3U/olyn4Y4V7Ch7cSI1e6qfMT4v75eZZv1rDI1v
whXnVcPoyNKRjNWoIRe+ewk+BHk9x6iCVb+x/7Ru705O+arlUFm9GBpybb/afdZV
mcSEbp06tAR3YmDbRm/bFRtycp2P9q0GegWeVqOJQD900aXTiGqG7x2SDtavMDDH
K46pupH964+QAZAFtZS1/WhYuoKYNL5JLBOeo+1OVSrDGlL+NPW5ckIi8F58y6/R
aWB8+BQa7XPHLrYgI68DLtmBHiW68dWMBQ+AS0tkAojk37EkqfFdUNVkPdYYSDsw
FHuTpL6VfqjRrg7W4itS/ozh7Z6ssnIYT88B2c7uTK19ed6JHGBXgZ5HY3THgH3r
0WvjUOWbTaFOzI5HnTEOZoikZpYsnwWj65q2KX3o3Fd6C5mUp/YIQiggCa87HM4H
Qy1DkrvLh5ms8gNZUPZ9q4unoaqUa+VKXeIpZV70o1DxvrPXfi8tbrmi4iGK7Ggh
VhpkNN82Qng2MPx3qlRlSIKNme/cnGvZcyCVM0we5OBpGjvcJ4BVJ+WX+ZFEANFm
nI8/kh0RdruYLPlU4deALVhauGm3wpbfIXSEdve2Qf/czvTPI2umlI+yHdq+K9/B
f8rj7qG86lK5+JJxj0PWyY2pLz8hLlvTxrkS19JYqvDrwrhX1Fsxw0ShaTVzg486
boDYxuACM0JVmUyiHFUxJYRTjVLW53GJzalLO4h/4s8W3WCrfjK3ZoMXIyEiHrCQ
plKdbUef4o8Y8MXFs73ck81lJfRtU+A/DTPRDLROrj4Qc+zKkgTA446FiqDqIvQM
zCN4tAv0GOGe2nytpeGy5HJ3oUFwmCa59Z+wK6mGn36E+EtBNeZgRUfDiK5/CDHi
f9fhgajlstDf+f5FOlq9RublA6TbmD2ZCEuGFEb7MEv1O4dsk4ZGue8TG6RsMm8M
e2to7IE0LWrEbHrGBGfavUvgxnKXqdY1cCgmx37TEr6pKc9sv/7IYtrz77K0+Qqo
BslMlNK3uuFt1JTYgU7dQ77Y5lj7pVbNgQ59lccVOfSfDRjh4Hcs0XptHUm1f3F2
uNZ1UYYDQBi9lKsrnGTVsuA7NeQ6zaUiNvCNnHUrx3pD5OGV4Sw0P/xsAfwAPyAg
UIqdyyPer+CpDNCwunoWIczbfWWTvSlrAPnOdYWJSTfv8SAyYTGOwmvVF8JqVSHw
Ks8GRueshsz2ukQKnWydUIv1B5rRIyhgmMeM0zKq797VnFp88CiPMe4SH3makk7Q
nNvQtDBxJz1saKodrYinjtXQI2zrYh6btmPkvi+ncy8A8EQ/05WjBeg+VEzconHU
gEcLE6T95og5BnpkXaJw18UvBHHofQTc2/l/o9o/+i1LKL2WVUDKGDXPbObsGPIc
RZUCVEcQSy6DyTXEiUOnhyWjkIxhC1i+rsUjGjepY83AbfimOKoFBTQ7Cu03sNJ0
eMr/sz8pVo/lsSjfJlVQ0uNVYcNJsDTaxbwE7QpHGuZiUfXsR6NA7xFnjO3pbR+R
xEkM7Q3v7ZlqTjWrtjKqCEJK7694EtL8INEhWv2YDVuh0q9jV/HdPlaVXW5Rr8G9
slLAMC5iAFtubeO4iYcA9llhPOg3gXQz/mQxy7BimJfTKGbaL5yTT+aDXy+hAPKx
lyq7NPvUf0R9YNtVUNOeHGl3ZtPRIcQwHYMF8Pnj6186Z8zWOwFzuuZocnXcjKZN
4i/mI/DUO4ZYkkthNHth6K9G/+Rh3mnbGHMo7Ajg9tUBGubu0lR43dlXWIcppaou
I51y9NM9Y5WcL0+KjZo69FLeYl/xCe9VpHfNwwHBisYzg9/nZFOfGQ9TC44V9Qb2
336z2E44DzLWLVRUp/pOCuaTmcYW8fuPIdkIzfVYNDBdviXvO0/IxCv5QKb/293b
bon/FLYUDSAiKjshfIQABFQ1tNENwtKKFu8M1mhC5XfUcnry+g2yCNqWJdbldOBv
Ckx3kLuC9uJ+tXK/xCh29iYvZk2lV6jE/Ug/robuplr7AJJ+6ehFg38QXRA1PggP
YWezpK8OsP+dmHNSUFJSafyXHDO7lSBUnUqJ6gWcDe3txihrJd9SQC4ahpRau41Y
VCZ1IxC2oBlIt2gK4ZMWyvST0TXIAikstXWUqRrNaGrzaMOJV2589BW5NbYpGLiJ
tnG4PPLWLWNt51pGq/NvUpkWAzrsEUL35zgbFh4vrP4XNVkFLtlznQltFKE17L9x
xf+N1vG0+MlcY+oR/mh+RKLkR9o8HGIVEuREY/q76/dbWdXeoH7o5BjGaCKE83Oe
9tsT+MbLeA8qYmxZL4aGLJAl8MPz7YIsPzsdRyPTAOWE4jL/Xj5RMrDxkaDBhbqE
NLc0b/qSq6mkSF5Tm2aVedHjJnWxpElVZ1HNVUrz9vYtV6mmxIUrDW3xQ12OsD+F
U6ygWA2mwmSzEmDEmlGXnD8BKFHmMnSh8HnEna4pri2G+vwJhi+CqeaGIiItUyqi
bIk/hOf+pLEq2EdaSycTDc++00FNnbRk7ynGNqQxF60oSXV/2K4iBZIa/j4HHsDc
Ys415KhdMeGDb4FWJwDA1PM9bodpeizB9md4MpLnTUkbU+61s0nJMu8fombfJo0z
Hc/AfZ20zI3nKN0YkFTmbaA4k1vA7W4CoodpQkFQE31ktyevqUzbLxCspoi9/1PG
FzzrIS89jd0YyZ2F6mAlClTUT9Tf4UJ7MYbgXxmEWwbnDTW4JihFmimWV/GLauEx
eSWL3xm/QOH6Jr+d31umQGCtTGC9gIZIupEUltTBnRusEVzttS87O20rs3kqX67T
nJg7HGbiEz2GBXn7Vgts7/qICM2zrZ34ADSRzC1HFTGbgEUbh8MTbp4+VUwEs9nX
ZmGY97qIeILinpv0ypLaTApWzvqH5MaLpFRjsdINddUjtsry53KN+RWcXcBSFXKP
mnwXJqatcgUrzaTqMCx0rmvrh7XNyeCLQcrxouJP+C7hNain55c7UJDeGB+uvbGO
oMZO2MPcNLN3r1h4+J0IRhlFaZib7oQeeppfuiBW6ymU07diSLSLmdKir7/YLWtd
ay/f2cArhvB3GiyCvH8zr6cFVatvErtfcCdMOMe/OkkFx5K/gpKUv4vIAytScAZO
r6snCWMZcSp1GAt5FcL+k5G2NuAOARWTySJwHGZU60E9VLYLoxaSRHPACZZuMf47
+SiqPPU/QOEMIJJ3gT1RjQauDP+O/9C9itMteY8GWgqFQuxrPUyHiR4+jew76UrZ
NCbyg2pM+vjngO98PA+7bkyMzWgdI3kZIE8oo67YyhXYrWQfPWV0Ye4Ahfk8/VaC
OqeMd85CqEWYk1VRAPytxecsOg+U3HtxnZk03oJoErH3OaPAUhWL51kHikHNYukK
DH6tsK9+qC/5QtUqdEytvOAIGNFttlzCLu0wKu5cW9xylIKVEwF1ZUdc0TiujSlJ
6NwCKyhbJqWy1MzQezuB5/lYwxJ0y3heu4NNM72RV/Zm/k9g7yh72i8OLCURWJVC
DY+NHbEZXwj8SiyO14NSrGp/BVsynMjWoIj52CaBhmxU63pefVZwK67pWKHpsi63
pVrkQOP75uoLaT7UZCpoQT+aGMRB5Us4AVcplKFFdeEqvW2sIAZylWLqCi3j2ou7
QaGS5FJ8AYPf0ukO9Z6vBjGNs0b8cR0ynBAHAFPNPSFUs/nyrYT243mZdzXqx3GF
I4vSUkMWb3pO0f8lf9dIwiE/w5iRLWKFKjfDOEFd8OGQ9QT/uJC+3HNYZ4FWz0w1
gp5x1K6X0h2qKyijISp+pnxPseoGs7M4rcZEHUbhDiq+sqWIgo1JC12p6c3MkCuh
tt/u/rHqX5dOfbFM7WwDY2vNo+FRk4jTR7XkPSe+u+6QOAhP19G5sW0g3PKBOEmp
awJVg9u5Rt4v1qmw95+EsIQA5priJVw9vcefdQvwclYY5NrKhudu2NHFUGAjj6r3
hEJ/NLO2Rj0V0P3x3my03Zy2FnTPni2N7mb2s1IZeS1OdeSLdXI4vxeI7tpNq5CZ
lJ0sKB/EfKRK5CE4evUexszOCIxM/QMfSDgPeRgOtt/UFWHLP/Ntv6aQkof0c6ur
Qpjc7u5Z7JWKCol2izoXzjTT6l22Yzu3Gnp5AS9oIixZrIvDPkmT33tv7z/W1UQk
uL3MH9a4seSaciHCqkrZ7M1fjDHwC7h2tQtvoZ/3pUi1U1sRhVJQrTaqHMHwWUC0
qntatdL7Fb5L58pV3J+YPpE617uQ9cIyT4VR79KglO9/1Nj5C9aoKadoyIuSfdM/
VlGg4Uu4rkteHhGgBM/wbhwdfBUlZ9ODDwOKOTt2m5giCdG8JZIa/bC0n71pXVuW
KKQlk7tMncAiEVPHv9WycEXhaWlxfr0WNbp7zTvKZog+7WDwOATqAwkgK38ksP01
eLhOSk5OoyzyI0wB3+uOLFgGZPRlG8gLVGQy0dErEHslux7B0Gf+uGq6bw5p0B/A
7cLsDTTKt7cPUN+/950jC5q+9lFKOOfEpP+rsRhWFK/09/dU1vwafs/YpmuhHrKB
oXZrV7+BpWkfn8qzKeffUKsAkqVt4xC4Q+e1sGlEs1cUwO5IRbuYcaHrNBIrFUrp
clQs5HQgEPZxyQQ3adyuQCp+O9ZP1TAQNLoSJi1e1sxeszV3oLxW0tZiGgTu01Js
qVH+FxvZ9yjC9VscBZdxWxY9QD4grXI7TyJ7j+1PlzdG23iWTV3Umlb8uNwuCvfx
8qFGgOAngdTdQUmJ6DZfNuNyQqbh2nJbZ+vMTIqhdHFHKdILjBCuPha//DvVVp//
g7JmB5K1HLuTPgs4nRV42ZLox3LDWHaUz6S70obnl1HAtkJ9GlGOO1eeWPXMzp2Q
454HoAiYAj1I0thyNTQMbpbj/OcwSdQnC9K5dlZgl2on8roxwENDp6QszuLF+NaE
RZPv8926FWnQK8Kf5GqGTuK0VCp6/Q9T9w3dJza4to5twTjm71Rmq3mpMlPdAN95
rrzJRaacN60QmPm35lhDlmLoIhXYFssSmw7GM99uIrZw/CP11i/dRHT0pQZrjp+E
V9uCQk8FK14wl3XvOyPIovCqf0XMQdACyJoZxvxAx1U4kdQpwaeLfRT3b0J0gGv1
gqevxdfIjFQNzNvRwhqXPzlO5xB4ZfpZItoBjRDMSSlSGsRqhUJkh5hd9vFMeU9N
yljNmeixFx8ntIC3X8x3fopdYOG6TR3oChjXgYwFERWojjnWKcrjZq/dfFB07XIR
yZXlFKAJKxKcMsEgLBMMYTeY1iNMqtHs1Wr5s07cH+nGa8o+v5uIR6k7HCbWEC2M
8fjFwEGlkXk2YSdWaw+l1h85JnJcBJVccA+S5z5ZNowZqQoqL8nj3+3aq7mdNoLZ
iudYNn6XcrSwABDGyUKgnI57svZgzTv+mPqbT0SJYVHLQ0Bj1bnf67iFRXq6AR9L
FQKSSoB87Ww+V0rZ2rltOCvT9/fy6y7DkWai3/9yl0yedk6YFBOvvV8yadDoP8vm
/w8zCgEqyO1D5txcHrW+JioMxFd3CwbGMPfSRUmFNVX/QszJ324j4J7WHUgKchA+
ZU7OJtPx32+jS1xGX/O5Cxc+QqYkalzswqWfwo9Mhpa0tKqjXd5kXD+5TBQexsmA
uQP2mUNL1WQmCT8EemoCunoe/6/LNYJB0bKSItvOhq1OlsNnvF61sGpV8tvxf8BI
cP/bYXSByMQnwf1J5jGq3L9TYqkkS4mNbjNKXLLQ8uJJKQEQs+592qMovEI4VoA6
IoA733RfTrX3RnuJZUlFtxrTFoqkP3FSlAtgPNY9BMnZy1gak6v4MSz6p/q66ldI
HDbcGoB/y3kDj6icKTAfsUmE6p6iZZifvQDgRk+mwIo8bcnm+1puQaunv0GzLguX
2h/8IuJEgHuPPVPNFwBFqc3QM1YZ1kqSBUmZmwYQAlep4qzAK9rIScUrN3B2vQRA
Fyjh4QRRJMEMjMk8cVNBVGYqwgDGepxea/G9UfluuB4J0D5lSO2+rHrPh6BhnsHM
y7pNjbCIdeO3PmTLcsyQ4h8lNItp9MiRXPna52n+zZupRTX2ioFuJAEYWro+FraW
tc/j0YtCxJ9c49A3ZX1bd1BacXkO4fp5tYsUWT4PI9g732tJpQlfBXQn8d4TIRhI
xwNQ/knEb2/aOwPM8vlt70YD/wO1w6mZRqRb+3COnVQe0EvjtaQoklim6FUNqQ1q
vPq3OV7hVdhm/SXQFWA5ZMin2WzkjRq5KOTbJvdRHm29n3WX0B+x5H7MX4S/SHPi
zdNGRhHc7QItO1tJKSw4JRcLRvEJ805MNIc96irPV7gChFCC/D8t1dygYU2UrCSA
WOxVV3l3RiUDB0Z7NCUugsd/KWAHQl2ixEnN2Rd7OM6VDeCB+DQqv9GdGDNrugcA
ckxHy4nCq5AAi1FKjy+h8B8Rb6eBl2VuFsjP8dyHQsHbHi6Az9DyYpxxGOEXb4gM
gSIB9FzBmVKTOwa1nbI0pFvuXIwayE5V0z8dt1xPzsJbNMzJ62VWT8c2Kf6es0OQ
HKOswGQDOFet+cn8RPwecRwQm0MxPhrcwhbo9Mm5kh2kVd62yII8Gyty7psXts9J
CgZhWKRTclQPQRJoPj8tsCnwif0oQ8CX4RLm/XkrZMMSrV5c6b2f8wcQBXPzCg5a
/dz+p1hruZJE5K9ApkWhyeg5VwWJN6LnDSCJrTBlx3yy08xtpaTmw1H6QCYK/b+K
yNlBzAfgi/A1tXcj1hsbISx+er94+rKHUaTwxJrtRuSyoXpj9r7HdrT0IiSC50KM
/Gn+BkgbaTSaWkXVGfvxJqIPNvAdl475xQYG4d8tHPf7muWrm1Cs0pxlTJBrpXyy
lpWt0ZL1vsXT2MQDSy7zPZ/LBkwpSh80oBH17e4HNh8lMVxfRazYN2ygBsPzj9M4
gAnzSsZWTyaKqyEonesLik42b33Mt+KSPr0ukXAQFpuc9piDRDuVo6/OBFja8Jep
/QR5OC2coSa029djf0XiAYlJ4oJooeR6qieytgotsGntO+SQSrnBB3i0A4pYVqmv
NPiItFSVTEY20zPGKM3bM0eJ7hDPcsMpOheQkGVWL7x9YFJ3y6DtETgUApDImlL+
SK1AkWy/3wRzvsNff7gWk2aUaWPk31FW52d7ag5zQ2TpF2BBmaZ/R4sSEOXYA+1g
XSc1JDEAqgtHyCSEm8yC0gYSX5AFol+OEwIgauR+rPltIoWdcddImYfzBzO4YQ8v
DEX46rEU4Va4wxnNP1TJQQd6E2fsJfQTDCHAUQbP2CwvlMbXgA0PBTw/GXh8zDnx
AhyUK5jRhD1iDSsqGoeDgidwxqvZNfKt9uUgIGWuHGMmc964MUbhscpQbBDCeI09
Kcy9yfYth3SBq5HNjObCD2Re6VuZx96MKqs1gKMGOFJjj7APJxLGBoaVMgFvKAef
KpgN0KbsxyhPA46qqwcuDrwbC1SS/5X2eJxsMSzKWqIEZA1OkbXbE5eQ+Ip1vk49
Fm9PAUseZJSJQ0UFM5Bhbdec4O44tJ0LT1QX6l/ATAOmzfZHtcUexDWR53SuWolx
DIcmIgJ6u61Hsz2b/uVdHNCXrTdie9y5ts8lWBIXCbXRXKuqgB43ic2/hMUp5SlB
+JQww0BNwYrwHo42AhrMldvXC+cW4qlYlrtfQReR2JVE3nQr2JpfJ9G3OywDbPDd
wveYsO/OG6U24GOISMiRYYH6sUUUISYqqGyHmPPEkNSR1DfY6UTteBhl1LTmelse
XaU0icA1XggP1V2z7X4zyM3/nGrA6LlY6iM0cvWlYM+a6Cai80Lh1b8m2sgkTTgn
RaUjnmUtFK+fqtuD3Dew7s0NLj5IlUyEceqGE3c+VejUucYmvuy7zV8mY65womS0
AWy99PtFbl05YBTSFSa6PlUdP3JHlkgqZhKZMHQ75fnOOVt1LSwv1/fRrH8G7hJY
3cITXrc4bOYza6W8dWEvbJlCAOJz63Ya7VBW4RHVmHerkZoP/9vEz36eQ228O0WM
i2H10T+DpgIOCEg3T+QfvmJGu6tVcsSNzwmyWWCWyBDdygbOKzfuCrTPBotcLU/7
VfNcst48do4Hujt1XwbpcizGE/2UPa1lHaMbSt3/2ejmezlTGOTcrN9YTLnnKpqp
PCwWj86eHZ7KnrsofSAcyTn8t0ycTH1Z/T+acA0xL8WAIRbHsqDHlLrNK2H6Aj4o
WfQjYd+5QEG4jAn5notUZ5gzbZHRVdI/Wz63Wfem3o+tsfjGW2TXyIOPzJN5MYAk
cF/1U2NkQcZtaizpz7ZDIEvmVr5NXLCBx8uxzfvwrpn80KtoOblJeo6+Xd1TAIXc
+yQ6rpHGsSD9OIoxsz0DUG9/pBedmtyhrF8ArNUcPKKEXQo0CqIH2rMsfxkk+uS0
bjD8q0TIsUdEFoA9LmwH/a68+OntBuY+VCmtc/J4Sw5ncoSBq39yF5C6Q5NorbS9
g/ktU8jaVRktwackh5W/dhlOVGgiDnO5XPLaw6bLU4vMeI6B3slWP5ooU4QyVQyC
pagAqY+T+fXekzekDGrK0BTOnRoqtYy0qsU0xr7TsI1NgYw3kCI/woLnKBKRQlfJ
/ntij21EMAB2AvkmG6wsG4RqRlw5j319eVv2NPEiAKRiQ22LP2DqRgN/fJ+tUl8p
uIWGxcWbWrOkLyX8pDD2Gt4Hbm2YjP2kDuDmg50pMl8clKeQhFyKXtqBmFkq/sI+
ugwaFLA3EEPSztGVONfhRXnznIZk1JixbrZ9A/otTuMhCquCngfNnB9Xb9F0I6K5
ALKe+hhIvyv/5rAjIVF8WZ4nXv+T5pg+jzUaGVoAl3Z+xX4ZR01wHq7YK340xdPd
Drbck8T+GL+VwLJBumfrANno3aAFPURbGuBfbFUHKjTYPhdofH2Z9lEXAtYC8bTM
Ty0ufIWa8xGmyVeh5M65K4Q+URoiu2eTEtmTgk5miH1xqiTuC8B92AGR9aPgl0WH
dyOXnRKr3+SJFEDM1Jk8dLkFZWNmBhjyaFDvwO0v0fWRvsyP5BzywHIEgte1otXO
7S6TmMbTUpiggUPU2INTwGVIFrs/zrJTokcxl8X4SHsXx0plcP0umyC/2OqVtB2M
rEEpVxshN2iOOKbP4FdWt2+2TvGUpcfQseRlMFM/08pTX9wZsd1Sh7c/n6li1t+a
Z19AwTNXZeXSYmimkPvbVsEAUGY5nszoJUBSXCMSAslFuoHXeDx6S49jpYlwDRRk
zIL5QbfoigVudsGgucxKYSLxJ+hfu/r+p1WyiAeidI1XMLyhEiZMbvkj7cs8cLpj
skwq1mDWzrwyExXHEDDqKyeHxIUHNjsTJvWpToKGcAOSI6yysHdP6y36SOi+sUM3
IwNwGllv+Wdu8CMgAvkDn8+tx7tzZNQIL11E9DoBEdhCiXpf3EnyWPbh7Rfgc3q0
dbCh8QlSGGPELCLTHLhUZ88M4ufbXBZD+dC/VjvxRsSz4bdqN9eJsyi6a0j4aHba
rI8FCrkj3oYnhNs+PlAJsMwxCYJAD3BpvcuuhHngLjLaAVjcS1TClDOT0xY/ufpd
tI4lQPYD3Gz+ISK1tZL7JLfDuNpyEs+PzfvagK0RmWt8knRlP1mNRZd5xr/2yMmk
JEoQUxetEZvFvAffCA+/+1P4lSOtUaHfFFbf9Ux5pnd40n5Fg9+z4rnVq0Gy6E74
bJlIa1km6s5Zy8ApvcCct+gk2pxm7gix6stZdXlIgoyBAVF08WROyLjU7xjZ4iCY
5qug+q7Bf3E6CTnKbDBR+MblI8FGmVi6v82hD4dj/uZP933k7igUwXt3z62kNhqR
uV9eAOdzt7o3R3JoilQ8E8TulpdJTE1o6bfEnmdL/1Qw0iv7ZFF3ly3e9RPLvNWD
3qk3ekMWwvulXuy0NGiCymJJbTRDoYzi6NzP2IzSt6k9aG+nNKZFQcrKmrWwFq9L
YWautMkJWPaExVpatB6vwAMJrPCmhJuQ6J03QgJVd3izD1PJGlSz8TTxoKwaykXA
or2RYGaR5D6qcuAYW1tn33pWNefLv0Z/7GcbxlSbHlAcSIoE9QuR1XLOviZvr9Gx
0tjaaX0dFWNw9dpR5I61DPU+UCkjtabKvv5XjrNk9e5GIeAip2EzqLF5+48nrkQM
FbGMdSLsJvRNPoDDdgnBKVezOwUu/0Wb+IA/kVhL0nlGZSb7MaUFVxF37oV2QpNI
xI0Ekk6YNtGfL5O5euS01zm304UmtXcOyBCPrXv6Ewv/X16MbprWcZYaZ3ua67Hm
JQHOMkdB/A7DIZPFkmRfQ6fvDLIFeja8mlhvSBKvw+F2d67kN0hN7FmxBeMnBAFx
mXGl54Ep8aQjlQ5y+v85YdbEnZL4romVuDUmZbVGQgYAEVUw9d3A9KPyXzBujLtc
MgCpnc5jsGHWaSOI2E9DIqryYfRViyU38KEB99A/c/3mN6dBc7nVVNF4kWbExwCw
g2mYyJHbBXNnLRsSJ6BDu2qwVe2CisY6msRFtp50Y7y5mhVKRg7oIcvakV7U7RWj
s5rjs+/LOewxJPyah3f9i0pu4U206xDRkgNED+INblryzGOEVoTyyPxwfAm1s373
ELusaFUMQ17sUYTlXfFO1rTNiRoZRUZ/t/NYrh9IxFOYHsGtFkKopKAfZmSFjVpQ
+NVJftJo/tKMwlT/8sx4wnYaIN/3wixvk9d6z33sI9hR/wLHS+YOF3QXRi6GLU4T
GekEuu3G5JF+rST/iDqB/GX92liJpA2ULtf/b90wzDetsmr+jVGGy3hofypZBVmi
EXTlWeQHrEMUJ/QInwyFXDQcfuSpyJOcWTDMb7/wkmZ6P9HYyNWNOJAh03g8YFbE
BUgMjJRK7bH0xVwlvBtkO9IjzNY3NzGehemVGos92aRIi7LeY0Oy0kjrMHL/6IaG
CUVmIkFoGglWoVZbu+diIJMsYH7bg0vmZCqWwBoY5kyqG2cfk204CWSSaceFJWvW
Sw7PeolcLk8C+fPOwEJtZvzg7Xey1wA38KsPRHuyaiB/b9xiBSML+1RYGttPVi1t
SQtIQ4Gx5FK/tG2e+BOZK5/ZN7ySKyR9XigiCQogNh3eUpM2WqGzJkXAgy9MmYy7
AHGT/yYKEYl1lTu7+Ytj1/dIgxDTLNovZZMv9fnikU5NGUDWWbJeNwcqGuewPvOT
n8yTA1j0sresR8yrpVbhzNMZXCAe+rinsdr1hh0hVMMa4I6w3QtNzl0rBcmiegLy
PmKe7D1lTAvmYlE2o7c7FrP8/EHZT3vgcn6beP2+RHl11k6Hojr9XM9vkHlt3aZ8
KlwTBSMTDnjjYX2zvIrWfKhGnMTQTJB724f5hENVpLP5welVr3Opdy9x/yJt/QnA
OuCtGVLULf72IlwddXiGEBUAJ/fF5vUwQ+aftmkI8pluT6uUfQ15psTLHEGdhB6N
jjB53oILNcrVvT+VtzSUwrDuksVSBqEsnUvE12N5+SH+IYgtKLjysdDWnybNDY6p
UViVla27tM4gZMswa7dqEAbZh9lnMEUS090sLkmcmqYTF+ILoCpAb13WzjZ4wP3M
1aA0L3tJZ1HTkDVu8f7uAmPQNuE6HxgvsgctbgQdYYRBelLzxiTuA47jIyW7Hsn5
PuaTRNbOTCBXOwW9YgXF48qEYvr8LQDV7tE0lFEO0Cq/X+4Vic0HgIg74Fdbf6Qk
/Ij+S5W7i9QnwwC6JRcnsJdHLqpAQMb2CQuDB1t214KcqUE4VViIIg9FA1hIOguD
gxoginxo2KPpt2ZWwlWfBxUbD5rrfmahV+n6v2XbNQWVSkuGHNhI6MS1hwg97u2j
igxW6mpOQRTtUf16Z7yOXhfZaDtqaucxB4kviCwS/i6pcujKWTKTaCjKWM3yij8l
HXy1W+oG/NhjZM1+44He1OFkE88TzERZXQtZYjwrjzu4udi4BkkTirHJ2EauxyvI
gEoHM3uiko9+rq4DodniaQ05K5A+KV9hp/Odsw6KEeoICLTOIaHHXYpNEBxtjkaY
se+ne2F26a3ezxVZ+6OkWhtR2rsc6//D5hHDOx7UDdXCp6+FUuYGS/xKIpWL/UjM
bovF6LINzikRJtqI3NP/hexY3s/sAVXlLCu/aVI2ZC1a0xOG1Cowg+ukS3LJFu0y
0AGWz8ajbtRTpORmrS8NVrFkhGzi3GcC86DSLP5hVOJOilwxrygkET0UkUY0KjXW
12KzbiJc1WZl1ZloknVOh8GPgpnBy2ZMDlsLmKTKbhT4VVRtHm7QFXg2lHnBsEzB
6VHP29chIuDKi0JOI8RT/623AOtb6VYcilF+4e7rofFPzYnQql2bAEn9jCOP8uwv
16Oq16fitpLSJzoUvMkPs8lbzikxu+8x1E5RXbB8uIbIQQ+d2Y128u0InUWRG0/A
RsKnN1uPM4LC2Ds+SqZmoik2k5izwD/c40t7L0urcQoD1ilhYrmmvbopLw52Vj6O
BfaaHX55P963qNgzR2DV1P9QFTsKqfpJiwehgZsmDQdP3IWAF94CeiXh44JUwZVY
P+v288M/jUYlMifR/dIcqXCbXxD2b3vZgsM0gwOhQN1T/dm5A4LYepeXpxHgCe8m
P5zSVw6ner41Dm/rwjd1WwLLT4Avr6XvWxm7WxnoqOQXiv7fKWyJ5HG3YYzxv33c
u3m0eRKfxTIq7jrMBsN3n12kmOA5xDjfaPX0kJFmK0QmKh09rUiRhGjD9W2y88gw
n/7L78gpIY+0UZWQgLfyByJQpu8VgvK+ubuuXU/4xiBCI5tYfRI4thGqahSEYwFy
UiLHXs+NcgWr0zyEEYEyGXuAfZCDC4yAXtu1P27L6mD9Hz0ZTAdxfGWl+HtuTxfs
Fu4LYR0U2MwH3j7566XishjcvM7TkHSe6XIw9c6D46RbNWAy9uxGRE4MMylgyhU1
FVfVgub/dikMxnadNditACuRp/CJl+VclNWJdtTgZFCLcyG8j9vUt0aXr+vrSiuq
HZ/3FlLC6H/sZB6IsdkxQIO69Ngk+Vu5bjwIOp1nqKhjHZzNswkPP/DH146X0oll
pI6pQTGvpsqtBUpYdJqITe07vnH2qA13VHCtiQkejzHpl4ayo6zWbJfghcao/73I
2PoZrXC/qGzTeypLm9mbiW2gWhHmnTfttvaScwWgmsJlkXLzZ/VcyKds+qbm52bk
jwPSE/MrG70/mJYXkOCgev26asgJ0LA3Z3ka9FafK4N2ktPqP1w78cAfA34AbIKk
HJ4eo5SnfGz3TWXx9R2SDQGp0bk0hsh35lDuNuz4GPY7zEoCozgtBCHmzij4pxsv
eo0v9b+VUIXaVf32xB6xfMQsgPFKxFMg0g1mR+aQSzX6Hkqftsa2i5e9pWp9s/2D
ee2S+G7NirRc8gmBMVj62n5tzgyR0aN7RBGZuP698kKW0wTuvefrvf0BRo9+1wfL
GtHAzkZY0iWj+bc+rd4ChIcz5dnRqUXNCZD2+eT+FbHtuG1MPyTlFHFgp1Q03R7r
aj36NBzoe7idLx6CVFV5s0L/J+rfAGN4lJ6tPxLkmIQYjsJVgZB2mdWVzR/NZbU2
toGNF8VPOtd1B4dxF96Vn31we0RxmRU7kwfLZpS18ryjn/djRi4juYqVxcmL/qe4
10LA5ydshQXhF6DQpMZOP8DxWJ9nmlqQYGzOb9WFVAsvU6A8s459ZM5Aj5nkfQvE
pu8FEOWsvAMkwfYfTMGwx5HAncDn+OUdXsuXokWQKnAT+3ds+XcQcnEhuRQZ1FJp
J8WrmSb04Wa378Rg4zYwysWgMOCyq0TkZalOLfEuPWsPEmTi8Pi25GNuQuYbzcf7
PO0yTSwX1J+xpZvzomL0nlqforOHBag5ufAnWMIvovuTaKsska9ul7ObfgpQAmci
uLPl8SMsKgG9ZxcCK4b5yJYs4+vw4t01YrhxonuDjSxKQ4KrhrUWsPUw1EwMKv+A
nc3te7q/P4C0ZQrpsgiE+gJP/L3IhYP8sM/2wx84IV3QAFoHDCRkdUOSNOPs/Dhv
sh5krjMLD8+R8ZT1ddH62Jjk5KX+xkheiCdl6ma9G5wYmzsO8lVvMvnaHMIE4vgR
yBrlF+XhE+9PGyHdfNWCG7DeecYlCrT5vT4vCwPOiixT54qMPTQHmpeIQ9X9FQxf
CC0jl26BcBRItBUGBQ1r/+xDWVjTf9lo44lS6fX2oaRC2krHOymqjNXCwjlsRlUm
ApWQyzA0JRgjoBJeq7ObLOQXdUd+ZPwXw4npYWQgeRdIKWDUS8VPoNwySG/KIqMO
xnkjQawPagseTEKBX0dmKBQVb7egzTIZWjdCoMFVBDaGg0oeF0AtqYDOH5HqBvmi
fCUnyvi8htptLAURFDADaawvDybyFLVEKMi6CEwqRnH05u2UCT5aDULO4ZsR9AU6
7ZLh9x8JAs7TMXKhVcZbvA0UhJCfPPCZ9l+dv88ocPphnrzwolWBq4Td+2wwvVpq
FH3VrFpxaS6JY3gZWcxpFlTHtu0u5Rzo9Ppy3PsKLfe2Kl60TJKdtiHJpkx4uvYh
ZkI/7wmgCqKaTPfEvHkKxLCW0O+zw/aHV3qjPk5BYSMrwYxoXpMSQNVf8yIVIgNK
guAgTXkBA1lv+XQRgjKw9IV4X6U+jZcEaZc4HsIDiOqsF7e/QWmnd+ziXCRYa/D0
wr+ltSqSrr4U//VGAMENOPD1gsyrleia1nC3a9XhtDoM4DssVVT+ErcdQb+q58Px
cRxmEHEjv9LSZfS23YtwhjBcikIqmbcS6inXHSX5kCH9RP7WcxyUiwqfERd1S57S
mUtBpx3ie6Yx6+fEutIGg3ooDqldkpHCL/OjpUIWZOtqmol3Kk3VwktN8F6r7F2s
svCKEs7SaRpapYx7vnq/YzTouN+FnThLlukIHxhe4T+J1qGXriqTBC/5hhdCWqal
afma6gnjBU72iayrVqxDmBubVZQmJPiITVLqovB6y9EUoK8AhhfrF0M1MaET5jSl
/MB8tE+fdn5syGQhTfmaKTW6Y8coNz6uPaiH/coMeRgWzcxw6suzmMBKukKwyX0l
pa3DvnyobUYKc5Swg6jf5XLOzD0d9PwVI5E1qv2tBFGn+aVEVR9wRcudy/cGbHiV
mmJ983HUNtFi+P9szvXILfMjDxsuQiPiQ9BCO70Wv6ikwoUby5LntgzatEqGpeUA
6pTLuYVj5KpWUjvDtDX+Pdzlju3qd/2G8xm2a9MYhF9QtyuZGXzgWDg/pVZl5Fb8
83EtveuV+2Z6VrvfeI3LElJmO2ef3KpQmjWCLaaYOS4lnTeI/+T0r3vyA/s7ZZoG
8FMyv3jWqDruDfBPj/6HbgBW4tefXP0ut7hocpH0rCFEn30xE11oT8+yY4LuAPru
T8FBN8gvy5MvimPpyS4+SioomMXHbcJMe/YTR7GHp+ZvjMEkCsEeeVwLxvGRZ3kx
dLDwd8Cyatu4moa6OXWOO2rJaRtjvFUdOlnmXBAHdsvRVVkDVaEP6qcdLR12t/1y
CTZArBpOHNDFI12kK5HLDpe57hgiaC5DSAq56pk3UqKXA04pRnGVyFkK7hYoYNw8
oDT75sHvm3bJ014Koox3YcdDF9lUQVAubeBQa8JuT84egeTN/P0FH/o3NPP3ZX2y
x2uWT/JQHT2+/1nrVYKheZdKHBbNRNuBCRjfeCxm6k6/6tD6wwFdDVG49mQv5Lrc
bARimo9EgtuyoMX216q/Df1pE5hVJBKYw9WiVFUXTkhbyMvKZzLtFL99ANUZNQJW
rQxg83V5kZnVeNut9wW+SoiuD6L3fmjb3dTWhLSxTlTRVnC9IePoog6Jp1hRK7wb
W1NFsxQrww/LzxpyevzldDTVxVsntZJZAZk88WXLfclQEsgai3WI7tnbU8X7WAwe
XvwmdwxXk5t5frjNRnZsqpdwU/HhulwvJxVR+Ucv9JSYhUjou/JQmr5quxPheccI
OldKPz+wEyp49lip+6igA2EinfZkOPBo3dUX6iN9UAbbJOFTVX/lUZLfnYgCmzef
lNnWDXSPoHnjYq4Z1lw8sNPPyFX898CHcX7aH+VmhlNG5DTIGrqk3n/T9c6XuSgc
d7IRnELaN7ieOUh1IN8wOwrfbo0Gfx0UllNeLoaI81abF7lkaxeubpMJDrg0Edhu
eIyyBpLfRgeT7/u3WfbpmVCw303OHJmwa+UlSE+Jw1qkbIayRKvSjYSxp3wq1cqI
dtQpCAZwaesr2re/xu4N0ecbqVmnKg+ENq2+Nv+pH8yCrZjxX7sH8QrGgmdQCXdd
4J4pDtHj7OwzNSbBw6h6SQf5v0mtrxx7QJ9CsYbwDVaWl//r68tBwbZpsk9RnZti
raaxLuwAvgLJuAGGXQ50EYPC5piJ7j1YobFCdBY8U81F6NgNCFP3aBKaWtqvKmoM
sqOTQQpsXwl41IHdLh8bk3Xr9hGW3cWPxz6mFFrYBesUDG1xcdtoM5joLfzVi50r
RzWWqv/8/xS/a824tyVAwKUun70N3j5c+aPGsLPZCltCgQXtEcQu3VYsyzmutcFq
Gt0sMpF+cFnCqqWGWGveadQf1iL/bgkeayt78aZdufAfH55oIwy0A66tZp5OWdwH
ogSEwrC169EX48ICevzDTdTeVf45TCKgeKMNAa1uvKaBZ0RFhTrUu2npf7qENcjI
ScdQdEZUiSjusG6mBkjgKhQF2TyteH+B7F/Iv65zsYMWDpmI4jMMpvzs4K7i9ZXi
413Sz31DNuDKxce0UrTexcGmv0Gjc1xlgVWMJEixRBsUHnj6sFEs8Gcf9JCVyj1S
UHoLBfJB9a9MPYTubVhDmhtw2Xf7iGON4CX01yJ9vWjT6wwWDWig9KfZCEjmxzw2
PoX8Z6AGY1BR67ebeHZ4UWWwO7tMHEdHMzS3n7Y9N9Q15UIxbTYzX6ylll4dYRz8
7lQvZdarqCZaIIoj7YlqnWmrTYn+lMT/MRHxZWEjYhkG7H7eXUGfqV1GMUuOtBWp
O3+yI6S0vMwTLxXml64qajLUoTXBPSHCk9+faMlRTWx68c3Tm0R6tB6vpWanavl5
xp1J9E7uq1fCwZ5Mr+HSXqf5pTIckINVW5ZsKnm+kovyIwYeSubDE4cK5So2C3GH
tYBO2SipYCgr+MoDM7G6XKNI8U3PI+iOy0pM0y+jsj0ttuY9Z+1euaUsenhehTmN
QlmrkpKLLhf7toKOdwm9XCmMSdbJdOivNAqaIxudwQiMVpz8ElPaqlsChcFzXH0k
zmxO1qHfOuxQKQHMt1PZg3jZJgLJjepz7kZJE0m8iYCG644Z5qYva67SnHAmKftG
LBSl0vNtqHEBz7UZvcRXHYsjHdF2Vixfb7jk7YRWBIWAkNysz7cjMfV5AGwL9xH6
I/IkoBxTcmKO6oB/2qr1GC7G1oVXacuiYJhggmKbg18rYjCBRRyvEYWNVmGFLooj
v3QYLXts8QcYxUxajE4v+L6IWTfRWYalno5P9oQV2LZg6bkRnXT7ORMHY9UE43+y
2L4JFz8+6vnokzaHpGhimUuEPaPHuC5xqIVlnr+8+2S/HDIn35fqryigpqoqYp++
fDuyp+dTB2PHfXMYZ8062Vla6ieNgTA0gst10QzXo9e4D+Qm32Bc8iR909m2WZwj
t6uQqerebRyQe/fn1eux1E7oC/Gytl0KPaBMg8WVMe8iwlAVBdD56NyS0sJA91XD
DIqx3EH4Yav7ZMEpyErfJT850XaVQ9mcxh+ltM3G92cscyiyQuczYqrnU2ntJ5Hc
iexK93lfOnwTcr9/4rVmZe63in/OvXLi2x7m4yvjSFhSOb7e74TE2rP/H9qGyDE7
vkq4M5lBho36O/VkYQenUUCD+STJDfMR0iGjhf7r+qECt48qdoD5KCi0IlSA3pIn
4dmcI1OvFFQfewKgkK3Y8KCz8gYOPOnkDMDG56g7IHxRkjHlLOrUx5Q1ju27pGtZ
oZ0a9uXA7Kxi387HDCrZW0k0K14kfVEq0jAeDuXIaU135IXz6XrMBHlbfPSbEovg
0pYfxmzrQE7P/eddvgMDxsmMctPTrt06DX0ip483BLFlbVrKex6NjEw7PDZkx2Z7
zDXgpJqCbNQWBsi643doBPYNRPkyV78RmUggOh4KPwo/VpLcJPpRHHG41PNoe6sZ
dFx/x/B33zJmzFSurauGbOd63At9z3cKRs7zQxeQlvgJnkGfK+fppneXJnxxoJfA
32JgPsRdgsGdfwlqU/hkPP7VXsjHL5pZecDxgP0JLDjk9pVh+0OeOCv7/wn5p3mP
d7VkCuq7uqTLo+oDRJJX9v/fcjQ7ysTMQ1xQyHAsKaWzNvIt2TG17DFFg2tAjgyF
YZrXYQmfakDxqajO1B58kpaUR2UF5+qFPynEM7XEplLiulUre2T379m7hFLALMkl
XPrqnnXFFrpAIxf1nIzH/qWRTlvxz1F4+e6IzbbNZnSI7qWmo8c23ppdY1ojEygu
Oh8b8NE5+6OnpfxbjdUbXPsnyg4Q63LfnHNpsL0IOVRLL+879yzkSz4LnaijjDlD
mU6xNBgGDlA/eJMEAUfrwsI/txqK8EvVw6EtbOIF0Bc3iVvuxF0eOnsCTH0L9Oua
dV9tdwsisyqHkIbBOmlWSpaEi8t9U2tysXx1jDWvvM3fTwe4r2dnbaR7lJsEtXUp
GnpqdRCjge8ObAMUKmye1/MQcRwklxVeZ1hr9UD7N76w8m0Qg9uuRa/3M9iEe+a6
OuYiaK4Kw2GkcLa7g+panOIOE1KNH2mNkBIJYHs5rZmecp3in5k2ndLRkQ9yr2p3
cq0uiPt1tRBUPEqth6vmeDqnLMgKADSoeR+NTooRMWaEQ0juJdmRyWyCeSdc+2NP
PgG5M8VaRlyBerUlSRqVJA1myzpthiylLQgDG8P72L8VmC0O9bt0Rvn70fXiS2/A
uWSwFglrORzI/Tw49nHNzs+WWtzy6rLYHw/9ZYGPpunzGCbAvWEQOvXcSYH+KsHn
K5LnGMks02I0i2x4O+SiWktEJVVTJayzKTQSjqa7/Dr2QbtdgF6RP4ST2PEkHTKa
AIinzJGCGBYtHIlcEGIAsF9Z4Inzs5pY9KD3v4r0OMS5uG2KUEXlt29bpAvXSXfv
ihz9zLC31p0eZYl2xbVrdkA2H0QOocNsBe+4BshRBZy9ity4oDaHRy2TJrGOlN61
`protect end_protected