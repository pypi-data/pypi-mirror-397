`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
GaB3xyH8WqmaCdxZX/nkcSyRvaPVC1hBwb3hp+YHHfa6cgS2h5YOemSdX8mL4aWU
VNHLNSguqYgz8A2fTubOFl5LM3oaCHpJTDjrS8f4Z9L6ZiaSz+QPg4wlsZOn8d4c
yxcImpkngYjupYFjIZ3wbF1MbWhGPw1ooOsORTAAdfMw59I9nd2RmhrWLivQ9Fmq
xTkpPyoLwk9MSqVMGsJYS6pA0iKHEQDpMTJiLJHf/Ii7GWIxU/Qo7HkmWT6nP9T8
TEfb6fpzryyzxDX4ybXUsuPJrghLblJcLEJcjQ8+0RG61eb6af9yg1GgH7kWijUB
1yK+plmpKBxDH4xAywNJrvuqS8K++I+2irhtXG9NAi9YOZElkzT+Su1veMzueAMG
JSzqAjVYyzqeivo4SP/rxoiYXkau6ZMMIrfSMyJddXV0GILslcfK2AZPG7tBTuo8
xdW4WxS2BPqmP4J47qOn97QxHS1YI1eDGEDwUQ5xttr6tZj4/2LHKLdAG1s/NkqE
gqP3VkAg+MNID07FduVfOpR51l6nPr72LXbtDiskNSt37qRv4dl23AfE1UK+Tofk
foYmPp8w1uP/PHb0b6KW0kY5mZAiu/mlmGHpfaMr6lVOIgYgdkFUb5CArvf/+F8J
KZE8KKDqDev5tj7fTjcq3W7nuzDhKX4zvnOX8gS26NzEjhcdOPVhc9ZDV8+pmn8u
R3iYnTBU4EBLDHKEQIiZfEyQJcX6ZF7O6ZY8nc2t5E1X8dRuQBhH6zyRtDwntsJW
+EhNUd53Wqw+YeveaKFk2bTSTMZEbtSEP9QyXBUrikUp7IvedImEOfGwHsX08QYR
jOPRUkioEEdbmKhNeckUmHK3M1Ikv8HA2Vfwp0zxQL02RP0y5C+qUBCjrkr2L7Gz
fVNPWrH8Az1pqOLFZiyRNIaZkvsbjbMbbKvLZxK+AcdQWqy5dcC5qgFCWkVHkOwG
jTwlLTo62fnO2S9Fi1/uhdVvbkMR7I7OBCQuiF6twAVTEGsfgHLhpIs0NvrkuncV
2aUO60al/EqLCUVzAzPEV9diZupPfRrnvkKVIle9F6DA7ObJP7DzmWMmikQGjBI2
sPgcru7nzavpuRYTyxNAEeMaZMiQHEscoYDpRaqIj+lWyq7a6mdYenyV0jl+3hRl
HdtlvFXaZmTFrID+jqNzW4AyANzi1cEaVWCzCgbAEpiMCTruQZdJAo3jc72sxJ9Y
83PUvJW+zdM5+C4ZjvXlj3cj3Bn5BOY3hrUURa9mTqKJf4OqcwUcUtfunz1A53q/
m2QSi4JKgY5qOV+tN2Uo2nU5evS/r7EFSA9OjAs4KTxlGfawM4S7lA9m7PLqBoBV
VEMss79Q6jjnb3cIjvqaEKjW0SFHxOylfhYdddtehbIltv8tlfl9MilhyZSMPjEk
WYpuEZ75h9iSXWRwDDOKxi1LvgA9pQeD1yC7usxwYF+WQGgMJcbJDrmR16WvUk48
65GpyCK+cpr7QOJt8XiPLe3YMGqjXLvowj8AgO3IMrNxfJMbF8dyz2obwPatnTdw
HeAakWMxzI5/M9En4Kd5KU7X2YQjq3btRDZbQZNTFW+yjNmM6T1bO9pWrM2xIAo2
bWzTugzyaG2hYnPZpJoTjwZXtaf53WmSPwKfh8d+jcIQX2m+oDxnZMGIE1WtrAsi
ijDyCown+FSmHcpRZikpAq6pfZWFJJ5LY/i8SW1ibXppFZNKFgylMka2/4IhTV0x
acZOUXeCk77dWT1THJ0cBPm4ONv2NMmHfCny/4v5PVYAtTcQDdb3YE/BHc4Msoc+
G/WvDcnx2DUe9RxNuWjojlQCZNqj72TUT8ZMnTgl5CRvpvzhiEC0qCylqdyEkDRu
73NkMQjLBX7165w71MaErqnlarKYb/tD11aYPmIXDr9cLhZ8TIiNqSLJR36cB9pp
SLlnLlvWRTwk/tNY6V9sauX4BGW7i5537xffSlZVRf8PXwUzbBxG1+aFmXNxWoxQ
L5hm9RL3h751bVmwhWb6e8j0PGGBZRe7WH5mDMyqg/K1ZHhEKcoLrVLkuQDynF2x
B6uCjabWKJGEupqEvDzplGqn+IWDj8pI2MkBDMCli8yLpmntX3LaM7ACDbndHKD7
HZaf4LrkoTmzqjOA+987lmbsIhYDMv50tzUFUwh/fvBhpkmDtX81dt/uSdui/kMK
VnaYcc4bG1pPIjhwahnSfRVxcuHOuA7WPerI+DmOpm3U4W78L71a/CWjLPrEKC90
H+JKFWSVcILocOLM3hQD7Ox1VzUU3Pq92vifZA7tVDjEh5omJPzv+mUvyqO1ziSg
Lhhz380qkwyt8xns8Q2Tpx4+0OSuXIOlCZhZoEq4GSx1NG6G+yOxnXbG+Qb/ifPO
1N1ZtcJu7vt3Rcd0+jZJCmUPikRFQW6anWtqTTmrdUXysyOde4USY5SDIEb8LMUs
aeo/c2+6N7EUW1xHI5wRSbvtMqkgFAP5QldhXfxVBBS27AcyfD2z6EYXwN7KONOb
oHwS2PVPMEXFvaZm2pXfDs2Dx91UPG2a58YnmzJU6xog96ekOzO/poi4DtaY2EcX
Z9C+heiz0U41l6l5l1y/Re21l3hHwzh8lncv3B80aJJQbA2NO6HuZM8rNn4KJvkU
XkJAnU8P4VO4ZUPeaUYU8yzgRFY/x3vv7lkKKR5s6XPOpI1sYfhVGPd/RkMkylpj
Lmijd0co6bgoY8sHOF9vAWMHoh44CMkn+CNOmstAdS/zdGLVIwSUZxFVftFkMlRb
CsVEkV3YU+29YZ09sYIZEzX3g1UQzr10aYY7A0aL6OrmbIDOPUO4V13I3IqxOgcY
BXiu628u91+5SZDIXlPHSMX2BFANLDZOCOY2Dbbla77p5neU2z6R+QxMOAc3BTlW
1MCB6BscCL0qb3HBKwmIaCb620Pf+vcRwfI2SxyGDQrtUBA1zPFf7r6iXPCiQgRb
s03LGwhsvuKrdWh4CXTMSQiUK27iAR+APKC3Q9wmjGY/bN5MomLMBgheLT7s2eb4
D5jN9r8c11C3QrHXVjtXpj8X4Xa0BqTZcYknyn1ISGQlZQ/WcyiuVfVmz5muJmkx
BkAHdbWr+dpsXYbTa1LPTd3uQSco5jP1G5qePvySHckZ7pRZAk9vKHS0BPzXH4Vk
Hj8GDkjK1Q3JdOozR9KUhmATDusvhIYqZaSj4eiwNgpENzym3OvIqIrnYo6I6cKn
4LyikEJJw8FDHw2V0Dc4hfgL1Hi3lWoyVVkDeeEOvHmo5f5zMvMAYJmA7lo75NsV
2uYkdUiOxpQe00feXwyNDvu6HSSdRfXzkVd4QJZeDhjXOqky7/Sbg3EacLEvTmwY
LmEgtud0EcwBcE+r7P0hZYzoZXhtxAVoi/uauY1z87Q/4UnN4szAyidTgpJq2ST4
dYJbbiAjOduH3expHmEzaWAY/Az413rgHjOJe29CAjEh6xchp2qVafwru+iSDytV
q8gpPGE4gtj1mxrgfYfzfR8EVIvvepTKQsmVgsDVdLMGblsWWg52IEe6AEd2689h
HJAXaLZyAPgFgF0FjpwhY/ttOQ0OTaGfvJaamvwh5B5CUMgk9IJwGev5Y7Z0G5iu
L0QIdZ/FIqDopf7cIBgJKdkSBds3PJiFnCjiFkxEH+pt8lLut31rcgnNwoM5w/Pm
m9obOsndWzOXaDKajrWqa/54PxRv6V88B0lpKikkUbmDJHvX6HNJW23DRIgICEom
xvwNp+KAbi0C2I35PGDfqPkCP+ezHGBo47zLg/0Hp6D8jYrwL8P/nQWVDL1nDhqx
2jkvPNsQUcXuxbb+PYZnp9B46NbeTXCMQolYFdxpDZjwVIo47MwZaPNSaj7S7I3M
hkjetOwNp5jPHN5LdTw2aE5uFvzROv6i2e/kR6jd59upVOUlEPkQgGZ3TIHdpCWj
KInw9x4T3eZGC6YKATu4jrrkAo0cYzpzG2aLV6cUjU6aLa8FI0scXvnUo94KJioC
X/cyXJIIc/NAR4AUQ2mudJWCSpjM5mkAcH6C98vnXsD4fY53c51fprHMwnKu/++H
fotZFHCSXw3ktKx5VR5vk0tlUo5pYzd3ZjZxmx6yqUq6pClN0E34EQsQ9pBDPyQi
yqiyTnjJqciGEscnNZuA4jDDij0lZJOy85pSbvgHnlY0xzUN3UQSn6/iQVKeoHc0
dzxEnNGRw4wgGC18oG/iNNvewLEYInkUxY5swWXYztHkya5+ZmRv8PTQqOQsOuWr
7Fj0T69OMijTB/U9UoMKGORno1S1GrfMaAHaqijW714k4eBkwpVTHUvObH99cuXm
AppdYglfeCxacDLOpMOYoMO3jDB+gedQcH7PduvEMovDirGjd3g5+LN2QLwsru6A
Y0vP2MTUSLoigUSEFyXrAwmF7RytjQ1czcCGHlSIIvddujim9RmwyaSq/E4Fv4GC
QojvBqN4z/a7ZBoqY/EJLIlH9/edl8rOHlehKPBoDD0ArQu3Ez8R+r2J9NG0wJsQ
9+kvPwPxPhnYx5aIuoLkjb+bcGGmm5RJGrM6LT0Upe819NmHpd7GlbrWaNCRzo1a
gaHFwI7zV4I+mKwjYAWw0H4pXobLi4GJRE1fXkELGaDxuIl4a6m2XqG9NO0orfxp
+FaNpXLO6wgtAhW4g7WQcRY73nCHm1lIAd1EcLivUmkgPiz9KzhUuNVnwUdhUE7l
wa+G9o3JdcW6PwAXMbr1Gqjswprn90+zaIJ53HjeXVjPz5Hgorl2SuyPrYzAn2Be
g57P5AoedTzU2taHOwSx4zi8T8COiXct61oM/kaU4fxc7PeZvhQoWcKwNYcFyK3y
+YBpzvb0nhaGRYJ7V4qcqvtZHRXZ93q3dNaaPoefJE1m0dZ6wkrYf8hq2AJIeR5w
+DIV0wfnbBvJO8Y1anT+9Gam9G1+NbUZkYgDo/Yw5DNe8A45eg8Z6/NJu0cwLQDb
JkdruHxxgHwrw/5wlQ5b490KyMPOKvkUhZAqxIpe65BneR9UvczeNEoCWSZRn1Nl
AHw7Uf+dlg4kyWuipZgHIgCx5LTVZegJ08khcu2nFNZhZAUnA/9VaAQty/9k/Ns0
/zhssrkR08yPMfn0IeCKikIr/ayH1ilqljyEIZwruMkSmEif+7tGMDCxC6+Ti0G9
1e36dX8NEASkjNFgYvkEMurY7sKQxPIzDJZXW2dazvzZBpGycx11lR+ef4G+4GOR
pTNFNOgHO91K3ejxTS4lKCCe9fmrNd7WfvYiCNDHFZ1hohBP0KXH0oUHJ2xW18xE
Z0GwdwB9BgHGG0wcwDOLIxfxls9D74O98154GhXsr02AFC0DbDYXzUf1Z/Y0zapz
GVNzBmD3kLwX5BN2ItB7P781b1PfpFJyX/DE9J7YdP8hUY0f28o+fGt2OpvdnoyQ
APsfSJVpZOwk7vGmKSZ/Ckud+z5TkKSnmVaTIocrEEiT4V6crcbTfaskC7nYMvQa
L4wvym9QeMjguze0nvK5I8/1NfWcZNTHRC41a3paHA9NQJJ26aKAe5U9UAuZYFRL
j/pOQ5qMptpT01pyLaVqtIxhPNH2AckZ69S6qJE7ycuF7qgE5K0Fj5tvfJA2is1m
Cb37+S2j3OLAGDBObb8473GRVGNWsEGPVB0IcJEi+agve2AcNsRWtIEJMvJvNpuP
MyCMJbnYsidLXfstwSIZ1dcxNojnNdFx0tXRNjciVt/ALpVNPjdwj1WzDINGpt/g
O6sO07/B/FBUbwU+cUMqE39bBF5qFH+lpt4H0QCfF83QF2mVsfU5X+8aDoSQfjOh
9n4CsTc+udVroVxDaWyHONRSRgv4PofGUI0AMtgBmYN3z40PwPndZW04FIxtrQMM
V3lPfhY0rYodxNyUrmrVVBAu6OwRVOQuYvO1nijXeqECELifConVbr7VEww7Fx1N
XZyc0SKnRNLtuCFQIiunbvRpZE4mKKH19XAo9XfdnuLUdTjL1BlJIlEJH6YlRuor
AmFdr5D08TVVosWIm+cbrqPG4nRijECOAhqcQySIaJ56zaTAVxmtjFEsPqAPGqSG
JLqXWOKkF+/BnBChJ5JGmj3pWqMLR0kzvUwHp1Wyk9AGmedhCg7PA2hkHXif7NTy
3bL6dP+PCAsNJaqEkeVpJ7KATdttFjgJ9rVUaT4nezRIUAXO3HM23AisJBMwk37B
hSWa9JNgDqmRy+0zCGaQNKil6WuNPu/IdTdw6coYSgruZa0SxWPt9zTwnQtFzYPN
dZGOlHhGzaty79A/Ybi/lF7UhevhTFXK+ySfHVW9lhBfCVSiNFebT4W6ibjVdaIm
1u2yhC5d2qNWHzi95HoGDb8YL29yUFHZhiiMMyDa1zOt5fvShej6PZzBz9r/uRH0
I2+HgiQX08enStsVSiQxX6lzpufZeab8z8EgrXtCNsjWe9kLz6PMSUe3OMgngmnP
AMlimj276OdT6R90Dvtx0y4ChcQFGZll/EcvaQXAdMHFecw9b0et2n3FCLdk9ksh
+J5JOtEgdpICpx0LowH4sKsnurKJAeHK/XkdmfppGv6XcS2HVPb+SaBXmfLBvPpl
Rp9r7RU3YzhagMfXnfRmLjHilE/5H/Fg5YH6dJE0SaQzkrBeR1dMcNCnwGqHrowP
/csoV0BL5B26aKLHcT3wFtiWXmf0QHvdFIMKGJQIEXPB5IcpMNUfvZhmhV8r5FnY
rQGL31LIeqkHoVFW1FdBwxPE1mpsmrw/ZrdauSj7oQ7Po5tR/jiVrmS7Aa/zfkgY
902bPo0A8qUalqWkucTw3EWfWG3IfH80471w6lcGUfXAi8WVy1sQFz7l3RZ6PImB
J0zzW1L9he+FdQ+qxGPnBqhTmgbXH2c/XsXBqyTX/o1UbDtpbWwg4tqA/j3+w4CQ
kwUI1yd1nxWZbkiK3cUMD6bxAKaykzcF4CsMksE0zFexl5BP4wQ8pJjUUwDFthXq
vBpRLScjWnVJTea/c5MCsDHGrhoucT//ez2EfZDlCB37cxwpY4n+ehyDC8LVLLaH
VcQTtxGWWkXMszd1zvhGNA4b5tFcN3VO1UDyFuX+G6oc4dy2ttEt6/i35IAWpQ3u
ohqrhYAPz426aGv+H+9IXlPDK0SvXPLfomGjkc+aBrtDxIM1PMp3kPy/w5/SiQc7
Xr1dG+XzqqsENDGbXYta7vS0vclJb2LSoP3uIkwOHhbnHnrgzT+WcgHmt1flhFyM
OdMSH4pR2svLO9Q9K5LuCWtJ3fcALbQkbz+bVN8sVTlGNWMhksHwmcp4ja6l/MgW
u4uGYhaQpq6V5XpZtkZ6mPYlRs6WY5hQivEFNb+8FK9O6Pl1aTADOUasAvZj323V
wmZRtDR6EzGsDzjCnsXj2b/n52iGvzQ//iNVfLxQHYnHKa7yPT6DVR12FFkOyAX7
YADpSI7my1QzYGcMQ2Hi+KgC74otWv7IfQ40M7PNKvuN5zgoDI/6XGhtKzw076Qg
gfJQq7KeTCazwWTIFlGG95LwXk3zY+zzxtIIunpQssrTghoQgejPIrCq+B/C3sdn
uZT7ScdyBbOe/0P+eFQWn5MIBIOHAJ418hXoCMTGJNoZVBSz/bQoahh/lUPrtHrn
oXycEke0LfWjWkd7t1ZtmCX95mehyX7IWyrU5HVzXgjHkx8f9KjbDB+mQZBAq+wR
mIaVZYovgIyjP3gtBU1r5bhdhLjqlqwZvrmHj3xUwsRptpcrVi4DEvpkUmHWUaM0
ea5NzIKcT3vdoeboT+nTsZWEXU/945lppSICZRwGXovmwFrsJf2sWbHd9Gt50dFl
+dg1jdpJpp4yBQrmGgL+edsrvsfB4xh8O6+4ngZpf/AIchBEVP5VHSU3fWfio66Y
xDDWaJmluVU0/YXW7bBlvS/aFU4uqWgh0b0Y2BjmqZeMXYLqmzlG3lIET1wlXDxE
2mOUEisYf71FIUC01zn6tJrRdYl/AidVXKo0ySQlMCxeJu/Ae03aSyVCoiwUZjSs
`protect end_protected