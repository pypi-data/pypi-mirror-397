`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzboRxSb1dtdRzfByyVgSOcX5DXpobi3CMlH33ga4f9jI
sJTleFe+iUUMVtSZDgQSbZn3QwGX0tN/9PcB8suuEkqR79201pUkzSmygd+fX0V5
HmPTT97eImlLAqMRe4gVvW+y7mkgBseK7GtbmQV+IKAMIbYpT11NdKXiHNgN6+QF
yHSGuI/X/44+OvtE5Fk91oxiuP0OYyZeUsIbaXo7TEaB1NBLXP49NsE1rciXtJAS
3vcJnnMCgOellb9y31SO0yIr18uKRS05ktJtgIw6V0TY29GIfdoFCUAFeDYY2JFd
hraHgk5ax54EGiEdboiZum5pgI2zsteHoguq7pAczjGAiYbdeYTLmb3863MwP1O/
Cnl0t/o61EeIlpUDIdbFHQbRU4BphMoV9ImOQGFNhnzSQVgdHDeZGwHYL95ZbhwV
zDE2VgdcJ1eeCBsH2kebjYtFNfAXHl7tP/phzJqKogUs8pEg5F17KR/+/kYcVZ3Y
rT1a13gyC1UuF1tXzRa0smUDpDm4nV3ZUR+nfmEJns76FNJ/NUVTp0q1IJKUWbJu
AiZtfiuLyPgXKqw8blygK2SO88wY0oFOq4yKSW54d5pMriievg/c9sp9eQy58d7i
nibZkJFeH5UmxsIzr5zfYaFDobogZbAJYnh2M5gsmcijQpZWcU+r9lzni67KLrHS
8TlboZgrqlvJ2f/LihWcsO5Gh/1RldJFxlmEc0pSiCWVTlVZ0WgNbIjy2uxGgK+P
nk81cJ4vxUqLAMPfjGqleZ7TF6Mfoxi621/rMJT9xkqx3MCamMfyTF2+PWxzKSH2
s+ItlaqOxQz9qzR+kLsZKtKOhvSaN9ULjStZKTT6ZEWw6/CEhkNNXboNGBmI6s8R
F4w/sN9Xr53J/ii752KyJrdCKHE/DK8KrOuvk6uZtcsCkzFrBcLw9BoptP34rdGl
phxO46BHWuMqaqKM/5cFh/ocSHfFvbdyb3sdWOX2AYVcpPTHVlUY3ETm2eJb80J1
QGoPxyzbvze25KEfOykLpZjLeoUeVQ9B662nQ9Xy0161Bl5PJoefPyRPQ8OP4esr
HvY5TT/D0/YIO7zCvuiZOuL5yCGngahr9+P8DQxIqvrNFHCPJWQ3HpprEKRhHNHH
aCj9f8wUUfgccFHyzohBvPzAEbnv3X7d69lX0j4Aqgo6srccgiNdrekQ6Cz+flXK
0+UFHPbvkkLkNoZzurJ690eSycQw/oKN3RSGHcfqCPaJw2hQF0tFgsyM8fOzXLYZ
4jiw5NXQRaaq3Gj8khN/XoirOEmos3zI6bLDUb0qL7N8Ef2x6Q/ZEOec0RJO2Idn
DykKBs7LnWlzbomD/XHDXZph2Uwsx6brQ26j6GoK9wyYHP7oLhHuyUHWRhY4rR2f
Uoea5VzYgC7wyWjXm7rQz5G1nL7ZgogEy2qFzoJjmjLuz3wuYpHJMd0/FNHKFu70
72eAQpr8yk+1mi5S+AHF+TQ8KwXeybwfXJp7Q4dCj9Hh22LzLtjjXNtnI65QayJu
or2IhkdRivYkjIq4DnIt5kwXHrsuCwLBwk+PaakHI8sa535oKnP+VQVuByc0fIP2
SUmAZ/z53dGuKynHVaoFr5uoZ1JN7UGlHd+1ZZZJPAci2vVk1BPQmiJhj9VdB332
YrBayTP5c0rlANJ2I92vnU/jqEMlpkiPGa13HAeHTQ+TA1ZIHvzXn+3RKCV238ez
zLKFFsP01SoPQ47uYV55Udb8PwGL9IH6UmKh1at+TmGH2mD8O4CdE6zguyVupoP9
ehFGWV8imSa2GfA2TVb3fiqiZ0F4ECpINLv5fvOfuSsnmAZkm4WA6RFohTOpkbnF
bSsAH9aAK/X5yWpjNt1oaCzDxw6I75bdJFBDG5Gj1BxANihshYz+iASkCN8dd0X+
b7d+aEaeKe/IXEQHtgM6i0BWo76SdnIXwM6maAC14CbaEm1Lx0XhmXfVk1Qb9Uj7
ripv/85gQnN3OqudRvzr8s3iTrXi2dRfW/902zu3tFllBTQMJJ3Zq3Kr2wJdn5Ot
9jeHcjUUj/3/hWJqODvUedV1n1Ekh1CrsmjnFRnXYGqSuAq7F0c0HCth1O/hKT6y
L68BQIVqvUJIbuJ4gdahQ+HA50mOcNyNjW5CamuqbKKKF3BRsdpqeZh4citsMQzJ
IqnHD9TmUwPjVh6SvDT58Y+BtZSL0gB8tfB8/LCUPDBQnWwoKB/42ssHdG+T6D4y
ZbqN8Fm+W3ztmQuvtgf8FWA9egSUAVOnMprGoc3h/K6MyVhIggfmTNBdiK+l+vw1
o07KiDTjSv9NWZp5EZWxWZakhADscaVBLdZzR7SGwVFk2UjsksNB5fLSZGHpXeqo
shVkKgVFwULZaoD9CvTQJzxlZ7EdbYkb7dgVUqRI2ZfvsF94paE7Lw/5nJ/xJzI5
K83GfiVBB1g/L9xJVcoP45VmMb+CFzn0qPG4VY7UKREjt+g/BvUsHYzOcxngloL5
1ePcPygdYphSJsM+sQb7EEc4bQ3nMnxdE3fjA4SLhklsWUjI9d0mBtk+1kjy2oIm
k6QfVKa3IP0JNWF8Qs+sHyWPnC/9iNud2y59vo8StQrVKs4/Ndwhp+jcf2vqb9Ti
OgURfDNeqe4OkgXJgOFMYa3B/uPPFCEv+HzypmbZ/CC8as3aGwohRf2H/vfSe7gg
Lk5zMFt4e9XdWl2PoMGTF656YYecO6WUMfIRPOfukOo2eq5uIMPKMzLc6CThnX7w
lFgpmfd0XG4te9Tl7QTNr/NuW+HRGFAb5I+Ws0o2f5GhDTI+3awSdUwpMUFP/DOp
o+3UAC5tsOzgsfPAIE3+2dmcrupxFaKRoEzzVumRlS0II10ramZ0LiSos5p758rU
aG5adagG6YFVjlbr9JfjnuMvFhmTGBsp+YY6rB493U1uA6SphLWu4TpnccuOwAVZ
SYc4PNReHwdEVAGGbLBJ9Uk2jZkE1iADATATzDPA6nNIXxQyhP67YPW/y7jl0vQ+
bigkwbXTh2wcFC7DA+7tcwTf4/5Fud+MLBYUYEIkqYR6FIpfcOwyXSOUliTELOCM
fxw24nnhhT81anZLN5j289m058cahgxbclDy0m8XFGjg/6vxXof7Tg/fgIN+4F43
YOXzPYhCHdx+de7uRt0enassHEAtbAEGM3igvXLdyOt8WANICHe4tIsdd2GTzF7k
nYfWc9/M4tD4EpmwarBzqFWTIS9OsXilEz/9omWCj4NMZIWAtPLhZvGCfFlfVbC5
DjQxY3rIvxDNldNCNnthNoSaIhLY/iy8HX1XJLpjJSafKHebZ4bH2IWzoPRPU8UG
VdNB8BLoABqVblmH0TRiB4kgY84QgGlm0sO6LYXxQnlHeqr6CvKLhPp8bn3CjEk8
BVfr9e7l6vmsddCXEGpSj3S7VJM2XuyZPeMZOIn06GSBXLAGyAaRdQQIpcD8FS3R
kYPaEko3JalHzxdB6tA/KNJSGN01OD2dhharMpJDj/g+Zbbm64Pu346ttusSjrGa
NQImgbF5hVh7NPjBDXQUN1H2H++G5bjecWGOdlu6LVExaZueT8JivcaK6kp6kjvD
ziYL2zPj7I5cNDtEpU9aqR1nV52Zn2C9c9fa00/uY+m5/ETcQYEpfFjUQiquAmoU
9O8s0KJDzqBcY6KQNoKAET7VRjkxPTKevb5rXO+Sy4TwkFzI1Aw4s3fiQEmCGy71
oiEcaY6m9ePedPGKD7qr1P3ilb0CgUYNyw/LqIhw4EbTOo8ZjIzW5IlRGCvkpZ1+
m3RGepSTcGRkY906QtvK6gFinN5ZgiwJkC4ZjKGCZhXiP5iiKzhFo3t6+XCRfqDI
5LbcLYzGZMGhijqmyTVd5dqKM6whsf6LIAfIfVdxFSAIy/UiqNTDqyBb5kSQtvVC
xTIcgB8SmCaf8OC5HZO4cWJqd9C5aDnBjMovcOikGs/x5RdpNed0HutHYzPrT++k
tCof8Od+An0nH5ns30jQi0B/zuadCbSKUFoQqKzjDIaSTnvdzaCQjQTk5yxy6MvF
7BqIlackFL2EIMdm8g9lDVm2sgqT+NgnA3W/b7gVXYENPt8OX04WdNDt39oKuw+I
A9gYHczEW5uqrzVUWxzjpYLE5dsXUgP5UVgLXHTPCnrB3I7oLCwPLLzhJXdckRRC
wuqDHWGt+ETeLwzxcwre3p/TaLCazXo4YxFe3olDbOsLQ4oayu2Z4mScQRz8KnmM
rm/HpA0UwIiWWjyjczf2ARkUc42UDd54Iz5FXnr4gTpPtGnZ+JY1QX+1wBxLKWHC
qg9tj8UMqOuAmF3iH99QaHLsAfpfjU/oShxBMCbpsjfsraJiHSUk9jDUIls94Gir
CDf8brcTG92W61jyVnUoLYVVERLWUI5BywoeBjTYqOC1NnS0qqUXOqORowyPe0qW
t5FXcqlpyX+9tvoezqyYU4E0sRLcaXwTtS/nkl7enMqCXEbU04BljiU/OEUG9AXN
V84o+9a0DsezwlLssGPWLnpHoZCKVijzWcl4ZOjCLUVaZVElIox6P4WvYH45r9RU
QiwtVzTWOoBCpvQ9Iu4yyxDITW6ibrdQiP4xXPQv3CTl73yHCyJVRUDGqRV6hUZN
1oWjsU9HLpbjI7N1Uc5rI2Q/Zv6WAbdhIHARwVriAkZvaZP2vQKvW140U3MdlHhE
cCfXh9+JyP4lOHRn5qSpj0xxqXbwdCCQh49/PNez6Z01wyLRg6pWhLar9a/w7tre
Qoy01HzHIWQZEqvDfHknhZxUMVuKkwzZ/m+ATGUMEvgXqhi1DR4VARBDovdSvPGX
TcHqpd9XSARzK19/CdRemyt3dzMhsEmQfJlhjCPPSt1yaELTaO9hykf8D4MKpSDJ
oO++mzhtaU0dAItjCdGfXaEZHGYMM8X1zN2glzGh2tL5uZ9N9L4rbyAZFg2NbZMQ
Tlzz6VWWM8aAUYU41jnjN+ni5ah42jraXVTH25UyBgxf1b62XvFTsPUAu/EQMLWc
WTk1DRnIVmg03vD27RBxu3Yn9ae5YSgGFkzViQvDuhGndUSn3jRxckA9vfOnl439
LEulSWPWTWz8nfoSqx0cY5qFNu4E65AO2r5qdgOQMbH1/mWi9lIu8R3IDQ3SqZGg
hyPCf98ljYhbt0sUkW+Cwydx0yEZDfx9gflBGpnfwzhGtl2qHtPTj8AeKodTe4IY
QR75XtFQj4DhK/8sIukaWmnckxIFmRJgan8D9BZhMWZ4wVnFcIqjHzKQZx8fq8pn
m6F3oAUIqv7EU0uA4RBAfeMTkpfdHFX4ai1xzPrksocnbdFBFz4giAggVoCFrCxM
ftMc/zkUxhlwSZWWA/iuJcxNbX8tr8gGMd74yNMue5PVz/51+zvJEBacA87b9FFq
C628upuoKGtwwip1bv2F2fMnaJzbZQjNgnIcsTJd1MFEY4DVEc5rx9fy6OvPmvRG
VEMDFxdgJ5o1VIAoBNRGE+esh+JIpV6IGtVenMInqq4Tlp1ax6g0vD8CK9MoRLoA
q3h1YizOjzSk4WGvDwXixRFUPqxDB2rsbM2s4m0JDUZR6iUKZma8/aDUtOsrZsJ0
3Sh6ZFN2xkj8kKls6sfpXjkI84GTqzEeVKu3exHvI102iA+QJjIWECZ4QFHbdkkG
0ROJwbIquIeqeL7cu9+tn8CmiOZGmbClLDVQn/BYZcfkPT5QxjMci59dTkM1jGId
TrJRSFA5J7FbcZnw400xGDXtBiOTKpi6So50kdgykI4burOwax+2HMVfMOS86hcj
bwt6SLInsNabHJe/drwZKjIawHqX2+A9Bn6vDeSXpYAP6+TuH8B1Y1TR598AHFgx
iuBspDzo946e9EQW8tDXO9ogentQqB90bFIJ9U3yWLI+C9KeGZ9RTsY6Yvci9DD0
tvdqeOxmjv1RzXbEz8jKMbzQKnhmtcseXKc8LGk/0n0bynWpyqSDf1QOq/n1FMBf
jygS1r6FLyr6hxLQY1KHSh49c2cdMk6s0H35MdACw8YRDYQ+tgmoBbhKQwSwloDs
ve9WwuRpSteYdsG7DiiL/k/xmAieKIQEzRvdeD2lmc0BliPIV1GUedxd562jEJUs
HVuCChWK2qWRAfK3U+gq6pGrIs0EYj211sXeB/R2pTlRQb1k/Z6okHkI3LxIMEU5
kynYwdjmLpLDipHuOtt7YS21jrXU/1I+XzOy7I+57S9gqeIxgSU7wQnr9cuNRckZ
WdvNUAvKfjc/Q0e4bEDO9WQR9KB3Qk+gji8RyPHVXfwoeoy5pSW71+VMoxMRms9p
zll8bcfo51hR0X7myfeP/HwkrWSSIVGH+D02w7uPQ+SR/yt8sguAL6dyfjSwb8lZ
WzIyU/HY7z/fFrV3M4cUgMfqcAKNgD42rfxC1jyb9Zqz2wsDXRJT9O613v6B2u6k
V4gad4Eo66m3VT/DwLmnu8vsjnSiS0LTmWVvpdKBcmTNNsvSKN2r8vBnH6+q+iUd
11w1rTwPVqv7BWYUF6XjGG0ONkq4TKBk46zfo5sGwFVoA5BHOtY5mJqHh2WwKl6P
rS254K1mmBTLdxcsd7c2iIxXCcvj4Rc8d2AV2uOIILbLmzJvJcdVHRGWNSLenxn0
75sZWy7nxcgB4OpXMbfPMtcTVF51OQX2Ditdi9xJkgjCVTvzZvM6S6tt3ZHvoRfB
lKsW8T97+WPf68EjVWindiAjj4p+tFBwyq5v5GSVisZ7Ng/ScfUlGqLn+i9KmYO9
BD/wKhVv/9m0vDTrPoXCz2ebJ6ZF+8BLP+hSrOxiOOGCAowN7OBSVgHL88hrT2gF
sBWPKaO9HY0oa3E1Zc8gv3ULWbeRgV955SjmLiEb4dT566eFE5VP9btoPOirVKYb
CAf7/X7FgtETVSVjMFJ9c5kMYpRJ9icjpNJhNf33RfncgyEWeKaW4nOUUnTPYPNd
Dmq/6m76lL4GjFkMbeT1Qd9hhwx7MpFokByFMDC8dHBzlGN/LbHInge+GSE4oRKj
jK0Usb7anIFQw3P661YmL/qGIU+v6TKCzpd9GGEvErPND2s4afDrYkvq+ANOuick
RYMGnEu02sOBb+UAxMkQtMDdlZqOjr6kwHdwjus+i3eoM0qlAAbu9Ni5FGmGjSMu
nVjoDITQvZg3YOgSkTGjFJkqCm61rpybvK9g1r+6DvMYgrzhbe8Mm4ArdCyLc5Z9
AB83XTEvarSnSYFokeYlTUQK3Lno9GfGYc5tltyIT9o0vTsu79iPocPMXuKdwMgw
oSLa3T1jgY4kwQqPGxBwWEcxd4MnX98zXnxNHSyRL3pbgSW7brDOj5koupu4fEnr
ZUOIQOA6fiGtWlkWndjEHmf10YbckCq1+tO/Fv/oTUoxm2v4hv6TlTKtCzmI+Lvg
3Z8xI5UbEauH/GDkxuiNRUVZwzOwUgqTlXWGj3MovjTfHPgHI3BaEP4KUIpg6hbt
CgV+IaokwiJI17kmzU2pWllBp05Ouzkg9nkSWXFv5UCXVGrAgwSnsdW0JmMqLPb/
chtCuI/87BSZ4DOcNeA3oDff74XeXLJM7iToJCLUjv123R0zsvogrsD8zmNOnuix
WH0GMacw4VkcRDX2Xm87GbKoRC7jSZJwr/RdPre70Kdclc1beA0q3U7eMPbD+62s
jNNxKBo98PBBVU2W3lgQrsfxn6nSa5GAVAdHAkYvm4UjZX9jX4ROKmwGKxwGWdOH
t+SWxvQREla/avr1CMXELJaHtQ87pLTblwGJ1Z32/ub+tcd3DFuXXS7vfdyJMwh5
IqxASa2c+dVLL2MPmd5zeAxEztEHpasI8vHmj5GuqmlwDH94nGGwnaKItcI7bmtE
X6lI5Wq4BT4Wfufn1ojlEsY2q78ZPqXmhhX36KL/D01M4ERvHYyW3nGHENOFjGD3
+/7Y/HlZS/0HCFEV/dpMi0y/b8gYNQhhPza0m16ENu/Fp0ccrE6kRAakDjPtZpQ4
clA3exXaad4kaDpfg8tCT6p+QaAOropRZhPLo6mtiGHJTQgtgP1Sku1siy/NUADm
bLmBKpzmt6H5FQzOCvDd26gWW+xsIW37XSwbOrapk50Jwm/r146LipmV4q6aSyXr
iIgetfOLAQ9+NXQrX4d8wq2hDX9svsodiaY0Wo959qUgrJ7LjJBbKPXLDjvoC9RG
CrtSDjw7lO/t8W947ShK8jWV37Xh1yFvwaPL1UhlgzctsVNdbZcFo5uTdNk1RdcS
Vjf+hpojJvl19VtKjnKlaEwQuVrUDw9K2+MmU2piYqZDylzduF9K3C2BrbXLmYny
pK2kviNcMWchNSw4Ats0mLJ2Qz0leVxOrJlvDTJFGC87WdSUQpcvcHz3HjKPFB5K
n8v/iTI02Qp+eVboqIXPL5gND98z4MqGVT13KT2ETChgXz2qw6+2m21S+wr8+ZPr
0Fs0K2u9pcVorU1kFRIGMF8KSqqGl6x8w9G2pgY7XP7V+zwNib5iyQwlcrLfhHY+
q0ErvSaMRxdbUTsWR6LvpfQrA/fjAV+/6rVFXdWkSlpby1fDM6l092hZHRa4jDqy
boCREG1K91ey81dEcR5a6GjddS9QXxhEC3CidX+249a7BM+a+L9ApwRLakp93HAw
9GRUGwcNTL1ylpshbl/0ReM8TZSbtK8ctuuCSQBpOqzXKYk79vkZOhMCmepCo1aR
i4HulCIMLJe5PpTb3bIlTVDOF/K85oSrRaTaevNo4M1ilLj7FWwBZhbguaycpPLR
8uxTSwlIZ8uBKAoibti0mYn10zTuZA2ayAIpXQcCr6NV7IZAMmIXIgJJo4f3XQLh
D9MAi44JJkoTiAtn3/AjTRzQs0TzGcV0cvtxzdVguVCNL0wSVwW5rUPab96gmfSv
5ZVlt70BGEUYaV0RLYBbHppyH8BiqSuLekoPe8vKuElsoUODQZsf+MioiN+jfILO
XUQxOvuaVt7YDj9YRcvUN0ixfu6cul8deQT6a11OqRQZ0YXv0ikj4ce2ilS5HdS3
Prj822AlsmcsyN2f8PbMKiqnIImE0K6F/s99abRfaOEERHrVMTo7mJOMBEgfFAd3
yZO8qSByxoCRKVHbxHz+hhHs6Nh7nGCeN/eT/tKFmHyPWN91QuOFiyvB95AYk51n
cZBpCDsPLzEPk7tEe8inM1aAq/fQn5ekmH0YjCqS600uD8OiOME3iOfOiWkmkNLi
9lRlgH2hU6Xf/VtKqMMpMC6OJewXFTSpET/nZ/vJ2UQNrqZagZ57N7cSpqHx5Qg4
uan8v05QtE0OpmyLkF5ufVr1yBAwDSVmB2HRLnIuTa1V4Xlym3zj5538MwGLsohA
87ZEhXzhRwtnpG5K/wtM8pJHdfOmx7yMZiF5KpU7fOVIpg4BvhQRoXGzBSVj61Om
v2d5JZUjyugLxFTF+qlH6Pdidtmwp6eFC+KocI8nTKYoIm6xOQaS0/VPNhJ6kAvS
GF3lMSWr9vEdvy5L2sk+uaIfOI1gwpCtKQ0PpUS05SRoVwjrYVErbBJbnQ5kKOYn
nca6ufMnIVn1ovVYJIul1zhJF3Y0beDzjxINQj6jfKeb6vaVVaDuuuj7qmQ35F6f
GYgxo4/aq9DEZhuvnr0M5sV6HZaY+vrnY6ZJni4d1Tm//fA9tSC4/Vd70mngHY9U
h1f3fC3o4Ff7PhP53YX6nBMAtwhNaR+m0Sw+pVVIn26Bh5typSzBJwFgNwh9sJzQ
cdsya1I64BGN6ztiLCMNWd5sNbyy1DwTrWVQnHskfeUPgZwmkjxpSi2cV5kx+Of1
aEgR3TFMo7Opwlpvt170SswgurtmPYzFF2Ta9IlK5Gk0FfGVXDM5zUDspde2k/vc
Z3KpnaLrYi0p2NIBg8j5akRoGrEvLI+M9EUOECFoCcmENMWC3p+bXFww/Mbjqe0n
YrmWuj1EyA6AyXN24LnjzfK4egYtxL9nsmhxCnM0CnH8Xc8OBvJNoxUddN1sx9Ow
x2OWMmeWFEaEhQIPKc9i4IBeCHzYzaEqnfglcRDdNmpvEAGOsJ5crWwiXy+/Zt6W
XMhdvOk/FYyIiiDRZJs5+4rGh580RvCyMgRqu8OQSxRrKfh1M0x2zYE13LP1LBga
YfiorxDLgT0A1ZUHoXbC1j4dszN7zXncKJw/kaorajjIxoeFEY4gqI0VKLqjSqfQ
lRQ5ATRzzikPyikDPodJSSogaA32uq/MtjHsPkaBwqBYAnhYEvrxCOoxiwSQwP0s
TwrVCkbtGtqQYb+bYQDddqJMzC5WxlFB510xaSqMjT1GkWrCwOV+s6QL5MNp2zbp
73e7A3FpgYIPbGSNtNvJIJHU9+YnvgOLDUsNMRWj1D5tk9R9OZ41/0pzBd5Gl+TY
VZ755e6JR6h62xFyoRfLpzzj30ia2jnAIQ/6g+DGkN4N+RS1UyPrIzxKcyS3+Ic7
y1DYtwlW9dPoEglR6WJEQ4KMUrUl+tVddIpxLrjiEcz/Smv5Ubnn2117HYZtBrCz
r8tlE1IV2eY9AyHIRM+nl6G+uAUzK9k5YVeb6Fqwytn1F/LpT76sMO6RVz2+ZfBy
U8d0vhWAKz028iVO7Didp0+RQkoUWFvyeiP7iy1gO/i+p97k176YEt/ZALePkDUj
e2b6oeyaG7gmeyWtVAquBHPCKU3Dr5nsnlcDb+ALB+tNsxxkAGqVc2C/7G3OIVA0
REFEOKMsqifhM/CYC7INO+LaBoCm6Xy9GUXksNrst3WdPpSndI2sDhKtFCQB8qTc
JEHS89zKkPY+YAIaHaW2CzQE3mUOnwjhHX905wzozPKcjrcB2x5CFbTmY0vkyOsa
BgVatT9sGnl/jCh74BNDkeoabo6NLqhrKFELriAovesrMvjL+urbcMNmo5ZZDb+6
66pJ5ir8P/ytp0d07cd8n+OuUx8Zg8hBQsHAm3iGRHUVWJ6qUTIbkBA8YEkoqk3d
dJouu3pITy76u3hd/oxDTyaYpzMaTqIgUQ0iMSFIQn4t5hiPNQ6Jmq78LqtF+tOG
VMe94yF8a95j9YLRN3MX8NJqogaTTBDOvuMa61RrSdT3JMHNnOdCVZNAV79KY4NB
1WfJcV1viwiR5cb5pHskEVlXbKHU0qWsWGESv6ncr5GxZxZnmHnm//Hpq+ZumGtD
WCnslPDwBaON8FbOF7XtH6eYCoUzwhjc+uB8A5gKIkJzWKpms/wyqYvyy0ILvUjf
/aqGIKbV0ZP0LvRL1p3FCGDJmHU94EwK/q9v7o8/RE+/OqHlBW/zC0bNs0SYRfib
JjBy+16KZIhpOIHsF80Dgb+Am7S8oX+wBAoAnE1ZyC3pJOCS6hPbj4rMFMsh2/P2
+JEsFKcAJiYMsTZ44NAxJzEJYoe9T62iW56m3MPBLN+dDmydul5lPL1JddeSOvYT
1wI0MvJCOuo04kcOO7mkqXQlsYztYM4yh8skjm4gWDK+rcGL/RmEUkkLfcvcj8TQ
Ly2bCLWsogaou+nUEARY9Y29uhvJL+K8aa2/GJbOS+1WEkbxKDAOhkut9XtMu0Ng
X/p0LjwGbuBc+/Ij702kXPg2+IzG9P0hMh5YGnIv8ng4QIjkuDIHciQaBaM48+fz
AH6NMqLb9flLwmr9CxeIJ5X/mrlIExNe7zpJx69JoTXknU9vhBCVVXDdXcLapb0E
uQHmHwtvMa5ybolTpvHFMvTa83KmcQxl93cbL1zLAGmG5Qq3/naiIG6cHjALlhnM
BRTJpl03Sokv5wAS0ZyX34v4FurIb2uR5W2R6liWN9YA3Ts1+CnY79FvrSVhiNxo
dT7OEZyVh5R3JmLqPoZlUNWVEAUzo9kiCYDLso9ZTFXz4YgRdMxPJxgemQytAxXG
tHIhjfoNJT1fHrWZ5sOHf4iOpufKJIPJZ4W4u2CsVNitMm45YH3CijQ/UPY+qfLm
9kIHNnFt7e0C23insZqqijafxtaM3R2xxWmY84xalu70ghq9w0HNDgb+WQMeKpNb
z/N1B+dV/3UyNNAFtoNjxq/U7f2pvXKXYR8nPEaoEOuQ4lxiQf/XJnLlt9hxqDqe
6QnKNQJj7VCk4l2nOYFPgo1OctJgcXf4GVmacae2n1uI18P+u3HThYOYo4CMVhnp
ALmuFmIv7SPuECVhtsKeHaAYih5ZDsGPs7q82EtEEQOP2N3GCmST7RTm+FXn/n3g
VyUNFfiTQK2EtSY8XsbIQk4JXPna1ulrwdXuVR5uKQJwGE27C0gyXu9djqRdBA+C
PU5vghMRrd5Kje7uGa9JrCAFtWtNWvlPcpcXQvufr7jlYICooHLDjToLtGEwg7Gi
auLM73Z281/dQd5FPAF0WJCfPYqfi840K90NMeJRUdUfTvqN+AkjjMvUTdsy4APl
/an0DtbWzyfVbMT5CX7fZDXYNaY+4uG2HxwImT1KBVPUbAzdgA8qcWYqDhkXTwVe
Ixq7/2O1rcByeyYL6IQHHgh5aSfncYAhtGvhJZX0e9nXEbfuadAqvaJ5tmXqgEl+
wQY7XN/FL0n97yaAttVrCVAO8YgQQDectxboeGUlhyGkmZ2XJqG5MyFYUjhs2M+7
V5WHmr++vwMgXG7YNe7edzWrEAqX7Dewt2r0r00TWdK0p0HabO+jEv3ySL9ZD4MU
UT4uYEDrF3Knim36gAwRhwCOw20NJZH1NvPIIE85vXySS3xrkJHgwmZBUk8aQkeM
tSQiVbaXlYO7PSyblw7t8G3TF/tSps/KiX70Sf5ynth+ik0uEaxY3IcXtYxJt9zR
bUy5eRnP6XPKQoNJh4Qdmmffn49q+eBlxJpKntUC2/xJQys++jKpXrnTwx+cxA3N
43RImhQsqb8A166wJof/CXYPOb6e+viPKxwLHhDoX9uhJvTU6qXX9Hu7+ayqYdnj
r39F1ZV9kVNvDrtClTOrdvzS+2ulr+5xqDzmnwimVTY1fQi+HYwuS+YIB7gKnoZ6
gH6YFLkgcXtWFwD7S07ZiQ0JJCaJ/RtGullPosgOU2PUAOe/RoIA0VWAp4OzGums
sqpC4e+cEdFdgmd2Kh5MGQB0RWlOkRo0izva9pmUqZQPscS1SwpSH25s8KDpl54r
rkWBMVJeHrxSY4a1UYmp48C+SrSlxJ2SB3N+u2+KsoZ0II5tCfbOnJoSRwudixRA
4yAz1N1x5R6ht6oVXIO2NYYGe1UR7YONIOsisn1Fxd7gpFDyNe6yjpw5MrqA4ts0
tK4oboGIRffhiYgm+2ppbQ+iAuXc2pCmCoxwnuoyMJXyWB0Hdv9Ov7NyUllNpjlp
cfbPr47OujwJoklUc40JyAK9dd2GC7kjjgiSG7L5vlHoPJF56h+nl2lb1UZsuBgV
Wm0BrFXzIOr7CO4s642EO46KvnQodLe/00lVN4JmJldcM3FwWplbNLR7ZV0X5nkY
efjWbE4IrXxW7QaKopI9dVtW7yIcpGEGzweIuEYYOGXxOtivlskbbS94zEnLhp3v
3SCcIMd6jN4N5/IYbJ5NJjjcfttfGTVGy7qLvfMNwgVShtIaYYkll2u1vQza0sLq
MRG2OAVo9RzK1W/am0tw+LIMOTU/GRM+y+wEILx3LiuS8LeYkLC8vlbOuvp/GDLw
yhfqNGz+lUVLZQYEZTb9TkqzdcLxaIhaEn2AZA34RDLnYmZmJmjE9SecY1OlJ01t
WMnROez1WY7f95VCnb21liN1gqi+/YOLJDAoIWCtl+EHuS1P0vBw3JHPgeYnPR85
6GpTwIlpAKey5DkUZ2+dsqJhNksSRp1UvRYi62RMpQiBF/OEzpDYUkCuiMnKVnLa
Ftbv26/s1LmpNqvuXnJGMKGbNE/7REvFOw5sMFlqKjOoaABncqH9M7gvjd78mcOL
i2kOdJhcHZH4vvzbWTnX2MKRzN50pKKXJL92VhMX5aB7jmR3Mx5SlDQVbFpLjLgo
mivSM9hNLJLjTuKeBaNVWoI9KyBqdng1toXEWUu5898cm+Cb42ejztNE7mIqPDGA
O8l/o6yd4bjseoz1AzjFNjMftyVnwCmLtUIYyctsTtn+7Gk+pZ8SsvLvhYtKx/Qy
gD6dW/Au9oPdJu1ohqRPa8XDEdnGlGirn6fkwCcKzn4DTlDZUiwvh0yZnVPpKxL5
YCTbGjIOuHaydgQE2o1iFPT3V52LlVYQnNJUroEPN4phss8EeJ7xWgyOo/WlZXY8
AoXDfDATU4jLQuTHv+/TcnbMgeDmBmvJW0I14UTSSIr4tbFmNVRc51AESxniixyH
yWO98EqHBx7OUADSbEFqFm8iAUlKKzEHs/fkJSyf5BZfnZQz8m7Z2ip8T+NAANIq
jOcYM6dAdeGsWfVIq9/PyNzOPBgsVbwayAKasv8nB2HVrXhCGxpwQGsMiUN5+SEw
CAnhUUKrMEeNqxl9NCw86/cDRFNggk3JXic1hBhNoiGuFovAyrk5xAPleglIkC1B
39u/tMIG8aWHZWpfjv4txqzaBfDwe9/2xO0hyyFo+vh6pBmkJj84iVWCRnYcQbDt
nfPCJo32wsfIyIiFQa0cGUPPu8TPjvHBc+UbKuyIau0ysL5ujf6hjtxPaiajlmxc
fYf2vlNL1v08dr8Xg/hBASYh245ySWqCs69sHgno+z5tWrcGAt7zOFPP5jQxZgKX
scV0AEsRZKx6QOxvCXrHnNV0PK2Nc+Gqc0M1Wam8yAzFfqHTTxGd/3FFB9wWhbyL
99Lp45SNw1c/WssxM8e8R5w4bCu2BlPxnkQfuhQTqjICxzuUoGdorvOF9aBQOgMu
eBxzgiFlBw9MpbOPMsWTjiwBWKYM/MXkvWjrgVa0gXP6cnr2/aPnb6po35plNmvK
ekjaBvZ5aKcbB4NsKxGocuZy47Wd0HUadeZsL6KqTQ04UTre84stGdE4nEX9K6I/
bmnLq67D4VbTybrk7o5OcW4L6sha6CmJsX+6IvCP9ipXJydMgW6S2D5K5F0hjjXP
pi9gxd8sZi+wklse0lRP+II/jFnNQKVM2PVZUIXqqC3yMHZrwqg8DLvYs9gMdlpE
dbDv3Qqhf/p4s01T7w6OMdJ7nAXvcQtLer/nG7zSVANc2/Iwpo71hOcjHgg/3Mzm
QvcHYeq+Bj6q8PX6GyDvDFbiWp5O31xYqQNUnN73qtdXNLqNvIdYPtRAXV/T1Lmr
SphyPBuU75p2V1OpXGu3lfesNst+peZvoH5QbeWzJ46KLbNGg677kwaDoCWAQ1im
VdhI9jL4mpvQV0DAHeZjLLp+ZhX/YA7I73BHuIpxfcTo+jMbe7EcaVp74ltItdFt
M6/0vNMpR1ROZh53fjndR6eeeY/7Uz9oHo28+tgOcedu3/oqWnVedZDLS3fShk7i
4Al3FAR7/wVZ0a9Sg/Ih9fGgroIuklRkbE7TP9RIEC/FPt8xeUQ/ttWx1pvq8IbC
v4FB6HPmGim8bb30hYAetnJSVf+AKCo0zJETA4FrwW7P//SGNOeGW6VHIDiMqPFb
Yl5deBUDxYYHkRIXiLS1ke3kDGclJfZU2jhfxFy7wP6zpVLer1Vo1hJmjSkBrpyt
UZG7A8iNK7Y1PaAdCzMm3ixqS0o1rRYLO5zQhkLNDqZPvTxZfIRLf6F4HA8B1pID
vX9S8ayan9QTa1ufobMUkr7EMpCaE+L1VQG02DkP2cG77ZGvwB/RGCZbxQeYScPs
+LTCmZYjg6bsxd/DvgcZiKb5+sVu8DqSyLLvJ+icF+uHbjvNn8XwnYdtSzfmdRI4
5T4WAIIhNeQ4U8xvOLz8aJx6UKtdNeRwbDEV+Tmdb6KS2vv2psvyvCK1cUgyL4ba
TgDfDm7Rr7GxTvDxLd/Ru3s2JOcp6RoH7MFkOqE0u8/IJUoCm9Y9184xgN/U1rE7
2PhWNr6sb0kYy9HccCdRf6QKphPnpVkkgt9ONUTIsKeSUD8EgzTByE1gsmy79eI6
EkwSvazDyBCAYnLA3Aj0iCcN9hZimYGpCuooT1r9VdDLgPV8G1NZqZ+7zKSSl7wW
vBklKDSjwcZS/9Kvz+PXg0w3JdAbMNlJWIYPsrkprLlQjlVjWCMe7dm8zhvzlW5O
2iHMKN7xxBz3P4XlzRhC3dCDdYexbcOGcrF5Qc9n3U8BhVhlDFb61LUtZCxnxC/b
3bMDNBSVFlHFSVuFTGFlLW045YTR73LPmRRzctYweuVV1gnRLm5rZ1YNSYWzRBXI
akrjyxup8SJPa8ro5beaRH3up5Hwje2BHj9n9BSgOoUr0D1N5mdb9vZRGAEx+MT1
irVxxj5ume5J2IFrbCSm/Cdi8tBvYQw7BfRUnhOWE/e9aP4ZEi4IUyQ3msAb8SFf
1bxwvIv/tIP5qk1nsa6tyoYiyZqIBPoMvbp+tpyH9AZIZnSYn+auTdSVEoFadT2x
zrmCfY8USKf0CIUxRHNji9U6KgDdGEXYY3AvijiI8+4EWlExDfSdENeYziTZEmkA
FYaJNoClTaNj5u1pSGnLcAqCZCHDmiyimhbUURQjVnMmkTepNlu6cLhcjdpzhN2z
6kbArJgZo3Evk4pZ33+wb3p5lTnWphVxAbN0kgEG7nqqOhf9hp1y4wZc/9nO+lyx
xTPnyU46izjL0q3xsBkRiHgomAMCNuGPWMPgkD4LrmoUCDez2QXvw20tRyWUndRA
RYvKXkXO1X5AM2XlWC5iv9FYVbNVm2FDuV9LUAqmENIxsLvDZcG5B2rmyYJjfQ16
62zJtqOR0evBIm7hdOEWx51Tfj6i3VNgolTDRNnMoLNb1nhjvIYh2k1Y0jxAobA4
8T/7gJIzvSAIOcSUSXuDZbEASxgTfMLdx5BJd5niX/MWRDzM4Hy7sfsQMC8d7RId
xs1PuQ4XXedIZV/damraxmgqDnd2OOf1zJ350gPizc7dlwkmQrYTKUvQYM4yX/Rl
n9BIUzcO+daQLH1Ou41rK6xgqm3dHbwf/H8zZlzLXHwDZhjuZmCDLzfSrv7SlYBB
53fq0pZTDzW7rLTIB6AcaHoX1DFt+VMcT/TBYc0Wyn1Bz0iIaoel9MEGabBdzasT
W+zX4/nCH8EcVOvqrB+vWKeWQlz6WNUFISrfwxTMvZ3CmR2iVqEczuhyBeVi9+oZ
D6FLaSSxLKhDKgWCsnDOuvwoitxfmMNbfuq1Bz1Hz6hPLepq8is0QXQT94nHOf6l
rrWt6vlJ7tHV0dcnz16TQBI3/vvTxMf3ERGWy2Lb5RjCUbPGBje5Ys1iuyKdU0NT
rENivRrCkt+1/5ZtKwp+VFF9dAVsMlUKbVbH4w9RC14ja6viHMeCG31QnQ1YjFaI
l+G1scJExuI4Vb8ujyVCHlqWGKKolk1W3GSal9I8Gh6vjp8lCebE4yIZM70di0yP
Pa9PuhiNl8Phx1n/b4uzEEEp2uZ3Gt6Dra4zul/BJc8nolFPaiPOJhqJQhzDlAbw
Lut+mlwBdTQJfsChMdoGK3S/cbKGdF/X+cpQb+aooUs6uSOBEGnfe3PVcPb0Ry46
lN6BB0uP1kZCHFu1dcADKz9d+iy1b2eGMjFrOz+7PJNtEAl3PB6e5cS742D50XGI
emh025xVKVB2Q0GsntWYq2wr42YE3f9kAhDRXzfHa38jDUId9v77HUt3v3tjpiwH
KS4Ft59a+AulOv5J+4HXoulk5fqtWqkr3SvnHHeEBlNzVajkW9Jd+S7L188aUdre
yvoTi0rHbg3o1f/niaPaCUfN86h67Wvb8JwXvDB1O0QfSG2WOEGCn+Nh1zbTu3+d
2mGlXUd7HcxP1M/b2XkbzpNDG5Z//C0A1dQAclUM/3JpKFbxPwMtjeuq4/AbE+Ow
5J6/qAowWv+FSbme0Pbotuau/RG0BUI0dHr/05CBX6kkWxO0c4qIWRk1MXtTkWNO
CNovgs9iIK55J32o4tJ1nquA4A05GKtk/6L6TW8v90Pea2wB1RNw4dSvovYqAZmD
IzKu0Y6vjVr9XLqzzTDXijIJOkEGxgiWNig70HKJ/T7Ea88CpqZ9y3svV+8TUdwj
RTUs3qWQamcGfGOKzR1bAcgIYrNbWqDEPAA6zVdzEIkR2hFjZBTVbmZqGD4035qh
w1hZ9dSTdNAktXaBVrSPUvzEx7C4ExIGbQO5W7Ba3LN76zkdpugbhPVqvHSom+48
w520uzMgpttptXr8+kjPdOKlILzudx+9p0HTNiI5mifV/77i/0br9RbDKnWQYG6o
yvQTCcQRDxhIJNTAqKBciza6gzgmKjzvaxxxe3G45i5ciWWrhiTxATRPK2F0K60Y
GWuE1DZlxvy7bLQ5awT9IjRVooYDgTi0EbjKc8/Oab4r+BVesO73E+ErxX/bpCyA
ACulSdOwCAW9W542XzjT9ajy2DTOdIi/941Pr2+AKT+1oDX4/ML42ZghwgA9Jwrl
M8bbff5E5Ykkvs67Ev3WC9JIMW81XG2lSYxbIvI7Ekqw8nOOWVI7I8TZMKam6l3X
DqScSoL/Im+611HxTA4vVkPNzwe6y5iQpc855q+On5/fbaCOvhOCmmJ8MBfjxL/B
AEnk/O0lOaWJEKEO6x7lXjOdMF291n23ncV8uW6p3VH34Y+K7s1X3TTp9EneHPKv
FKOt73iupob9QYoaoeojBoNsiJo6Y7QGs5eqeQXKdcd2bkSG1wt5hOpc20wZJ9EV
mDHXRT08Nn8D2xGd5Xkfv0m9Syy5q9V8gEULKLDAd1q1KkKtnRW4plTdMcfuiLOD
dDAQL31c+DwnoS6XoPF/4JJT1yipe1IS7kTxQ0Zi6fIeY6W4meg9UlD5zuxHLsJH
jQuzRVy6sELCNnv0UkDKr+sA7w8a1YPuA2PO8P/niyZP5fwlDficSMm+xKh145OO
+HrY+7GWyIvh9uUqfaVvplgnkCqrjldYq7eSNBnzyjzn8+f4UdpF/vUEpSpuABaI
znZ0Bd/sbAZ/sCp3hKtMv3wpVTy/MqgC9Y1rckE3D4ohupRKX4TjheqI0FSqbAKI
kXFfylFgBKq9fUrpbWLhsZR1p+oOqmzskfDVkP76X3zWvsdd71S3qfvPnZgapSis
RptTOMEa7afqTzsMBQFVxHavbTwAFjtiUgqgiWVsm8wmeMjzRNg8GfDRd/QCw/cR
eVO6u8V9rkvSdKxb7MpvgqcvsG4AJo13i9beQjf0wjO97/cPbirScuo7ZE+QEBCl
1QiWKrIYiOrr6A6hJN49xE8qTO8EZPKICTN4G71srgQcQ8D1YJTEwb77wIPhRJa6
8fToEnepVAAntgComojFquzB48eH9S9h5ll38bULWKVwZ+/PZ46N5rvUfHtGQ3/E
7wXysh9SosmQYPd7wdSxsBkVzg5UIGI4No+Cv9KODrci4nIdr0NdDn2omQTnS5Zy
FtDuWv0QZnUZ5t6S01zaQTcAxuU/JdBI8gERvFnzE46pSWRldeipSHbw21mM1O69
OP8yqS5JNXIRzPehILMUJonwSpoBxtncyOVe6IzFAjJfcN+IhJIvjL9bOBqLtDWW
yZdKg7iKMthlR08ikMcIAAnB90NmtsgeaQYgN81OAPfh9FNQ/+hLcqfB4vsBk9NU
OyzPLztvaRV1zSs5Dr7mpqym2yBazRCjM1GrKGuUev43ZIkbg08eUnwAnu6mrpXm
GUX31G4Us0/4lqKp04OU7HWserX2/mZLNrEGsg08P7SBRjkCXu7ZCqGLij2yC+3s
N/WqY7Blbp0N1zD//bMPVOKkhCIu85NqbA+Km0P94YHOJEMb4tyGxyrngmwEAhuX
N1s5DYv0C30QETvGMiR7S3aEonv7wk3gHZekcWTFRTI4K/bWcsULiQxoBlV8LC2F
d2ZCj71u4CLwWxs+7N1ZtvaPUbzKfiKLi6fm5tEuYIDU3NzrfctDv4GdGPSZBUuN
qEJ2teS0iC5cqk7zbSlrZGWVjtMKYdS11N4OoleyFr8216nN9com9s2AKLAik8hq
nllQrOPBknReYB1vOEbR2oF8V1gYswsgOERmxvpK3EWLThjEwO+1p+/M8N89Vtij
VznhHRmSw9yDBjbHhmTCW/0olBF2Wk1CcQ6CE/Uw2aWVj8Ka+ev+wMZzWxiOcVGt
OBKAeKvgKwM7zS2+llyyXrHpUahMitC/UaNdqf6kRlI3B5rivu1YuREO4qwJCNEl
+RSlJWTyftmvaCLxJRSVKCdOOzdafT/ErCNUlaeJr5aSYqUsAHaqhGZcVVzYgY5q
+04XwdT3EHOKpS2/aAb56rrgXM7iK7v5PAoE8/NgmhIJg8k8sOMhynxEebMy9l8d
FcCVV1Lis5OC7BEgyYzeaoPubk/Hnd+ed1f6GoHSDehKodcDYwC6fOBci7AK12Fv
e3Sh1RscLTG0ePWl3RI2ShvPp/x4az0vS/K8/DIUx8gASj7J7xQhwd61xxFf2jc+
LrPuOHLEZkMTJFk7nj/L9oRALudCLgYRTiUveR7wBdGm3Bjd59ydDIbhPMeNQRCd
W65XfAUrExO+877296uoh9/vRJuLE6mPQNCJ73wRvFewNCo3J7X1LJIFxTOej1nn
Jd6U/r/IEJLTcDo97v+vNIJpdxWx2YRWAtoqxt1csyCI03DfOi2IWHI8Uv4Tj6fO
Be34yNSPnV74x7oF7Y71pPYVXBge4QTCL39eYbzfbtpzNCN9Aqr/7Q+0rli9FEEM
D8JUS0eQAczECNeNrO65S7n1h8NbTgmwLtCJ/XzoHXXtOEetkKI0M1X/KH6Wbwko
1YzzdUAc0d9y4YPen6eY+TjQahOMin10cDs9fAmJB1g31KcpYurCltYDNp6d1W7x
jT4zH0AOrEJqnWhMyGYQGvdjUO2EpceUNC1bpyKoT1/oVWgmOoJ+WdQIuFINh5m4
4DklqfQetQZk0DA4951+w76KBB8EJyI7DIHazTz3zCNyWmBWAHnBPb2OGaSYfxEc
QpF8/a//pxyqJ0bUOjKe9CXnwiG5dZ3NeCI+uqABN4hXVJi7ARgf/cfbdR5/72bC
V2C8lMfDtgpok5FlPRCOs/9Ijecen3KF8f+bGSRWRpfk5lTwwmgvswUtxwu+MZal
+y8jTjCMg8VZIX9Pgri5TRFRYjmQ6rgMM+ADp9aq9cSZbKnsqqDQsokPur7T/DX9
OdqN64LjZDnEATF+FdODzSQ4iZPm+D+AZBZhhEoqik1vkGztrpP8n0Mk8YPoLSnj
AHf8qZQUMR2gAh+7Z69l9KDmvlRF2goa3/2GQW+7tu3MwnaYBZ3NxjkQZXggXV2Y
kCUFqE6YhyNhu9q7+lemmox7b1Rvg3agvTY5m1zuLbdA/0y6oPKHE0ESpeDhkWsX
ZomI6LqNIjmdoMgraEGNSOrNBxDkcvWk1IoBoFRSXWWQrkBR1uriS0V6csz5F83h
KjfBiXeG7RMyP2ktFVbMbjN4r+b1W18p7liKzOMMjxCYSjBCT++ryl8m3k/2yrnW
ymVBlmPoJFGwSioJf47X5zmPiIzl1iQGt7Sqruq+aYJ+ZMiPshZbsMmC3IE85MFe
C+c712D4M8nvvgJr8jdLbUKOqwzGsz1bj9Ii03kZP0R1DZBzroQ77jXT6cEvMZHx
xwtfG0KewSSdxd3MRzjDA2Z7h7bUP08DeisXZNthc3BEMjifTxekqDMbBICISfOE
ah0lVFrrqnyPyC2It1eDz1gM/7Dc9ZgDcSjPzC6KwkN0lpSu1epVpDFLmDwZpAjL
mWxu2zzR4wvOL8T2RKgux4XOv+M1N8ZZPSi3YNT5w3VjZoo8Unz/Hx7AyjoN2rC/
EYrbo44sOtEtQtyPwXzFfneH8VhBnJ9gZFL1wCX3tI4zzEJKBlrnD+EBr/2dDr4J
OIThaMlMqIxqiRre1DUTEmVsyL2aOQj/ZN7jvEfRaFAALpUmDKFaKaK8XdQxk1xW
iM2LapHNJt1ootjtFTCwQate40GFN2CLyxVGKmDyE090bZlYZcES/W2HSwkMOh8P
VsNxHXFIQyhrzDL/fpWmWukLB354nnG1SF9O/Wyb7KpBErk0/7dOoqsm7rsVooBG
E5tWz2SS+yUaT28fi7xzltr/koF25RXQdr94a0bEUGhqLoNgWTXM+7vqzzeMsMvB
vqSvozmyvPqCTfES7/AIrHK70zbXCsbreY0oaZQG81HAqWZE0pYcr4vKu6U37fuR
9mXU5v5pYiqPcQdYx8WjDo6ejkXZoo6fjrrx2oMn6C1dFaQvGVA4LdqhCutV+UmM
EMzeBe9xYNi2Nu4i2hPfStm3pPSe61BInFQaYaRDr0vEIOEyQ0gD3ECj7YUsiIUu
Sp3QkdrS2qC0U55hgBhr7R8cMmc2P4ddVVg5hZg65hww8CGgvVdWlkYcsAl1g6H8
OuHZ/++4nMQb/I85WzPVtFuA3xyQ+mVyHkNBdrnzP1wfpjCXi1XTyljSA8mQGhFo
Qq0LQFkojUq+GuHcYHi0ZJfU8bY43jOYJeDnkmj++aFg9U/oDm0gdwjbv4Q4sxUN
YyYvLThoCXMXuxkEidHH77gDr8Ea91mjlRZYodCWGf02AY64/mVp1NsCTd7GQZSJ
iak04iGYG7DzfSGPtH00RPfVVap8lE06nBXbRh2s9EhMFRXa+WmTrB9Ll7GGYdk5
YNKZES3G39yGSx2OnRX6rJG8rpKPn9VqUMGAEid9qjrPVQJLaGu8O3i1Tg4v6LDL
2oMZ7ZeBaUrVd0Y96yvppfegJb5vanYxwfZxCn2aV916SX2hxgJDYPi9w0HLlbXX
2iZb2vhD9nMAjdChcYAkYt4oLtK19Jsw3zdK7eP2O3k0OTpA5tUdKdaFQZTSrGk6
LxBiNcybdsRPYnCrYr3+oMbGmqIy+isbSoZ++cxXj33eXq4tWmqsJhfS5eCB9pui
R1hSEuXYy6T6jxQyk4nKrzpHPnBgt9DVJHZ++ofaIAEcBCkk80JWr8gn2kpkqo/7
Pm0fBKStQuhXS6Q5E3sClVtkN8VuCGKJuVpeq1ngNf79t+GTBr/DxhPDWgo/Y3ml
LwkdO8ZkynxCK0nkPa+eH5iE77mo5L5oRSN/5eC1OmkFJLh14G+0XN2AuA7+TjEI
Po7Hm6HzxobYLvqaED4Bs6UGowP9RwVgIUam9vqMXecRmF0y+tBshYUNpPRaTzoh
yjczKTt9RmgNcooNnV+/nJsYV54jOT6Gog33pqmQx/KRylGnvvBIe5Q3hM9X/tIa
DHPEOlLtUXitxdk2d/0AYJIDLFOsY6ipkitGAFA3LIOXD+J6KgTlTjEg/B0gGip3
AHQ1t4b+ncacHORcDUbF0YpKyuGTcgedCaG2C2Xuh2IvdOouvILji9hvLniJBEVi
lEqgyL6i8MkYVYAD9EctXy5ZDA1B/biO0Z3TzQkDTe5X16YbV15VRec9qlrmHsBJ
9F7MULU2a0dDAOsJTpJaXlcOKuPTmGbcLMNy+96tuj3uka7j60Dt19mKbZJ5HTNI
+GZHzUcae41YPQzhdwtjYr8kibLmi+D/b85GUr1/HgrBC57XleOehr8QUZr6XtvW
q7uKFgLYe8T2u7RoEqQW1UD5FCZbGbeElfLensmvVPJcxytSIrSSytunGlrn+VWH
73bOsOR8cEiNsjiauv3a5Zx240zrbrNaKsGePNihkA95csqQjn5MYEVeIEL3E2W9
YWH+Z3rxGxYdY1ikqc23GAtvZcTdIc6eoQS2eAlvvbVGPGwERIn416LOz9qBZyR1
7rdyYKjwoUnAjjmvIyENQRDxyJz6BMeyRwLAVGZPb34Ys4dPIG07dxWq2oA9ynhN
/paaS/E3iDONQf6u1ZbCrbGpDrBYT9T0IPIwGo8GIQaAZE0YEklfi1SDJC5fGpyW
af9XvrZwKCXFUWvI/GrqsTgn/ySj2eaLYXerMEUmu2Q8BoIE9hScMR8GD9k4AM3j
6syeR9RLjac5dd3zeTSrj+IUYXQsFxd5BdNAcv1R9LMh3PClcee907r1kcNHigUQ
K4zEvr4d+GMib9hRSFobbzWqV1yTCITLfZGEsWYWNe6ajoFIR1ERmmX64BaA2orc
OTiIvbImzz/3CjL23yoa2OHgrxdfEBs3+susNM/srp8EL0FYp7BLgplFwE5LrZHx
GbGx4N4kgUgR6qKyj+rnl1jOVxugM4VOrWNZ9irHq9qW5Pi3UbP8pW/mGq0otFZ7
UOJin6BUD3z+VeQ1Vi5RAAVqLl/EikhbAsBS9pzE43GsDt99bewFKDzvYb+QB3cc
3haJDs1PGupJdi/3yWanY4F6Fyd9bBCZExMLhrs23IX8PAI2Jo0s+NrbulRnZWWu
XsOYyLKxj04/Go1J2hzTI9hePDPEy24VeruFdUczZ2d6sdFfC/LBgoCDHHlqH9I1
1/yPfT6052t3lS1tvPYdCi4asqdAQDln+7budG26yGEDfLjvY7JP18kHgwgPcudZ
RsPA90fitsdkzhCJ8/N9msCtE9oX6WNaTDTvIGREuj8U/qpB6BljxdhMGlG4AQjJ
7I6EO0JuugfFFyQbSp7Xkb7qL2ql5AjVw62KBZfFBRxlLSo/pNJNjdHKdrMULlhu
Db61AjJayGLFC7QOuKl/y+oyvnq5eqBggwfgJg+EdkppmS6nmMczPV/JmORkhO0v
5tpAzzvQXQSvozCtFdc7xDNh4dM2rjdMX+jv4AkvkGIm5w4RdzJ5GVeZKnF4pcOG
XCLqcE+G4ZvN4mKgZqPmqG3gViCpU7avt5UosIDuTs1N6L8RnVnWSRGlz4GoeybE
9w4xia/qlyDTG3qbw6U0uaesYT1NIgLAFPhgSG+vxVQKhtfV1xUoKn2aTHXkQ342
LSixzb4JhNRq1HK20heqyWeABC/Y0FxWOiIrlyVPwaPbANZ3BZiGp35HAUCvunop
CnQqpR6KuOzHDCEPcCBN/yfoMYGPgCfMwjZwG/DzOWJtmHb9qLjDySqdIk8C2hHv
0neQQ3+9o4L+Id898oV/EETuro+ta+hvRy1H63agv5Q+Y+an+zvIMq7V58TxBg/u
8zQnw6GO8TKyEBR9xtD3+hxuSRFEl7guYB9hl0U856ty4VKYBuFpcqsuDga/enpI
1CWPd8LPnAz6IAIwRenZ1KJziNMfB/dvWy0LAcgSXay43FLfhczndYV6Yib36jP8
3m2nS8ezlbhzjdsxPcIrfkqieKUZOsr6ac2uaWDn+kHCIlKQ8Fft9pzAO7QR07EX
p5PP4aFE8OCCfQNZFvT3NIMYlcAVdy1rI5VoQHqcA8RrDE1Dlb/csVMDYNDOnX0p
mWOtwkqiM+BJ/5kcdjruRbc6sqCiyCV1ijwb7dshOQL3raBBPeOYkXOCIqydYpMi
GBeIKF7Gtyg5lwbB3JNvGqnpeNVg9PlHqyJdbclNRs2Ld8XLecan+ec+Vdwg7CEr
k9csApnQ9xUbd60V3+Cftes98Md7cN9NR0+lrxVyt0HASaaYOi5jvMlvxvqowWlA
OhYUferMhtomoy4TklOV5OcZg9YZmQ+RzcK1pWrldVt2fukRIr1ItFTogrDzTS0Z
cVd3Wfg+7aGgZZ/vevGAcNida3wFF/Xba0nkskTHvh/AbN51yAqM5mYHMONC+gNX
8B6qdFhlHFIVDof4vIpSbilkmKB+PrxD5R3grTiGo9TeqMA/a+UETLGSUgpi8Ch9
XIliSvOvStruA9MbG2oTuu1MtXRKjuFcoHDQoUgw1JURX4dMhXIbGD7TdaAaO1lW
XRrVNqS1nhyPEPUHFbOF8Ido1GU7jZtgoEM5FbykbIqm00L1yhYHIIbNfRuE6z97
YL4LYfAP2Ib8edwa46lQyo8YzvAPIqzSt7XiXuXk5OQIkqPgO5ytmZAXyx3ryP5f
X9BBMfZ8f7rhBGm8e4D2vOux+AcNDwo5bjAtWO3b2PRJAKnY6P991Qhqd2iSrKz6
3EerAw0GJZ26E63mIhLCb167JOtr4G6K7cWopbGXkn2/AqqxJZveWftLMFNg0BVT
GOZy/IyON91SmOjxIugzVJW3+NAsLVj4ZS9niJBH/KZhyVPStbiintNLZxm/2sSv
Oo6Zmtmam6kqOEcdwQ5faFuaccHFKedGfMQRnAJneLkOhohROXUpR7zgVNhAsUMn
4kf8mFRNIaHFGQBUeKefzd9V3n8ADUnAL5j3CT2lhiCamv0A6IRGiS0u3Sw2E3VY
JWOpR8Czn7TpVChvDzLMODxBRFA+I4b8pDAo6SIgMupPpdMr/KBsabbWlgiRm43S
FS+Q5kKB69cWhBRuURHFRpt7aV8hz0sZGdqrdKdDhXdaasZOlo/Zv/HJPZocQh7Y
Mj3s9DzfkUeO6M0CzSiieOH2F40xvSrFAUxx+XMHagDSS+k1S2jpXu5Y69Ma+N1S
mkYHxLXCyP4P+IP0XPoOYjsXdcRPWevjEkiMfOX/iUKsqAf863huIVXkeXgmaiG8
HxFeqzctnqcLycA1Xhmb/Mhssiuw6EhNp56xhxx3ENDQYoI2XibwEN2a2vgaA6Ve
AbKypMBqb4D8CJudUBXUyVYDJIWz2zNDwLHhW6evsgtGDiMP4TY/3v1eNG2lTQF6
qjmCz4kfdh2YxbxhBoTXRpOu0xUvxGv1JXzxMZXH3ROw7SemIAPR0qo6u0BEldWS
raIAG9zrKzlofM7lwkB4s2+UFfGOvhBs/P0dhb6NhtB8Y5qfQZ7vxcJ1GD4E+rRc
4mSE6JUXcPSVumcFHG2puGz9YORWwasTzU/rnkjvX6WofFxmAnnHW7wNGxU/MVAY
8kBlKTB6+3fAY/RhGM4tfQDzbdU+nctgTFBb4AGKYsYv+KgKnabCxzvheKipzHC8
E1UXGgt7o0M97LSTiqvosN8lMhRNROqgst044Jyw5S6HuMQJtQR0Byb9vHb4Kl0f
zCSnsx17Fxr4HobLuRN5cBzLtU8pxIb3N0mMPUZ5io92mbVgGyHrRcjLNfqUHh0u
QuM4JyOAe7mQeAKP3G8zZVszfZ8iMAxWUjfY6PVoLBi2AU+PE//lprnut/2hCMvZ
jzDK3osSQiFsP0O2yvswnKWbTS5uGWqG3pbIhQwRY+s7r/CT9lqNKSv6gCcldKBD
pxaGV6Ay7cEtKfdQsixlWgzhaFW6xuV6khncLUVslu8YClBzKuL5Pi5Uk0HRVyAU
6dSQ/3Fxwhv9RydxZy/nD7SX8DEEGtk9HdawFQc6ngTpddi2vlb8D7fs0ySBUZy9
EhMT5CRaiix/+/UjEEp7UmSUhGmfw8dgCVt2IKHyQCekAIQN1XTtH8am/EeHv+uM
YOSru0/IJMcXflALneImOXFi3fwerE5bDi4UzHdk9nUySF7vGuwOh34GoXzga5rh
rZ39GGHWJ7r/FXu+m7XI6T9WKdwteHLaFwKIlo3VspPg9+ASYFn3geTx1faI0/CE
jycXXugwr2Bw9ZvMmF+JU7ksPBb6YGIMzqm85bRwfsoHX74cIkm5vpgo3QmE1+YG
NUeDPrw8dXFfK4Oj2Sn1MD6UVIPbIaC3gcmginAWlO52AtbnGRHtTqym08qPWe7g
fS0dYPppIfp3+WbyeLniSSSw80aGdOq1ZCBs0+g2y8d8xXWxtMnDPQRlN1mptB/6
djT8NEeVCBFBhQZANGDZIqfCiL6nfKkQjAYsPoWPzPtbqDVkfRm+N7sXdjvS0K5n
vJGo9m0BtdQFoXqeM5mkh0uU1c8RxKL6y1sEU2OHA3CLZg00+08Xf/HHJvHwytQa
e4xz2Lanhz0U1mg/bHChSDNEEuj2Tie+il0QbUrazvpdn71K+EV8cO4+l1E1S19D
4EeP8PXjApO4RR90PjxPsqeNONPWtMpAgbEfYbQ9sz5pcyRWcwrqUKvApv1vDWkA
vwaff+kUBL6UL+Qb4ue5bnkLPf0G4vpB/8885GnNIGwaeuLV7DLrls40D0fefShi
Bb0ox469sas3XvrFc6+ZAwi2MecefKuprkoRuoDDkNfLY7ZVEdLSAlD32zK+N128
2fk7G7c/ZMYvDhoVymxqcL/GLm84x29loSxcIwBODYkfu4+vj2EEH3lne3ZS1mOw
YiC81jfzCdGHDiEGGjdd+8XbnIczJkeNELgmhPWg2Jbg0Wi8pDMExTaavU4to06k
INjNBYszacfVhvEd2962RRGq/Gesgb7wI1ou6xH/sMDjyMW29O89cnMXLV8TN5w9
DA1udUJ/4pWoSLUcxMDqpBtXCxl/+7eWfFVplW9oIePuctDEFyPcaDJ6p3kknjMr
abJua7kIG3SX3OHqXrhDGVX2OPJ93iBUSYKcKyO7MLW/sljeysRvZJsHYskTxalK
C57KGESUuoZ3aycIuLExMbaSw8iV7tjXr/xSq4yMwHEjHkPTw02ZiYjcUKEMM/yO
NmZeR8U347pb1z7CrctpDKMFqeg6N2XD2QjxX7oVnPBmKbzpazSMyL3/rpjv+1GU
IomccqsSqpsTzwisYxquDd9zbNvDDfrLutiCQytk0Boq6umhJycwBYjnzv9/6Y/L
1QwXWfUeHlF79cVzkJa2SgMR/sV7XsBcnT2X3XQ6ML/3eiNJnU+ui2it/gpjvgJQ
fOEqZ3NJlSAL6WXZll0YcfNjThSlxpj9/E7bjm4MxwwNEJDD6Efq4B34+ILH1vVi
QHN2t2cIuvbKRAWXFATx+IkIyBY4Af+LhmJJQDDHDwgh6Us54DQ/CUKR8WuoVynZ
t7DvIqGi76M51fz6G8lq5Dc9kY8ceI9HnIraYTLCb+fF0HDyMKp9T8DiW9LzacLc
UnAM4StVQVWI+22XR2xL5sPr/vIwPyHYmdwrvsMfADajYHS1WzyzVrDQzBRSQp+R
ZNMooVWe4BEIFYQ+NGKdy11FRreJHoTx8m6UQ6zPggmXaVxy+K+Tmt2zIwhNRvEA
e1rNMW217Eu0nRlnByq9CebI+2MF9TJgAfNIrG7gpSlZxtR4qE9hk4PhtWwk5FJH
78Wy9+ECNT7tLRyiMhOrX6XtG2AS2XPtVjyCAR09Bwu2ql/5TIfnnlkkECmr1blt
THNkLHyc/p1Lfl1Hf9/s/kFV/hPBJpODLpJoADMlqYhV5ISODgZ1xUPTdde8J4cD
4pxbW+TtWiYFcb+NQ7osCSvtUhpmLDd4vfWfvXih8UqtVgi+8L/TPHOAr3pVUnGM
D9Xjbz8tMI2wZMmBgpV8p6OGwrrsiGW3IahRK4nMbkTJuwTFwsYrdkjhixeHTnqv
MNcuDCz9+qHD/RggFHcndAJa4pds6Cm4EVZhm3TVDxSMEtxzOB5yYdP8VXR7yn6+
+Io9YAtWji4fDdHwiyHcrNeJdKrZd9l9x281RrC2XjwxjNqmlauNvozi8Q0jvf6G
lymvgB8bZ1rGqBNpxpXt86GmPddeIz0WmViNoe7vcvnsguwzRbWOMDz+yF8bSMDC
R72Lf49eCiskwSLlnhYc8MP9ReFXYRMvY7AxfbgVprexewty5Ot7EvDRGdNnhmEZ
Ux9/L3ruf28b/+iAYlntNRuMi5gWJv6YS8QhoVKdBSz9rDoJLXv1DZJ4P8/ssnoE
2M80jvdp9xPiJm6USZ5dFb0pDT+Ue+k8hmGNBBhk/PSANO1fBr/vFlUWBvsfCjTP
A0qnNkLdL+R7ttBocK8pqgviF4B3Ekpx/PyZzQrXCzo0ngkfe0qaS3Nwvgo3i4ys
I3iY3qVXxIkZhC3M3iSlL1mpZqt5deUf+c+X6zvEWUd15BrABCj+SJFk+/Ar97JU
+ZCUZxGlqOf8MqYBEIpEo2xGoARS/17IgFiRZ0OfISSIcv44fOmbfXw/hNEpnpVU
AvP23XrB65ZCfHcAe3DDNhDA2Lt8/eccbA6QR0pSFSC5+WGlPn4PG6TocZejj7W3
pSPdeXRzpCwoUXoGd48Qc8wL8iRfIyJgzqMsM4R7O+jGljF+NiR83XaikYvF25Sa
Fo79eqWj1HQlP7kliaXj8v9sFsAox6/D8ZswnM7EWSFkoQtF9yrVAxDKnRU5dJHL
eYi+XApoH5boNXkSH3nsL5nWK9NANeES8NKLPBfYR/fsi0t/B71Iz4nCfB2/Ooa3
mBRcDT6xMAt8PluqYHk5JlhTW9c5q97RZ1J+IdMvafEAc/EFOuNQAIEfnBUVzksA
QdPDOGvS/CDmDajX0J81Wp1AZV9j54hdoVpozxMaiam90RpgWry4xExLxNsuzq5/
+IISoZicI4kpHseMJrPfdJUL4ep23nTz1hci1kqfs6upjUH1xbaJQhJxF9ZT8Vyz
JL2HHr7p1KcPNI2fmLmOOqzL7oXqFPeB68+xiyTT5zUFEQD4SfrfcZwtLLfn//lH
NewoUiBSP9yA8HtOzLjeJCyoEZ+oWs73t+JXEbHFmjlzm7lZNWvvDIx3zmvJD79z
pYY3poUJj3cvB8OFLkQvdStxLtnpaYg7nPoKJNnVFwcNaoXYbvYrejq2Ik7vTDb9
zlZVCDwdi0vIhbUlUxNjHsPjcyhp2wTnXJuO6jfr/0bzlCtQICFo7KMGQlD+O8n0
IJnn9reY3wBQDStTj7TXM35TqeTbAQMAC8sOkAEFZ3hB8gJz02UWtneO/NVFq9x9
s7KWboJEGy9I2L/peuGPIskXTW4hAKTuyv8/f2b16qQqiuG5XY/74xe5WFvn7M1S
3wkmORa/bRvC001dKREbFQyyJ3TJIDxaZFcgB9S71W+twWVLLOPCodeI5wAIRoD7
itMnbPII5hnWC+Zyf4T4SrzkksXbdx01TLiPm0KRlzip+rYMUbDiAFOjfo7RqBbc
51JQ9UTBL/BwQjKxAEC7L5XyZf7nIxkOUceyOSK2qg9LNO9MN0CKRWsirNuSjWxB
4AVx0zowR9sHupVhxmxGb9Y83/XvvaWPcKmKQVuGy6qB6Rf3g6COo7lhUbnL9mQ/
C1DMfG4L7bB6JGY2Yqw3mrPJP0fOdaRDIUOMce+IVj2A6AV0CCZXDwtB8X4hmliK
ZuJtIshtYBWSoh5Mnu5GBwEY94g0lWs2gJ8uYlAHfzvUaswSPuXaBCatl2ZAqnH8
rZ+O8ef/ly5FpOLkDFBbHHr2mUEICQjFbLvhh/UyyYFinD7UZ2em1WP1VAhmEWAq
DRmLMuRZraaGgmjR0K140ahaKyxzVuddbRBzC60IjpnBXaoPEJdJLVD6tezJkbnh
89PmrnQJIWoYIaORXP396gVJdKUZpUF5QBlgGCr2Yrd4KaxTZAxE4wU/KKXb/G86
U3qbkNKDrfe9cKd6pk9xono1QJ2mR4kqhbxiB4Mh6RNpiqhBnn+V+8BJlu9ffPbY
gu2h9qxtwf25EX0UTfRSKeSeoGuAmx7/ylKQBiFw7PHQi5XR5GS1h1hAotYXRWQq
R7xr8FdzOEiQHFsfEa5S2dzgNPxKgFJWPtVVb8Squ/M8E7RhVt9mHViQLNBEXV7g
n5c4mVmDbBOUF594Z4BhzsYVh9dQhwSiz2TxNKGeZl8xJ5izosR2mnRJtzVSSLu4
ksH0QOIDeYSERUZ6z9xYEg0/2kllU4uAv40um22wZIC+5mKPHsda4E9B5058slEv
IfvUmog0PLHa81fw4tl+HLzZn/7M9jnjhBjOpVtvbtS9/I+O2ms7cC+tSVyAu+1U
qXggl5I3xawOtnL7e1W2UkLqhwWO+V/8ZZF7WHHZ0ekxUWEtx9UoGNvD4AyDGn9S
NXAY7ItejKNUHS4Wyr5huecAZy0r/lnLWKl6drGY9LnRZnUwRMVzx2PzpYw2DkY4
w8A9tlHPxrG4Nkl+taU58d0Hg4ShOcZT7qwLsTrE6PaBIP/kEMOrjQfyQGIfxi10
uI3mhznZp16VYknpRiQcvpK1p88YejB9zvtjGrzUxkcFa2/wdVqNSGCEirmOr9Oe
x8pbDXfgi8d7/7S4qtOfI9Pwznz8Z3jsR8CtCabIksaSrv0YghIB0AlN6QPwfEhd
gQNcIIiy+S0xZCl++/rt7O/ia6b586fcl/FOwFlkA2q3+N+nfiTxxW6aEXS6q2J2
qWY0lkoAhnRTvBGJaZuGI+c8OSIu8eFMtW84OIWt8oRpfarVBLLHyJcU9uh1QxID
oWq6KysXX6Hqr6zGNwatIbFtF4oC5Noi7NLGnM08SzRfl3qqOm7UUcFFuLxfQUA0
YSKShU9tKgVmvZd3CPN1wFkbM5RCDUauo1g5EkrO2Lii32CozutfsWvEuf7yRWn0
4EvhzaWBYeChjIYtFtb3UdKaexq15Zw9Gvkzpira1tlhbLotnHx2PW6CR8YHF9f9
ZwCpBsLQoUByZI/r8DdCxsiHF3UWipUzqi30Ep85mqkjObpYbpMvx+dWzut4Yktg
aaRj1jgJ0bGZWzQ+tCTXSdU9ScysUPf5AuI32HwuZhE5sAjvfXon4w5c/k3/E7wh
94WQpDGPM47jIGGnLIL/DyeDJ13kMl+S+YEy0VUPTja634936sxcPuhEB7LteLTb
6aB0hZ19ObRHVWPjdtl09WMfVFntNNF0mzRYLjKupA2bHmK/HmgFTN54anmTuAB+
iRMVMr6vaG8tFxYUvDus/ozdvEi42N27tMTWo52QpK/dt6Hj0a/1ho3YOnShR/nA
hOMBoHeZZTH2WaJsAsuI6gQsZc/mR9gVGkePwrKMIl2JA6U90KNUX5Go8bORb1Vf
bBcaMKoTZFvFX3n+6sce6cPbIIGpLcIWPJoAw+nvKwdrGYRPH4Y4zyQogeJSQuHh
FAUHxemCvY01kFikfjzfVRgSQLIQk1PFbY16VIA/A2lbFIaoyhxWHM8x33KqgxrT
9Lw6gGwwn9QyRYEkHwYlZfYGiM6k4wzbTuEctb7cANd5vxYK7sL4pgB5HqdPT1lE
Wvbn203ex/E1Q+3FZIBZsFf4zsRMk75EgKj0C0A+TvEl0dH3MawxPW6dEqZQIKf/
FfubSfx2fbc6eGtAcFHhCAtTBo0+Re749j5ZWxJU6de/24GVUzE32mpW+qFvg6AW
jLgPHtXUaDxoupekG2JkcwGFtvoOC3DN8biO9jXsrnY8xbbOUJ54A/I64BnMTxE8
TP7l8pzdCY6lSa7us0ELMe3+q/RwbAREIjEX4tokzsgklBA3/N0NHsOWb+RPbD0h
LWlaSvVRwdQpUA8NvnrXD9Cam0UUu/MBMRSPM8Iu1y2G4n1QDW8EXdOEfylGsXc7
xd9g1i9KidXTjaB4xTehXmUHj/OVKPC4+xZWzNF2wOVWKD4Un2Bf3f5H3tDgVf2z
3ugGGWV1/AOewyTN8EktXseAmDuLMv2NkPgVUcGGfDGSI4+FGL/iNW9emrTBGpu5
IWNsVuKM3Xr2FplFwJ/CdrwzJ8HEVKpvlDFPxuC7L6GKJJNAbEgfa3L+wjE2BWli
ACWWRS5WN61Kqi7y97iYBAdgNm9aJZorXunfBs8fqcOYVPYml3l9eqCq85TN80/t
DeLKaIXHtp4lKtPuecAZbn6AA13HteJYR0VtRo4RTWWNHLKnVPZSfmgpcTQVCTv3
gYgXVa1uUX1PVPhQuRT0sVPaX9X1mPVP6iatzvL+uzSGrwoju/X3eFe7EEzG/Tww
kVGG+XRckMFq+Q7NkwVsfkgnEUVAT/uzMfEgwexGneHQmsSuwXZkBgQQl9yvThZK
LxKbylv9L/Jw8DO8Iwlj84W6ew6KaaAOFiYGWNkpHs6ntNcEQQ/xicNhBsekkyU8
+mz72MlXbmuV3ugPRfWpadH7Usa8HtZ0kn61ZubFO3r8NEZjGFBGb+3UF6afUYiE
Jd9Xu5YYd3myiNEJixzLvlfm/MQvaie3Q4MXF/0cWI5Hp5rIqb75EdU1CBCxxGb+
ZSp8+/bVzB8+Wuu0BMgI+cywBvFXrfLUnA12jyhZVyJI+UHgXiMWKZa49jOAY6cg
UFlmbb2j1kq7AMTRAyl4mMpshI0Jowq6hvKqa2uX0Q8L7gkSNZWdjHOn9hNCF0rf
fPhwvp9xsVQLDTRP66jLSkbaX+An4omyY9DUY2aOe3w71gHMrmMk4EtVEHxUI6ix
rpwJXj0mo2sbkNjYZVuUrxqZ6qEBYKLLP0wn7yykgU6C913vXGY1Ar4Pc7RqYhWS
k6KU6VvWLRz1HONBdGTtd+ovHXqBAFRIgkcLDVaSwX0KSbHPiSnYlgbtiiVA6nqE
yy9EV6E4RWsNkrtfLrCrsYBob2vK2HjrL/9bz7FVxU4YHT4QSD4Vr1vSIC1EbL3D
61LMwiGrLL/blU8Q5QWkXiEOikGWt/coi9aL60mqGje7SYoE18LXot8PhEhLuQzQ
wJMr1pXjwVI7vS3PbXG5xO8c7chhsMKoqoFlJZDLhYAlWS0l2j8Dp8OVHtyv3KaL
GSMDulbV5LwRBe46J5CX9NzEeFxHhAdjsHZVCJqVAzjjH7Wfnd674VD0uhg5XGJO
K26LLIrwB/49MuyQxlJeRjAfI28K8G7kLCBKWJb/EoUvYMAFp40tbH/ZMS+1S9Xm
/6tDNg/EbLftcoDgHjmo21pfq/ZuHIO1ml+1ANYaNnBakBE/wFApLWeZmUUmlxbA
GkV12JyLoOFLS7M10xS6260atONHKMJOGmd561zkbA8glykU67iF51TnLh+m372K
yDWkw0G1al70iGsueNzcLRBnY1cViX/fWIAnjQYjkpBGuUMHuOghXCrG/nrwJrsm
3eFEAKiQBY7elHjO8P8j+gi7TvlNKdg1tPlVzq58M6daZZ11r6kFQRMCYUnZm+yN
oJWetZtkOOG75Y0mWSPfr6bwX1QcUFG4cLOxSX4y+TLMYMGmqh1y6a8EgIrGeNuV
f4YBdrv37xii8/0k0TtERxzxt9p42T6rvK+cSCYIyhYQQHTJjnKZy31EOzDEipk+
O1RqBRqK0J4oiT4Ihfr5xxdtwc8c3rrs7mlXN7UyHXTxcR6vLVcSx5aZopi62obS
Gyy7s5kj+Dbwf9CAu65jELrMBPlAAb53g1zP/oMdrAWhjL3P1psUGXLxPhkETm3T
mD3BID8ZXZrvuDTjWvOXWqzvy1e6nrfdm4Ev6Mp1Frp+Ayv34zQ12xUbHXgE2rmc
8SJ17wfyf9SLZuL6laMeFlUESL/zMAwCsOzWhaNz2nUs5oFCPgIZM44cgW5dpVIx
uaER/Fai77vFQdqJCUn/aRWNxgIB2/Vz6mQcgtm3Cp1PlK3gHyyynqj8IqHvq/n4
HYdp5+MQGA0OSsB8lb3WGVorMvTPiice7Qxmg3FEEWfpNLT8BVLP19hFDLGZ7f/L
0SJU5hTWmV5UQdZxl2JMpW16wqd0Dm0T4Gkj5S24nJXBc7E1CkkAL4MembOaSknQ
ZpD35Z+/TKxQS1TuIFd7gaKFwQSAomb5gL7vl1UST3BHunXsJKsv+jRSeoBe9sbt
rlEAxwAPlh3RE4pXxsRJzHe1//358YANBNFJBpnzQ960+wlpEmrhHX6J9LQ1Z8C1
qxlYowLJS0rgtkF9+hMIXj7FI+nTaWLnfdoiqvHyYtLEBtMeZaQ48eIU+63AtSmt
AurguI1ljPVkAN8qWyyDr3DBSbNDJTXrRR5C0D1cIEKmM+HqojaYoCW0VBD30wvs
j7+uV86lBZf6qc1ebgRsKN1VTJfgZSs7Enr4oQVXjj/eajjlRr+b6GZkoQvPx+T1
PWyQKRuRaQ8qdLyjvzrh7Xqn6XKRWeB1lhlaYbgiKs+tF3E31AR6XYA0ge/Ly7WN
Oiz4M1mb98/bc8+/Vi7DaEETK4dobZoXcofYWa1njew+fp17M0+R+F+DKE7IBBU9
hpHKPK8FkIX4CURiR3gy9RHNGx4faH25X0nQLfzkr+Ng/xlcpLa/kxWU3n2SCSbe
fmSH4GkRkflD8aKzDFvBLHDEcWQud1PQ/BzBSj6BB4BavsJH47IbKD7DPYIX4ffv
Y3fWfQKdVzizYEqleq+vRAeDE3S26o4uNoH3JfMr2KBk5W0bJ7bmRVjYpBE1w/Db
tQSVQgtsxAGgAYB3+co17i2PCcF/wPcZOcss0oW3cm395Kp+bN9It1T3B3g0j6Eu
3b2rlx6sPNNUEDMQNR3/H1PQqbA+4FF1jyUhbgW9NBH8dOvoRLrSw5zpGjVBCnZY
a242as8LwrHZ05X8nxOvQBz/0xJClaz2D0hujedhCgKYqAiMured2kydn44VvsmE
nu+Lvt2Mrzm0A4BNY+ebbWYSuSIWxpjsu3p6du97WUads9zd6uygFEp5s+nmlUC6
ZQkYRNOLzCSpP9x2qMZJf2W+nezc8rbb60kbDYN0nAnI28IGBXn8/BOUG5+vJ1FI
67HcRTELRHdEKBSD7fGUuRP6ShJgt7EG1wZaF3P33GwbD8JgTBzpQJftZGZytDsh
K/M1Lza3KQw1c/9o0zFwBQR8le+sP4y19suYH9N3wltUiIh+eZNZS+4/9yfkfMUU
e627SQDvJSi5K5E+xTIXd94HB1zbw6u9SGtsz2AxgxZHLv81YPd592VPggCsGU5f
/ymU75VivRsWZjBsTIQM4e1EcIWgHfKGGAdX3jrJ+GNOpZ46PIPNM0g5eJ5qFwo6
OYMc9GfR5zW8rLud4qpdVGC4VJLYOAexpVulZ6sZkFg6ma6w9c+lH7Mx4B0FzXHY
a9FQu5f4jhg5Ro4mJvE1EQ5qa21xp9yH1svA5yjjNXCoew4KYkE6SmOhkDp+inJK
2ZDpuQ4/2qkXdTYCLgK47ZC2pDs0G4enW+QEWKtP2daH0Yqqmws9GQ6AJqBH/0wU
bJk0t26sv4veDF88OTnz56NW4FGf2L8ACzJQndeJlO93+x+sbEvqUt+EM0ojZwrP
GTNyr+h4dLvItktaZAos+c2hhIs2nGe+GWsSuK3kCjcxIZWxaW/oo5ZepudSgRf7
P5GMMdlMTeyVr42NHlJU5Ucqa95HYiPB1OSG1/vSb1/WbXnkXeLS8npYXSTHMTvJ
6P50YeoIGt5WsmZ1qhnrCkwBfz2+h0AZ/ohXFHziGp7FJwS38i5nNUiahaMvY8eT
mprIlKqNN34h3VSwT3vmtpyQT0VTKmvHGAvQM7v50ji4IAQyRlgXXVWrLDez84Ut
H1OQ1kSd7/2QhEYWy+fb9f+12TdG7SHHObVVn+LS6X8daw9+oQlrDItZLDPrk1dz
GOy1GPzASbXvZUp2J5GdWZP4+O30PJ+8GMr1OL66YktZ5ts35JMV2zM4GqIHHcy+
7MSrxuwpUN3E9u+UWkdVxE11r651YqogGVEbsFNt0/buGDBNIZtoIq6+d0w00Cqc
BbiMYdQoLOtvf5ACJGNPal7IinLSHVZPKYBLkQXMygqv/XWOCGQaUJHEAwVpGoLO
Xn46O1PvlPdVpuPsWsvcOLQn44APIZa+7RPRmfC71rzXg+AHkKml4rk/Evt7UV/d
cVxttCZuyN89/faRY5SqjkJgQLQwvP7CObVkvAgmR8+O05htX1++8g4rn5G2BPGB
17JMTbGCVZf0xl50vz3A5QUlT81R7J9H1ayPuSWIFy7f5+VN8Dsn3TaNUhVsUY7p
JissLxwLaqO7QZVegNkXyj/C63rmLMhYEekpPfBmOzKJcD94nhtGODn5eBGcZOjQ
81EiFB33Ix36EWQvHKbKiapUdd4Lo5EFT19RTyO0JIa1vOTDeesidhvYsvfAuA8a
cU8gWx6UOY8l1wRiRGlWxivZTkcLTwOwT2FwkYrrWEmDXEhk5X3WyXKUTyQnt14E
6GH3AEOik/q3PsdPfRQ08NtCcgsCk7IuEKA6kJxgs0ZRFBZXp/1pkkQpKw8UFCYZ
z1BtjJWcqNpCPDrrI7Ae3f8SmJQFz8682JHEXOMzxjiiv5jMF6odRU1aJ27S2zhD
oYHhHkLm4wp3qIaJQfrAJuUrf7sUiIv4evd5o5wFee3mrhhbF/xWiWa/zBhU8y4k
UH0kWSxbf5xeXIbBJ8hsw0tama9fbX5ZBF1yvnoVJYtsDimwLXyXxZHp2OfJwwD6
nyhstjTQbjXWnGS38kX9GoZaH89JUOijvLeqs9QlFf81WsfSqTjsAIJkMYxP50Bl
3IBNHZFDUWhD/vl+A0uF6KFtmf9urDGOz63pm8EMBedOPjPU9friR7flp5AW1hTM
3o+qYKia6X0OlqG9iv79GaA/kbT8VqXI93EQv+jM6aPdIwYPfYC4hhjGSUQMeN1l
VIFyUySACCj7C6yYWbHEws255o79Lpg6NfHN2GNSzcCve+xJHtkfUCwxclJ0r1KH
GKn61jylrLKvTw0c6lvMwEIuVw4YSPvlSZ8YaUGv1kV+5cM5Nfb7KUCeFroIJqUQ
oh3hIj3I5vYiNUFmCiVS6fS6YO88l+VvkMrPcuHJ6dCUD91ruDnXfBsAHoZ3YKK1
kVWt7QRYP8KGHCNcVD+bDYIow0IUx1mhuqDbacvR3hAS9A4g0FCIzGwZiriz9gzz
QxXn325xMrc+8yPHe7E/WuUPlNzxWvZlYPXJO505OX/ViJUOZp+VdpHN/y7pvMuT
TcMSmDrb001tTHdfnNq8h6z4L/WP6E1DyazSfnIi99N8TFGnNOonVIh8lvXhYVCw
r3NDJYk+fSb1fZCXEyXI5Iuhg2FwXscED9j5noWwB96qnGocK9+1QngUmGXp+9p3
kbNrnaLPNThI8VwOs1GfGaY33LcHEw07F21J5DtBG3lAe0YjJLMfetrqYb/319wz
AiWZRMgFijFl3BZ7/ILBQ07cCdDkT4qNF47tSPwi6+URXDKprp7ymoLKZVhUYK6x
Wx7ynVqahsiMiZeWnIHZoBnQo85RAn1UHP2GlHzEEL/D+aBN7+Z374GxbPATiurU
CmiUByNafc0uqKFVQCg2zBUZHsZ+YpUifOEQvscP26bKo4cc3cXwXIxA8D4Nmhvh
UGtAZbrO+H30EQFNZHz944UAvIKsQ5yMZAAHT6aXF7f4i/emyy2jSh0jadNWkyo3
vce5gJk2LYDT0Q4SPHsgB8FkaQ9LgLmGov6SvYxqD13TdReb5Lf3D44S1D4QCSM5
hKno1mCECRCWo0V0gIyOWa6nY2KgYstx4WBmymRSbT3E5s0G4eY5H/bBSWORsLf6
cl/MM3xyRCA3WhgWXuylyjPv16awh/NRoXd1g4GxhgexXyMvv4dypEicQjV6VIHg
paZ9ph7ArUVNHspsKUyaIsD1lieefARZYPZOkcRAnYOeOPGFFJi52fB7HtCKSKF6
zW/WyyIo9wrGL7CJOAt3s7WRvr68G1kKIqGkV7e6OmR6MuVsc6TZQlQPe9kzNvRU
7oobnyEEh/wdOYncbMf6pRyKfRRbDdQnVE1mHiBmjjAtFfUfHSqkbgfyXyWdx362
KWwkO1PiY+qr4W3qDxfRbWY9wRmW4uXJBiRSBLUmeV/mCdiVeNKo7hCvpEKxI7uG
p6JHqNekOqzB37nP6DsmilqkbrUYYIzIopx5ejCdoMTIHTdc1bKFuQ3V2y1pfQlA
CVNuuwFO5uGUKWlKFEYM49fKaJgCcVELQQjH9dYNuFmrt9Fzds9MI+ZHRFdPfvLf
Jkw2UFW8NLt91IRnuZE3Ps6Zo84lOG1v1myV1P3RvRRJwV5SKyQPMKju5RP3hLGJ
j5k+NLum59vbF20WJmVycj+bwHbGYgcA2+GXcJuenmhooFs0Gfoc/J+ooHgM8nGy
6evR3IGWddS+oH1+qCaOi2VHGJwycw9053cgdybVNyt3ocXFypszinsSvbFrPjbH
mrr9jG4mtZofTvEneUmDe/BUN98uxxoM1zLQnxhsQqUkFiSyS1rV9TzC42hmLHIr
ByMS8DrXY432yhoQtGzrDwxfc+t34oJxG6Sb/Ms3wsJshZIixkuZL2Urab96iLCp
6TdWW+nd5HQriXqNPHAYGVoyE5LZa7RgMHhhgw+ArM+P3SqZnOu8FYI14tbyLHzW
wA3Zb+bov9SS1uER1CyZDDzKcJdkcNNsgxn0twKy2JmpYZQk6FLWMrBSiDcf0qwD
oegndPsUe/diL82reL02vhG95X9cRkFb2k7wFlzk5sWGJEt/7j/orTGKtTIGto+T
c0PLh/SY+6Ga0Msn/WDPk30BaegTj51XUw4YPEKkIauMDNZNKS+ytnLsjNSdObD1
Lsc+VrZ8QkxgjBaGj3vQzYvmiZ450tdlLxvVJTWcWpoNTTGqae0eLHhL7Q/UtNma
cxmlr00My+7V9P90L1T9whTp9BTd/Nd/3cAbCDM+71Go0IMSfX4zE/P8qqy0OEsV
WYG/mIEPn3TY4jlKGd81mTp/7ON9LMQCbW8x2bSaRr6tQBEnnjGRuqq/V5V4CMuA
G1Vx7dRttlhDBOh4usTW9gXMMzg8k1+UxbAnacBMdl5EAMVyMyF43waR6QqUvzU/
b90HnD6RPFXGY40PUNrOiSauqB5RD7LyrJbBl4cd+sMzcC+zZT++abMvmneBub1B
B0BLGFO3vyKzdEju+mfUEFapGDTkany7Aq9FcOB5lVID/sxvfDnkBcIBqh+IGMzP
a2G1UROKHOs9+vL1FHql8/rYxR9IvnrUTAah8zCpd6aQnGW2TKCI4ukkJs5U2b2y
TY2xgnRYcH6f7ocE3Y8IszuFOQFslB3XdC02Oe91y3gDsZiW5lvA0Wqa08dpGTBV
hcuhunJfQKteciYCMFMwFVzXH9g9uI5S9AUbGoC3Ftbvzeia/TnYYAE8YDkDf5tH
qnQ0FT4mR+pGAesMHnN9aasnkC6OzhHDlqUw9vOhxsXt6T1ubADGsUZZbMGgQDqK
YjS6NZQE8xdp9TIt0b5GPoiBqOAMOBDzFqloTOuCN1lYIl8Mo+vMHxWRwBlaTgpB
fcuWWbduCsf1EumKRZzdSAE1ijpxDqIhnMgAONkZyHWZypUU9u3zAoL79jV8O9dj
oAZel1s+4RENRmffo2GNJvK5vAS62nfLp3+lBPA1zZ14ioFK2Kp3+JkGXDkCfar3
cqeARcPnWJvH829a6jdFbWRaGYnFzMv5xA/3DmWbKITfaHVKbty2AYb25CZuPj1z
wUTEedM+geucQZaXGSyszA8KL2KUr62MafSw9yeJiMvrcE5nA+JOK+ik769d6NA5
GvpCRFAt/sMZXosb3dCOmbODco/5aQoVGJfweGktoG9FJbKsbwzkn1lrQez9NICr
yA4pH/YSLgAa/DSEUzGVQChq0X+nOeSfKFsIAGQEW9FjHye1ZqCN+9ooP94xjm+k
nq1wCO2znCj9gO4ih7SVJYoA1p661WrvlsKjYPZ+ffdE37jhtaKxVMGPq/+qrRAm
On4vwH63EL9QzxU5Qe6XXCC1SvRlCSZWhjdWGhN69VFbvftNfVuHjAo1fgHzzJ7y
Np5tXXjUu+Qx3dQ7mIATwxj2zd17iZ2n+iVxj52+SVcixgi2AK5s1akSkbYSm9AO
GkTshsDwr9IkPIX+EptQJNg8v8d8TwBlvH0lPIwZSdFIGwYWa7MaYZiFD91j20Pg
eG95Pyx+zhygwd8bnzP4RlqCwTyYz9ltsYiuMp4mDSq5SdaUfWDKkPChZjTEHGHO
ZJ9V7kiIhbhArZsjXaV18GvzibltQ2imGrYbC+NsKuCl1h/MMmLtL4/RuAZb+5VH
w6xAguup83jWBl60TsTwNBiFGShoQ7ll29KTlpF2bUaWiVVVsRwrZu9mQs/ZvqYQ
VUjoFDbdrVzQJXzJRWpWSQgZd9k97x1Uv6liodrNYL8XoERYWrjCZ4Q6CEOnC9ip
sajngc2Eh63fTQWsG+HRIpZfbx0PyoRwEfce/A595yI/r9j0Tp0cM4m3kzPz9nJD
dkWwoYUN+VZcuBx+3YUIO6WTQ5+EztK8RUvr0oIO12lB4nFoeO9yyvtwiwhyVvHW
o2cyz0Dz5VLVZ3avdD89NyYDzsI4CECQJ0wDXjhNtezARhWExP64/jJXlDY/nW3T
skTUPlovf2XlbXburQsYQrNJCtCywtXyUkyWE/2GRT1R5nYGzVkdI7eVTCqSyJYK
Vij7EcNydiXHuHhLZFzqi1cVBW0/n0PySxpKLT4BzMx4lXgLMQVKH6/aWFeS9nZk
U7g4UV/3U58OFQmcEVLSdHWBeajOPE2+9SbnJnofum3ZrSObUJ5DCkRwf6dueS3L
MAilS5OGmcvNsPaK0jipf/jjMvkvy3F4cpEGiH8e55nyUpqcIZ6LdPFiLdLz0jx2
OctdL//hZS1YyuUu1Yc4pwV6YcJSmZFc8El/VXoFZlDZ9vDAiqVpLPQFr2QXMMSw
PijwWzMtHEd6QcKWd6kbl7WiWV6b1NG4ogzwy8gOdeoduV9KsJ77TWJ5GaIidwo3
LfrfdX/GxyH/Jk0nH6MRCedhDrH/oyFWA0hKE6dXVK3NfNKX81iY+Cgns9Ggo9oD
pFHk99gSTxdIJ+ElDGZGnYlyl/W98MAaHPcd2GoQH3ltkq8xjRPonIfX0hjitEyo
WIfsaJDvTPUbE3oI/k496JKHG8/V2MB5LuzgG/oMK5Bcm1tk7tjo0RMKivEUA3Eh
D4R9x3P9VUXPYkTKQ4Th57LMIlSd7ADWeKsenSBl1Gmpho85b9nk1fHEjdmH8g2A
tJomIkfEBnVnagSvz3gOm7JhJPdZxDmHBk6pbwMkxL43ZGa1kqrfzAbQHwDcq0p8
SQw+axgc8fvGui0WrHz0F0KcETXnTYhfcyJdJnlrvhnDePyaMLFp3aSNtVFfHATN
83FWw67yYVPcs3DQ3620Nbgi6q+p2akNT/0279nZ67Hfw+f34TMqB34x/mSa5+QP
AyapfU55KwD4RJRBxTf38t4Ld1957XHVd15UvJNdn3jrORJAmCYXvajIT0gmmi7J
STY4ceU2JkCHsDzzG6Z0kIvCSM3sO5tgvCa76ZIxgzpL2S3e35CmBqQor9sbWQB3
e6alZAzyW4gC2hj9NO6/S+IrYq+J+3h3m3l7nObXkB2vYwwp4nOPOYWiHrpGAJoN
HRHySUijZkmU126QZSrBKyMgmoj7XaHGI0yu1ZgX1jCYklRXqxJ6RBfFX7+oWs2m
KbUtF54/p3hTraxtoatPmwtVXPw7zGKb+IM1Emi833BqreWb+EPqUegj0ccQbG4V
C2KtTp4nQgD2NnxP8558pEHWKafVoF4qMshgw9JZ+C53CBmHz429I8q4j/+mCIQj
gdLEMNwjXMvnl28NjiSywe9Qm8O/LSfrP1H3hLUgELRWfKb5MwIk2mKre09cpRBp
767+R5Ox/RMYpYkMplNkYgQ1T5dVnK24ZAGl6g8jpPhZ+56zGfVb8HdNwLgEJEBq
8+Z+G+qaKWPpRTTFw/uRJIGP1fBJFZ8VR/4hBWWBbSPamx6QjYCFO74bTPgXywId
V1My04Z3jWdYahY15r4N9Si59UKy7LIN0U7pvtVpSK/ZUBai0J9TArKD7CBtv5mh
QVBXPtJ+UpZeAnr/eIKa+ElyilCZtXfjG7EzNwygL7jVB/7Yy1VGL/0YJKANQhpf
jqItPSlJOB7G8mwrACWPwYOGgsnOO3lP735bLsxiEDPNmYKmbYVfsWifyav7Tzv9
zK9fz7DOIfWbH2e2Xz2XSl8oCQwv2p0I0syPMK3UfNwuyU+9U3IDT0tNbhbQlxAg
9pPIk9la1eK98S9WgLV1JJTooobXr0uKvA6UBBS+fH5zVF4U/6xo71seitxGZjUj
+SWC7qisSbrWj5A4DxMbuR7d/eMN1+VYfarRQoGFzzipTq9qXKDcx9RDKfw1vy3V
DE+5rStW566SfxOfGyBZPg9l4hc6+Imi0gzv84TeteD6eFn1nkAFDsZOUZm0BY2Z
B7EyH4NGkqeaHNEKv7QVBLX3Lfk5JzY29Suw86iv1QX9Bm+hQpwc9BrT+NOA5aYM
RENGzRTLkUeChuERwAGoz+k9P68A9ezVLy5lm1i0GefT2RwmIrTH19UCwdBm7IW+
dbVPAZTorGaYNHBMfC33uiCFFQTc3ClR9scw3UOHzOJGLIlW1Ae6jG0tyRtmiP35
8jhLFEnVd+nb+oqfjCbwF9xkh5eTsWDOHZFO7A5uwXXiSkCw1nb6K/vy7t6xy1Ve
0P3TrsokkD+teOkWQ0LaCS21UsGAKBV5xxtWIlznSRMf71CbOJYCwexHi/LdaAU9
9mzygJaFvE/rp3qnRhVx1cz8bYjCnZvuRv3i86v1VjTsC84EWUETUsGyIK0sf8Or
PicYtwnRVnVoCTI8CaFf90uE98X7jOrsgAXbcW0CAmKAOVzWDm0yDTBYik6lH6dy
BhQS7oeOD1e2rFk+3yD5qelzdMpUH3ZwMH9t/tOgFMqU2Z6G80JkQDMst+89jukr
cvqOdCQmgtxI3Jkzi2drI5J4z9Cf1B1GV7fKSUJsCxD06gqnvUDHzZtOhlvwaaIE
VfSAKVb7U+J1dxq1HSktgLgxwuaI7B+K3jOgPwgxQgkzAP7MB5j2XXrZ5P43lePE
81mvi7JfGnRINb4pqC/ahZUcKkBgA/vn+MtAU0CCUBYLehhEPiddeshGHi0bcNS5
+v1ARRgRyYEtgKf0PBGvcuec/eKwBuFD7EuWri817LrXqJSsSY4dd9QGnzcu2ucs
czHzWZe2/ZMpUwhWeGCucXI6fjzNpAMI7yjFA6/W7AMRfFIJ6H+Lv7X5OVCHJB9b
xc61Z9FqYYW+lKfEyb6xO5j+tVEj6vg6onwW8WuK8mLh5FcjAbxyUuBy3QRfhXjO
yKoADpMhyvy0ZdjU3tM5N1VwxAJ3vDrvz5t7Xe/5zGK8GoAvWVP1lkLXLQUbtKCV
IzvvvuhUo5v34drLhZeAcsXGsLdhDLrP0c2FK8zoqSsY78PDEW/oIAmSkZjxDRGe
H7M8NGQuxKa7eQte7fTk7k0gVLU6AMw3eRCjxgUSeYcSHihYcs5VdqQi9Y+L/z2i
zt+U3wB7r197UMZh/gWgqHhcRUc8+wXCYOjAweqO/FIndGkpnkNMtVomqLSNAVqe
a6auE09tIhKHYUiz3UwmIpGC1nPClGoBTJx2X/mBqNBk7PHFckKcFb3M2ZN8cY7b
By6AqCm+F6AUKwm9+2uukuUmITEQlOXojqFMiR6TZYe8UZgaUdGofKxb7vEFPKxO
FVS7clHVPyKFq+zzU6ajW1t9TY/rNHzAz4P7WltLt/IvtC4mjgdmZxUEnVBb7uCg
E7tIMUoTRtQsipv55svDI++YDtc4HzPjjlH7i0V0PbVgoa5EXBptwXy+QQEpCxdi
oqFMUOPXMsimTW9bGSKVClg1ov9fBoZhtTHrrdo2kB/ca1iFGjofDZ9NOjBVoch8
9StQ35QUsov43jugrvShSthBYnpB3YybvLtdq1Ta1wGkuzuBmKZKTp0nf4/3XS1j
9b0cYIGzZmktWyTHEWk3MHSVZBlvddFHAKy51QS5aX7TLzXpcfHcY7+6xySYZ6P5
NNI2agHVV+QxzguMHDKYJFX4/0j1qxz1MX3fbK1w8guPXnFNd9Px52UUXB6GL7dn
6pLyMr0UUyD+fMISd35RbyigAJuoRTSKUy0SStITrKnLLoU3hl6WDnR98LlFWJFk
kX3K8MW8JNtxMWinyMNHX6gGqX0o88FLzN5uBXbCLVXmK1e+011tzgvTZMc13moD
tCzR9sLap8Fh7JelexXT5BJ7ehwUU2zSJD36V/KQPMbvPNnLaSJLPz26Tv4EnBsI
YRboeWSBQd9LBCXxlefQRw9+U7qiYShpAA/5mvLpGJe58U1pdFSYw53VQa8t8W73
ShjiBRTdlD2FXg4opDK6bVd6mc175feqG1WHPK0nbgx9riZbBco5FBNQNjmkTiXS
ab8FUD/nk6Nb2/cFaL866MHHypLkignZXkvkm3HocxsxYWxlBD281ABm4ludI2C2
NJaWZCeRMeMxpz21OiodsZbbispbJPK9lPuE2MN9O56/srCAWkxODaV+fbEWb9Xh
PvEBCaZpSyqQ3lYm4cmZFyyzNBdgaUgn6MvW2YkipXbC+rNrf6o3GeLab/P9WEq3
rDNMtEP1LF6BAgL7gNiwemeQc7Dqo/rLX/cdrVwrlhAxR3tCWzhuGTqQrqMle/eq
0erH4g/FvEuHiY/VdENebHrWPs9wVm6RU3yxDzvXeWZ4BWQn5RfEWMccTRmhZbni
2e5hAHwvoRR1KPt6PC9Fe5LXGh8KVgu+FyvLsNNwuZNlc9BTAXnkLTOW/2TR4GHo
+jrAJI5pvUvT47PaC6KLzrpz+fXQZWq7QwEtZSKg5HWqI7eIxccdpekMVT7ZFzrA
L7x7d2BNzUUWjeliZBo2gjieAZ+VpqwyvDmXisbnfnry1gvl/dicX7m0OTbAfcws
aL1InF8hSmcOThB/wptCnNQDQhqgh/RyO3yw+rPlRWBkHZxa5OvXOjuIkLVmln/E
BZUC5gzhikij/r1q15EomX0lHFNP5h8uetuKwAQT5nnyugYSVKWlHi0NreVn0/rA
uDrjztwnNPvxj2I6bF87Kn1aG4hjBffimmqNXei6AKux3D8U1BfrxBnItm51v6Ua
6p+KxWCerBXvvUtAq1TXuYZ8vggsgktAh/Q+ug5RLopzkShnNkk4KFHf+bSii+na
eE9KNrhRyS7pZsmKUqUYtZtqGT2OkQuKqCab9A/PS36sCtzFUaeVYGDaLPApdPQr
Sg6K+RTck6na/IucN9JuFJA91dayp2MHG69QBbLKulk+MDzewtKXLONfuguKbM7N
IlQou32N+6RqTMUskPYOtWb9q4/WO8loEVwo6dI4S4oC9lgvTmWuz90KmlAZEu0V
4vRBErFTrsNPU0NmhfL7dDyD23GEyc/I8xIVznFUk1gXAQRh3+b3Alvji9/P/pWS
qocTzHP1Gkp+7nSqdyKo/92ulILGnPKOUKuEj+tN6AEKxFpsXXd/kxc4unZkC/jH
+u5/fxfJh6cguH7q/uRAVXT9eiaWmtYDDPOn8oHMPOt1bpE4nYqHJK7AhgKmeU1e
Qgt3LqC3gMihsR63mp6fc5BMyb1wYTMPK4tX/lG4paioG4pUZD7omwvUVi00bjV6
VodesEIcJ0VeYt+U0dS1i589XMuS/37FzV583FZ7Uu+KA86fohWQnwnc5VZUHwHZ
rkMm7nTfvILhXwW29YSRAzXNqxOgLQ7Pozi5a9aQ+hc3CN58Uuee1wf7KlC1pmhN
h/+cmX2YF9VQanFlJUdwvrXlD+Z0P8o65bcYpa+SbKrjX6ftkuvlypL7zBFcLWeG
fmraMDeIqHXxpTvOzMi4cQluTBK7ICARCQJ/bcieNDfzXXD2v+4vkRjaloY5LHa7
+/oA+/2UWOcyN6TMMYoGBJmKAydVBLucAI9qMJEpGZycIuBpm+pSKr1Hw22QkpH+
qvJ9cdCyBJidiY1g+qMUuFT90Ak2MoMheey5bah5iShnRWNnglybnib7nfObISvH
f8xURZp8UpYRPvrSzu+yYlS1uPh6byCs9eZQeJWaB0Up4DhVb4i231gEvGrgXvB8
ydImQ4hsJ5bg1trUBLEO7J7nuAGkNb8thwQBSj0s8s2PP9PgWzXbMcsyNMuurIGZ
2dEzMSitYs0zVgkwB81mOgzWZ4eWz+VYVil76rCQNLjiCnO07iZiYajCrmUsTl7o
Er5RyBvrm6I/3txZhvo6QPu14g1pAZsafxJfGO+9jqxszzqMwMCurwfaRBedYasH
t4URo8L/oUavQYSB34ViKFdBVEyGdfQ5+uFfVoLUd5YzPh4/Eme6YM3oQ2lp7D1l
+Wexb8Bb8D/+omP5SKD8KEsaMIhEDwO2VsUqf3NPP9z6BtMUZTFf/lnqKVis1xs1
/Aa6r2kPgi/0o9xjGfNigHmQoiuvJN4wzhaQ6qTFmzzkiL1hctHrFFP0Z8EhFHwp
cWXtAD9sRrfQu2Ih9hdsDBYbKyb1FXOvVhX5eKyHXBusia/doHdlsMHrFFLW0nqa
0iSTTSY6HmEUXXylXnNTPXz7g7Ks1AyqoCAwCBOY9pkekl1x51v/W+4COeqcXpme
7Nn9xG+UDEXVEkGV7qEnpCoQlYVMVnnSxNy2HgxIQUgYCdOFN4rTNQkq6GYO84B3
cMkF0MV0yuSKYJpPvJeS+aQgkDYNn6oVSYuBg8EznuW51m42rsc1e2AXbylrA+za
bIItjCQVnnbI0KCxaah44Awn909JxNxzv0QPLD0fby8GivgOzhvP8raWJrlptOb/
7ysvgrxQpP2G2Gdw/daWC/UQ/NnJVS6u97GqGEBRM/UKC+iQTDCxkZ8hKJ4l0inf
xYrqEL3MpeVXqoXp2r2M6Y38uyJBBnBaqiWsJoHukfbXjIfujiz7pU3AbHwvrdc/
NFDMa2aaLlx1qoNXwXru7sVp9P3xST0Vyk/q3+Eyiagwqz5nmmr1KdCjmLVyzw9b
jx5sMGLjLpgUuuFu3FoIpZiUMbbBCqxwABZMIDA82p3bqnMPSw0mTms2shMYzvqF
j7SFZ+ToNFCC43tNqcdgx0P9cdGQt+KG2l0RlUiAS+dhtbRTaLaO1Bw8TtBusqXa
vYFT8f++yOEUwcQzpyEqhH4MGNEC1c2PSivkSuT7bbyZG9gIb82nxJfazPYgtvN2
l9gf3SXoQ10uA87YlI24/E/XOecEy4Sst4aApB2DlrO1Cy7mHpJctDVt3yVgpGzM
sF04pg7mJehqQYGaV7BxEn1VhCgmiUfy0LcdKHFUGBgcrmRxqjcijXQ9W0IfihOa
w6oM1uZw0kQoe+9llTs7GeyBXrefrsPm6qffH813vRVniDNy8ZLUBd87AvpW909f
WCUW/seFs8hqraQyxnfuN0sscS4+0CAuwpS0HuRfthkruAsij3HG39DSaV4dkTgT
x1w234E6cMPdUFQxVqUwtuc8Zjk89D362sBQ7E4YPQrXhrm855LkzfQHJIZV/c9n
pI6kjZmmVUVctXY5sRdghKO0I+R4U1VZVJki36hjeyw3Ge9ze6Bc8cIwoGXg+1Eh
SLHfwBvYzROEzbnDbMoGIqFskSP6zjKfNx/O9AifhFsDE5iAjUa9zb//cAqOFS0+
oXXgW/nLYU6CTNAgZZLAyqq3Vq6uXPy7N/BnCfC26ryuVqUs38/rtobk/wvo2ene
iZUBg3IM3gBcEZT/Ans+9KsAW8NaI0I0qys7SMQSMKlYeGSDBF+YMOBXQ7ylsuZ5
JRFYEs2lbtvIqW9K/AAQeieewoG+NcTidqXaymhJoGIHxczNYnje0yfaSzutbC3g
qQLB8+WHXp7E803mPYu2nINXsCsp1UR41ouQHk8hziBA0pci5c1EWi942sAYTHZw
SVNVKTKddO6WR+HY8q23p12bgALTqj4lOkVL7WRLP3dSj2ntY4Qg2Zkh/ooARUz7
rkl6HlPeOcg31Irt06ihuKE1VT6gxtjkc15SB/fvl/Mw/XwvyNvFRh4ty/deL+Gi
JNp6rV2+NzSu0g+jOu1RkSZrvsQG/P57wkt9oVBG9XgjmdTUTR5X/UTE/hxoIhT+
T87f8e/f5NvRHNmTX3G4TjxINsDg/TFp34tqbl9+hzfNeb8Bv+aJLiKP8Wuy37yz
e6m3RwJpdZK499OAeFT7fIykdA9y9IlSt3pch+hcS33jkT3rPqdDE/V1kOF/SvZr
PqYcVhbkgzCN724ex/OtSdMpHJNXs9yJJ85bY0d7qKuep9ASEhylbGQmuJKNFoJz
Uni+lM2DoiEtHC8VBCnPJcGsQtSc9SEiAs2gcPEbgCpzkjCtv8WRQXjHqw72uje3
YU/sZH2WZDYLOPmlQ3qq2HuSVwEXxp/nI4XX3ghb1wi3bEY7cFcIYe1XlJQ1Nqur
NIRN4xcw4zVssF5WqQHO23qaSmbs8aiO8DDr/OiRH5+Wz6Gw+aiiYFevMpKY/FOa
LjYFN8gYH2gYb3TdQVjLBs/BHscZ7rrAZ3+f5bc67Ou5XjParUQBJWawbkONVfxb
6fZQSR/IfD1g8uBoGsd1ejoDSirKP5mRQ0pM1JzKo/xiMuAPKjxVOcJ1eCuFWXSO
pNooChbVhwJLEfjmtxryKcjZ3LKcpC0jL1n+9kXRwdoKaoLoPMSehGcmtkkvCrxc
4vIpLh3bWoeZYbKBeMfRNX/EgvlUoyjp8b/9/UlUu15Vm/+yMEVdxpnSVytvXmaZ
Wv7sYIFpWxdkJeGCXrhOERPse1842La4cjx7Yx7mr5zBO6dwCfM2QPbwV7q5gnGE
SpEAPce6Vhs6DmajycAaAOF9EJ4PAg5hVfTPc2RAqd9Vkl+uksE6YdYvKG2CiUWu
Nj1/bk3+Ip3GgdGaR8U9bUtPdmEgKF/0f/gVmqArW3y6/p+sYqXsxyWZnmV1ptfW
0UZjwBCIHZQEBXQF6dMAbRB8Z3zEUyUM5PE+wS+dPs8LqIn8neHIS3Tau2YtiQV3
X60Otyf7bl8XlMtcPpqSui9O9FFxNjNgkMPEM30y1DrBVdwEjZHLMdCZQlvVILz0
BWyJ3sxYCo+5lFauANFX6j3uk8KRQal4alfssvkWSFokPlsXhf77XZ0NXKF1E/8S
a/go0BN6astMI9pUa/RwNcUwMJRcObl1KyUqR/EOWkc3pTaG2RC+JI6N+nSzVnqo
C3GaaX0AaazI/r3ywKRXHpT5gfmbnX6xU6IhPHCfdoVqJovRy/71Fy+2hGcsvuTu
DY1bwJX4RJkL/JtfWOa+eYMb90aBm4ByDrpdHXFYCVQe90fMd/DUIqZ2oKSRzCNN
5BLhnMasgdpQv86ySYfjDnlEsDBgV57Qque5dHpJO5UCIHeFfI8LnAVuff7fgqJN
ipI+NTrlj8rGhLjS5SFZw11GjJR8rgLNRixal2iOYv4YdOHfZxpxgf6wh5NCFoxh
YkXpeDnUv4siZYHm7lOuDYFhoYD+5beJ+lbD2vYIhSqSJJGRodyxx8pT1bVtTbzh
mJYd8i82TzIA3gyMiPtc9IqyO1moUXb/McmxEsmx8pXr3Mk/ie+FSxoviao9GiYI
RugqW8I0pt5hQUuWS7Kq51Hkap/r821Uu/AGFAHgBuAYK+XVpUxFaranKB/Q9z8G
5oQ/oQGtZtx2HPW9WEcPavsALp/V3X+VF55hQmr9EFeq1auljCv42xKE7QhAKPl7
W24BTW/VMXmCmqTo+HxpBpNd5y+/sMsab1h4F1pbs3UkBhFycpOMMxKPrj6e9kxn
JHaVX5Y1Ee2O/p0oQBR6RGdNeTFSpR9hiY/4g7gIhSlIpka4tH2KSW+TQ5oyP58E
lNL/t9xju4AIwuGMn1oqpU/Qt4pkc7h4oyIHi+rUdDqIxbNyVRcirylOfCQvVlXj
VHdT0pa3mCYAjHMXuUaE9sXAlSvr1ogC0JYfzjzlFh5N2Y5HxVqxofoZi7mfgnjr
L2Ma4veFKrkPNqkTEMSoXsVC2jBGAsNU8fNso49U3UKtxGQHgopx2GPF81Z/Geix
YDvOr8TyjgZp060ZTwJdgn9n/07TEdUG0koCnwENoS4c2dyIvQfht/7Bwb6njzjh
trD6vIgKFG+OZnTmvNDiw8qgcx5DTTAjIEk/RQ/lAh9ntRGTUawf562pHXC6sNqQ
7M/UC9NEZLT7IebZHTkpZHcu1k7iwFhq8n3vKolQo4REiSP4UZ5pshLikVmFGVF0
esUJIq1kFG5PjjeJlT9/lDDT7giQm+U9HVrH3pWDI5AlXyGz3GFPQTWvZhfLRUrL
6ViRShhYntP6NrYx6SCbnhdo8Tvv6JOdXLExg2M2pUKCc5qxGLvxa4+sfba8LPkR
n6YR5QMsDwciMHdXvJiFAsMsVLxxaktBjitGJOaaIKz6cIf/O1hdDSHcLmu56spg
GXlKWNLadu81zvP+RZWY0hcdjswE36etH3psXhmMQkztbsk0NE3vzjVIFdlSXctM
gNzIB69aFcY+6+mpprtyMlIp75h7lPjpgVSHjo4ooIVSPDhSun0nx4r7aW3Wu74l
0wRXYAP9SgAjDZZLLgft1BselCUjO0+bXk5xmCkpS6WuLVuN3OE78xClp3+2MoyF
R6oiz3djAD4aDgw60iJwMvd2CETWzbOf5bD7Bvs2tCPZKtsEjM6lpFRssvsrQuzU
jRvG+oGjEXbTNurZJAZLWqkfG8vHMPGc3TVN2cV9IEb5cFEYLFQsynX8onGwDU2N
Vu7d0eWTLCIn/h/4NfnW0qSLTxoIAHFKcllfRxBTzAJknWDZwKZgR6uAQ1/bc+jo
xmuJ4eeropB41TS1bjTn9s0T8AVjD5hFSHtPgT8iAJJX9OPENTeNiB1TdmimyO03
BmbAU3ANjtqdM+GSrHCODp+zCGXtChbuuaCkkBWaTNAnF+Ao8RVVVWyojDdnjO0J
Nr1VzJwwG3KO02KgZ/j1J/f0pLm0gR3jl2g4bNnm7pjutI97Lh5yuVNjVHZX7jEr
VIcxVYe/fLloNmmuPsyNXmIHmmQ3TOovsFStTklIPA4qy6E7oSJwszkAPRPn0LaN
O9HpTvlOCrDGYqknlR1TWxxTdEYOqZ1GRPjeXEvbthbupASj6HjelgX7RkAoT938
ed9LzAiUtTb1C8WE1uKUMRmM7RBKT8yOYONzuF4ufN6E17AHagm8V7RsaaVhtYv1
vddw6Vt1qmYS1vylszj4amuoDOk3r4GpTUvn/90cGALMbtL2eRmkkIVgfLDj+2zx
HpFvi9gLzZ+adzTcfNjUQ7ffiJvSX0rE0ma7Jf5FUXR18FgPQ3E/o6k1k7Px/wi7
pWt2fW+c2AHjDoz8MNTil0aD4SH68ClOnuS3wZUbclftjX6BfIJbi617buX0hRu6
Kh/N4gH95jsb29EfazDU+jZprCEWV+mqRy+YSRALfuLmeXUMywvnRrkNITbyCY6k
v2Dj3qscSU3exmlL+eIwy0tSoUhYHJaZBElUs+a5f35QMto8Q05Kh7MRh6pgXBld
JV2bhitJKX44bbbIyP5nUSRbkLNNnwnb070C3Ewe+lb376Qi14CfxnphiIJXL+dw
H4QRJpO4f0sBZurhV6L8CLIooedIHdeiUZWXHI32vNMH6yHRkfl7ws9ihGb70qeT
gedHfRFg9K8YvS4Dd+nhWYn1dQ3O2pM0tt0r4HCFIJJxgkkc6hOuclReI2hl1/57
wqDZUxuoIrNLY3fldaJxvo0rSW29HRToTlIexe1gfiDot0wpGQ94uU/6r/O0CKtS
28fwc3E+MFfs3+Vjno3hXDL0o64frCymdxCgi5ElX2shRk/w+Ksngc9rFC/YVkL+
veuCQmMPCDgV3L5oGYGjVfJerpzL7+WysU/0hrECuF1tO+Li0Sx0ij011YGAO5eN
KOkzjGnSc9pUWJwO3lEVO/e8wtWNQIFU/FHBfMy0AmYXeIsCIs91CMRYN/KPkbX8
dV8WrOlDEWZsV6KfRbbgooCLV4MOxKv0H25xDlS2DnEWIw43KzIwebTfciFIaAzj
ZvgfgaCPu+fOtArZ9HfPD69ViqQXWd24ypdky1eEUlKAnWlwSUVAwwgiZj1rrqIn
4e46Q3l9OQUo3qMHDcwFQRw4YTdg++I5XbA5ywJezutaTwD+ynM/q+geP7blXXw7
UFkI2RGkgEMXxfDltGDH5gF3Rckzpx1dUHARP4A/a8G9GmZwU+vphe56l14gkZ+r
XQXLqyO/c8ih9XIBtBgW1uNqA8OYnlMRcZALuQl2kDS+Bj+zpuyTnqPMipyhtiSQ
NHV/yqmNaJkfH3Ae17l6LsjKZVZOTu0l2dWgbOOIJeAqqIuQTNGtdb2hWvL3luML
u+0EGVZrmacw66OiKGRJa7DmhAqNx9w/5CexfUvZMDK3FuJlY9bTgOmgL0BaOy+f
hqFtHFitptw8emCJgynBtfyOFVQ5MB03xzVgEixM32i/4x1Dbbnyi+rn/eu8UlC/
gLOk4V4h86bnn+St2cxYGcxP88Blytm12ZndwdzNMYABOTJMGwuMhH7BHHy0F6SR
EqMJoWvAbZysoXOEntLa61CbHpS5qgz6yTPrBhr7jgnC11OrWPlNF7WRw2zLkWcw
jerOnNMFNAb1+oY28hUR+I/p/5Csz93CEmJich2XZJUZRTiClfol2eBQpiwxJq2K
EIxTzjA/bn6VqisTfgY6SuM80Xg+GwRpQV6NagMM/lrOfkdR+K/vF0jJSDbv4JZj
CW85PPWbzRfyut4vC8cFz+HKCbPqTYmMRyOdw1UBfr2W2mmQiE9kaadfzF3MAJuw
75kg2mOCsbCyZJSVaoc3QjQIh0Yj7vvgGXHPuLaIwZ2POVnzWp6fhsq499yBIHGi
akBzc6aejc+TwnT0nnCPJFTVhchG1jxUuLnEY3isHCFlM9FSpzFr84JntIUXSLL4
z9KfcpIP1juOwoiDQ1WY+9wUeKGtQP6yUiUOLeVmMJfEZn/yDiSYWOxVo4aCIfFM
IFvofy14LkVboptgBDONdxb8vCANOBGLYRv+2bzImag5fjM+50WyxD6WCNKH5xTN
nE4Z3DXEbnjuVLn0KtdliHpJQVc6RloqF9a1wl0rpokzmfJ3LrM3mj4/iyBB55Zy
PP5ymJj5GUbVMLFTA/PVKxVJIWBGXR8w0fMLQ9NUmVKA5i1oT7dwdvB2ca5XL2bO
OXjzqDX2owBkwzTATIEO4sAPaVpyCZLzirH+WTUiVNl61QUo/MDvVLXgdpjc65Qt
vMEw4vGlDtYbpDeobtS7mwB/aCvJY5FT5bq436pF1xTCA0ZuBI/RdwmDPdONOoYP
pqAhcR/+SU2Vro1WXU3Bsm5Dv5VOTLhKmrusQjw4pef3Ep/zK3GU4aLS7rn9zHg9
+DPKFbOVJxQNjdLR2NF2qUg4CyWoT2uyP9INRHjGhivGQmk+EQOyqOgQAQxK1j8l
WAaIG0llYrkB4bDBx35Y8YcYsZpSlPhnHj1aRcSOfR52RzVvvuP9JizI7zVtSutW
HSjVRK6okhBDBQ0IrJcdgAhSC65gZhQqXfetpxqqtJ7enR9jdgXfU+xR9O2kv2KO
2chG9mbEecpSdE8EtsAg+fnRiWCKZsiMxQW72z3quk2cx2MzRsbMZFfP5yxpV8gC
qzVgasvzj1wJALBZAtuGmNqzN4MRoO5p2gErs3YVmPie3NUjI6G9dQ1T4yJ8qsos
h46UHqRys7LOJbb1SgKBjz3VG97TmJ0K341IIVa9S/4312ORRNy6Mx0eFsMAG4X5
5VSLIA/k9L5C0euktAstLelhgMToIK/LV5stROnL4V6Y5FwKulq28IHsY3F82dsx
53YhF0CJHCUcXxnPLesP6q5BfcvIpd5wRpZ8uuJFBiiaz/AUpjNyNvhLINbcXrW0
B4Gb00UUe+pv69waw71mj6GmgoOPDpfnI1jWX1PmFmGgJ7jZX0BqDePiCxCIuWyj
lJG4kzErXEX7Q5pWCZWoFZEmxSBLQo0yjLsNB5YZrWXLkleWSXXgbzljtKmusHSP
bV/bnLSLrv19eeuolS0bmiOTSwKb9LjdJ+5r9+3LMsrj1DRbakFRlLxjsAHijIFK
Vh2aWD4ddCRbSMMknZGz2yJjj9PwGzUI/sshgzPdUmLS1as69kT8eS3GVVijpu3r
NdUa8B37miduNsTPAxoNEYs81yhLracXKfc1FNrG3pGBH0yE7/YaB4/vwOEH00DV
dmEV3d6tkt2Gqx89J52FHPoEsbQ3dIBp0WOv5BY89pu1kLch5dcQUsW5rQ60Pu3N
QNHV9evELDK8/NnedJ3oMlr0dHrdBMut2D2FSsYSJRbtyr8KRomU5Jl8NTVgTyO+
jBdEKE4r4nIDkFb0STTlAKuIPeX1YQ7u+VBHVrc6i82GcNqo+Mrku++mb4QR9W0C
O39v2tG3B9RvaCiWHFSwDLaaXH2dxKH6VKkQGfZ2OukrYmnFIuQr+OHeR4u6LGpi
WGtKRsYHmxJZ1ANfW+bVstv0RSJ1s4GVWosdQ096wyQ69Y73kRUikbzg537L8MVX
HyMD8PqpSR54NX6n7QxBf1Yd8HC03hH+FK2SBN4nbNDh3611aaoRwYSwB85RqJvc
31Xe10uPOYCqF/sbTGKPTqsJujt0nS3b6/6IJIOUMIjNZtGRw3d6XAKhwRjuYVwu
03NzvCaI7CNwFAOd3s6Q2uhXfEbJLqumsY8tEGTUUiBtDMxmvHC/DcE3NLW6UiLg
78aV2eJNTNICoP82S1qE2jxtByRsK54LkB80478vLoCE+wbh4D0qaBsdE/dKvzS0
yxdxDlobeGN9AZ2b4c+HZJW+H8j/+g0K3IPeOBj4lbcmZrhqkTFsypRymgVxveiT
Xg25nc5hEpCkj26csyZuEIJHtXLKKf6ZkxX0NPlpHdpN9HEn7CmGcBF/Pd0k/Zuw
Hi9wtTa/+YG+NoTrG8oYTh6ASh3KV9jDh9bexHpU15nfDReakAxPedWnfCAXEzXd
0+nkvYrpxRM+sSNWoLPdCaRiHW7jj1GVZ0crAXGYqa1CTgGNhTKYlz/cc/s8Rtif
FOPuVIM/PHN85qvJPERiRyiaQbWvOPdct2UAlbIGc4nAnJA9Y6Xx3cEDSM7yCHr9
MGIEGGxn9dke3tmmEAz5mizcP0Mj/O+KWZZVcEFA0bFjKEuIzhPj1A+yN+AYfoHG
w2ytFmXhA2SeVIVItg7rE6SygkHHeKgkK9x3u1XzWlzxcu6pcAdxGbMJ+YasNcvr
1+LUiZm0cMPuHCJdEIP/h1sYsmv62f2K8fpxnlbKEwuF0+YRvYxZ2/j4KY5jRFJB
HXKArZZw4i99Fn7lzxMcOweiPk8Qgo1ePi0/ugi8w2h7DcFfnDV4jyByaQWIiDZp
Rm7ASi8XbtPjrwp3ReqZ7mZuQuwKR5uZbd1gi53Z/QUcbUmqMj+sugWJq1EDAB0h
BZB6KzZKPGrjSDZjudw7tSIeNu8/V0BDdIqDXmYGt8G6GYGXACkQz5noLJttgmbC
0NJrx0K2v1JSxvqq9aZQTf7wKYXSNNUCDFJTnt9U5nrlC2HPc2ZbZtTjB4bdajju
IJkGF01ba/nHw4HHUTEn4NP9yAQaU/av5NImamacSBHfFe1QEHPcq6UvGtU8Ugfn
G7FiuSjtLow1tutQXmnQRdZYPuznUqy0JD8QztCaPJz/UbIc2CbY58YTBwpHawTz
m/6dcL1ZoPKcpqB0dnWGwtzYTq+o1x8xYrhdRhGQsj8yMdWcYzsw2XzHkfNclMmC
3zkk72qp1rEKm56JccK22XROBZ5yNpoO/692CT2ox2PgZ2ItENbecKfQV1sBy1PN
Tc73AcDNBQd14JBmNZIqAhPbZ9UetghCQw2CTVsczAuXsjER9Y8zrKZcLP3hFJen
jdPNX6VokPHQn7wg1gDLO1TsXSRQ79Vw5/Pkz79jG7MbV8dB8DihUZW2qDEgQpuP
kCk4CAXkbJnud1elklq7HfvW6UwSGbEA/5DXqjOeM167PtaQzXHPqtP4lKGy/wvA
UrlBuLE/vuz+5CoopCUlcHtPXowMWHwqjLbZrS+TTn0EHOb7ZQL7MaLrSEFdaxjR
wChaS7YHiH62vKTm9Fz8cRItEZz3B+Wn6F62VNrgbuerZlZKiD75lcUCtnybDwhq
60hSElEGnYFfHSrQwALHIryJCFbCEFUEqCOyRUkEcufLAHTZIpABzT/K4/iq60W0
a5VAN94Thtn7JDXM478T9v6mQixANz3jYwOii5dESWfhcp/DvDXsztU1ezn6othU
WpE+rTe1Nw/+d8MatXH1htyZHWVSeDJX/pTSkmAl2XCGM0MygGbWa8RNpbssIO6u
aSgSC5jNojFNb1qwP30ZuD7B3qxTq8fCeQap9IddmthmF5QszeAQWj/e9EHcdgAQ
ptE/wyzbWb/OPRuBtWTDfKW2uXIr0gaWWDUDJXIuSYSD6JucI66Ndzqn5e4G6HZO
eYthuVoWhlylxriz/PS66fB5DxkmG/ujQcxLKxy/EKt00l+jsptD6mg2puOZloDT
p/Re/A4E+gwbTihlOLkpnzbcoAIkRLqeEruo51/BOSzh25nNnnT97M74/oxYPw51
IVNJJKLwomkxQTgG1ARrOY5jnQw9ZOGX65+77JxigMKUepSQzAGp0Lt6gSXYMBBG
jXxwVjcWWlqzO4iOpY1ZOoURQHyHxcktcGyr9mhlia61yulro/zkyNmyF/kwBm/9
1R4N+6kbM0J43cnfVZqoJxxMB/mZ4+cDo3hyOMsLFOdLxTBvibwMv7b7pTU81w/J
d5chzjpIjyADRo5X/tjlv/wFxJK99l1ZCu+++Mu5ShKjujVRuCRbyALal6THLwPL
nGHF8jy9K/2vtWVyN4UWRsuz2m1DCrh4upWN3PF3trA+DU9pQgxAocejXgm4JkHB
rMwU9zAygOJviVxxBQ83kCejXfvBLQS92AapeuPXE1cpWl7fiqHexmVvAHZN0gmc
yUUsBo+F79wc6lBooNdxXT2AiwAHy6NBpPVU80UnPUvSc34RMvOczL+2Ex2Khf44
snc7A8TTsOCMu6MPvQvsyyXSIgmo2sarBde0hawqgyBa2QE8ffBJj+zUYgtJ7dpE
Ud8FYAshvRfKxNAF6i4rs8tqibjo1nLnQvD/l3MLDztXh/ToUnyw+CK/yajw+GXi
TlF3c4QUPsdT0NCBoS4oo+akKH5ZX6+qiq+4u3iqHCpCGne6SW1wWGIvJAa3Mg0n
GdUbE+ytMYm/O6eRnenEYxLT+masYtEVrCL3xrEImOlu7YZrjUJdKYZ5hsmXf6SU
/j8hSBHQ40NMyxFLm8H5Us/sMER8hyFYU6owjZi5GFdTWd+RPigu3BBeI3YeaBqn
CZWwdYYfS3npZa/WdIyang1UA1XCiIjblDv+4mmA5FG4PxQjZED2R32CecfrBzdI
h3B0H5guJ0wVqIyzhm7X+lAKnQoI2BfFzhxIFdZkkG1afCp2Ov+J6i30l765DD74
2I5bDMMFpcFOROvJEp325AHySr3En18xoegIpqi3AH0kzMrNu46gxFPqkGcyS36V
7Iu40itjTRMHEqZ2Nb0YLHZ5e2N2kv1i1ynWVQUtP3nNVGhLCooLt4PAYwn2Jiwk
QLAcpnMztp4zhEyu7wJDc+/CP2TvJKxFxeAW7rbSuWVUevIf/awVLEKTrXmiFh7R
8H96ByJzFmWy3Cy4rPjdm7qPwQ8j+KHnJyZZqdoV2ZobHCnCKbOOYkRjzbAxxZj/
PWTQPdS3TqiO2arZ+34p3R0GSlEr50ky3b/S3+MhKjJUDzJVbqgi9mdEbBKNXedj
vyZEtOSOenTqk7aoyuzgfq1K0Dmt8E6T6WYUTxHFAMK8wP/A+26sOTSUn2j+gUDq
h7WTUw/ep43RxrHiuSCQihfVL1qCgEtZjfJH24Pc4JNwTSHHeYnSh6Raxdda2nVb
rCfUkaU0hv32tYSALu9SXRopx7s2x3X1012SPRx/SlVWBbFtj9X27y27g7r8F3eP
LRx3efhcBUG8XdYsDLvLfbHE7E1uZDoXf/VIhB4Wozpv5FyA2eJVHEL0CK47YIk4
GiwyKf9aqZLALVwqIdCHeLrs7mFoF3mnSwmtqFtzVzBZG/gBPnNbx194Pr/7Q/Uo
4ASo865gYAzeFiH5G3zja0QmNMuUSDktuR+TdiF0yoI7tqf90JX0wPwWnEZxnuOP
oV+vKGsNAfKU2Ew7J1E1jBB4ZlCifcZPq27p6vrglDlWnhrBCV61Qrcw4nmn8+sL
7I2pPaw3HU/qzoNXU8iPtq+fl6OCtjYxA/t/kkzp4Inf6771E4PbSX1vhofdw/DD
WmMtC0w60PooUFEkhjw5M9DjQ/BD/Uszvwl3kJLjjb96TRazpzNG7SgxGVqsJ/AH
bPjSBVnTk6/c49aVEbZEl207RceUVJ5mG0eUMs6QOjZq3SIi33DcuRpHwwB6IrJW
HV7dkemCB+Xyg8HDtB5h7ZS86kbzrLcKSuUdoCpgp5mRZGHf5qkIZKwZu1PZKk5Z
mp3z4X+/iq79mF6SDaayxP5Asdqa9xcD6232rUycrxJ5N6J4U4m9tTsUoeInFDsB
C69DRh3+2KxabjNsCP6vcX0RzFBAjkZfCLpZAxOA3ikw1HOOVQ8iVaCDHwp3+ot2
bhNPSP3KIf/MyA9X435MTLddMmFWita9B127NPtINOd6vYF0Q7clesgkX5ZRC58Z
dYivjCzmcM1RG1pw9BDeTnFuw7TLrFncEupIPLJqRahO7ZbmkP7BEir356a3fzzn
5Et50gw2jwhlstBeCrkT4H6juMLNMO0SPg2NYjtYeSzqBozfN2FHVTHLXx+Ml5Lp
UBNSrUlf4lvNkm1O5L1zjN0VKRzWgfJC0127kbhfoK8FVuZuevqBEKBiz53+1fWP
EuyoLmAv4cQY7S+bIQgIpRB5ruK4Lszcwul27URulCIam7i8OMUfkIIMoIiuNIhr
fA+PKjd97FbQTT+2TJIlyBPuR5sp1S0kCtxU1Xp5dTTO6/MJ3pTfGp+7WgVD+hYm
8Nkp0cvZcRQaDBDGxWO/J4qQnzvKqyBZObHIrPhQLOZKnHJMSOR8hKq4eD9ZJL/T
Weo2f09bWu7CeJrecAzdFse5pX3xcB9nIOEjESt1PWfiInV+6UHOEr/Jc/QAcfJv
B041ppz0SuBEasOF74xzuis+Qjzx+sLQB3uZa7GV1prhVjTEZ20grbRNci+J0mX2
BRS86AcSJdsDaANHuBK0YhPeDTgeyEIgJGlIEE0TzBeFfjQ+xRE7+X3jahHMEzP2
gY5WV9qvtINee2E1ql+VhUwpbYjqBOlECG8tGMXJ5rCtZ05+w0LpwKWPJ333x/OZ
Gj2I5gdH6aGkWBhvecW2irMvKlppq/mgAOvUuCwsGzeAwlkL6UDk/E1iLJRiQuzG
/vkq7lBdklD6mus9IS1BZ1GKefCLSilMqcoHdd1dzitfhy1tChLbh3jl3/dk7Fez
r7s4b3GhfLGGv3rpqyVAxiNXAvItIyUZDTdaXBO7guTepHh9tCdEHBJ4LtgZx13j
HK/O4Q+drKE2D+tA916t/wIqYb3gbl0cE5BiLiy36WwJ8bFwTKUsNIRWYnCwu5LA
3m0N8uYIIfdMHVxhBH1ticRqwBP2J4GQblQzlkJ0K0gcw/XV1M2XuCH0nvMuoE7/
abuMXXSxP3MgUUvmcYqSP+5+by0VSz6m/cWI4R71tXu4Pa7KEkbpzwcs/BdrOeZh
v6n1MrKcPEVemQ5HoTeHwjNUDIWUxChe+F6DJxRQE4Ow5RLNBTOG7zrU//ZNSqiV
mL/R2Tzn/SPOwygDlPXfQB6Cv+rYBjxsBkmhe1T8jDdpSpzjkcg9ykMEQW+kSiqs
VK6Mhtf+4lbz7dRr1XPeheEST9CwycPnkk0fY8LfV/9Fwq9gI6a2PdFAIodaM+tm
cE7jmKXstjaR/Y7w5qlO4J49oISDWelDauUEhnRoc2gkaj6U2QnL9DC00+vf9hbW
9Ybnrgru40lFXYrGPWOJf7c810HtN5mdIYeIdf03rLcx3f4CeEfKlpSILLWPwt/P
mD/m4jIBfcO/q94QzEv0puEfDcJagxpRxNyQRJiphY6GPRLLceIMOKUHLVC9imwB
k2iL/OenvGCH1IOwLhkamWaOSv0ysSi9FiF3cqopehdx2vwR9KU7LDRFHupw6x60
xHYuVTTSQlG54thBDHubNPFk99Glbw4AfisFs3eLjju/PV3MtBjEYQMh0TzCIBWc
yNY4FtsMN0OcsWC1R46XJz1QEtqgGnrJR54y3TfeMFbKtfdbjLbk7E+5lzgh6F07
5EpEa36zVp0entWrwBtXfe8p4EZhTkG4tb93iaUWpEz42zeMcS5gNN5dU/w0u86f
zJgSiyTY3APu2Xu9LhAWdAWZXt2dRF1M/q4XqIwwYNjfcszEnhN3VvSAS+r5yJWy
fTnkriWquqG60pis3UxP3WnvmxhxXBPXDrdCoubmbf9qxbeGXd8m8tR92Rf5gAHZ
+8dLYtiU3enuJ9WYrvwyUbzPa7IrpUbwGEylKDbBNXETZD7MeYTEbza1v6PHimla
kKsw9dI7RkyKtXevLQTC8BdE/NDTo02sHB5I9dRUOJ8tDh7cwmgSJQ/T5fw1nsdv
WTnrgN6RrenuwVetMiGuZuyVkQkzNuYNUYw7OunLT7kkm6p0c3Rj0HNdkb2o4Vt5
JtBCqlCBHEMOpyQDHXGfRjx2N/lQNCnbJsuFk6U56dMaXCPFxxYODwCFhFvdGnBO
AtaLP3nZgknFKsXMR0bWYYH+k9cVmgX+J4FrYTyyLrkhHQrHRCW/BkuhMGv3x27M
eC1NaZSWYrmJ2eZHEANc+LOSgeSmtd10Qts3H1McjIqYiZljBLPZlsp7GXnBs+GF
mkOkehE914f4ZsLWIjU66p3gY84sPjqqbBgj7ypVqSj+Id2cwVafY5CaHidV1iem
sPX3WJHPnuj16w57Tu+pUIeePtsG3NgoQRC/PV3QqfXV4b2R3nTehBMFe9vyusio
+NDbv79xuTqwG1NT8fiPhAAstp1jxFX22Ah6p2FtU5EwErr4gcfRzg8++G32bUl/
qOEnPlL7D0WmN321Q26lp5taFgnhhJzdlVMZewrwftmBwu2nH6suFiWn7H/vlTz1
LkSFZbM7k1ID7iKM8Vg7fc044u6ik4cOmZrupmm8QUCkrTSuhKQIrva1Udkl5DBz
0Up1P+2wITIMW+mOsPzFVo9AIoofPXUfm9qgWAJXX/W2egkRdZ9MfHaeo5jI1uNl
dQdfuL1fP/LIsvW8yBdYg1Q6RyJibQF7yp4n0QgwuOfDIfExeh8dhG2i7cDWTvAw
nihY6DER/TegGpC1cS+vdWDPbO66z7Ng8CZJzt0F+gnIQeD5Xa+NHw4eM864VzPc
PZGbxQvKcxR7F7mpQ3tFgM/WY1Nx2LTEbn1HbsErKWo8dLYD/GpAgDN8PLidlvFs
NDumjIhMoMPnYdkvLkGrqFYZVQwph9puGC3P8Z/HF2j9HpCc7QeOzajzZn+QD3rJ
tLRcjqBUSk/HHsmfWR36OBOVvSun9D7jTpoWDum+qZf0CJb0KVBQVVXoteti6R2X
1AcMNCOaSMikpSeuwPFkrXvTYTU39cNJQBhOhOsXWrVp2+4Rl+Rb4Cfj6sB08ulh
vVD0JIUdu0MjfWUxJYgmVaIXxKOUA1BPjMbDxBT222Po0nQhVB7cdNAp9EdUUI9c
JeDihQX9uNUXtP/1TAMpszcpQA06FDKpeo8OqdmMvijQGWYDxP+/BNHKuDf3Ky/P
ED3OTp7kExsnLHvCzU3+J4OzersOTAhE46c30ZW43TCyx1bhFZyCwbYbLmx5gwCI
2YNmJxJ1lxjcHpD5DO4219SV/NdJEF8WRJChcaRrOdtwfShFVGuXgzfJkjOq6N3d
tR1IiT2EHRsbdkf7QapwuHssg/xlmEqjScYWl/0uATqgn0MEhlqXiOpKwvWotqpq
EMlLmY4ELJPXL1PAGABML2MDjf4OIbwyvEfT3lRnwyNM3irLBDczcTAYxPjw8emB
fNY2z25FK3h2QeP/SDZZRSXE7IqRPkwuF+ARLDPipFhajMDxn1GZuUhqT2vYzBw7
Gj7y3Vr4su3vCtV6NgDnEtVGwgdmEXKoN8fQfsV49kiVpACPr3T0S29r2jEY9WN5
lJDJwia4K6dQ97ieCPmwWwrFyQR07tJxUQIY4lSVeM4urAU5v80o9YYKQVMJYzKp
fPp+muw9tBTI7RUZiz3RcD0xDo1sXqF6i2/4UzqSXRPP3PY/ZoOdT+PL9fouK6BH
1FiLwlfS4r296tl+ZeRwsqWDXt2cQm424uyf+YNrRbHGEz85qHtLb9nyaijfxa00
dfGdgbHayx6JkzOyQi/TzyaaU7ePr7EcCIXIQoqUH9eh2jdNEVZdteeFrQ4MNI83
r7zeQqsw6XuCOOWbHXthpGmFabyFWkxQpvwNpDxe8HoHz6S3bdVYhZiTh8aW2Duc
JxT8VQSXRnB9wH/pWB65WB7bLYiwT1q0z8gextIChDNJ6PiVXG5ba9CxtVSmKnjk
IHgiQDKG1UwHhQ3Aem43qk/MjJCIa2jjdh/HwV+0FuSBR80JZFPgfa7sK1fAljcD
OHCyIAoaEoVduZqMdcKBAs3XGIRyD1jLmMCha8Iw2KlMo2VL7wJqRFYGH4+wfpeb
JGtPO2wRny5sMtHNqKOU1ls46xngZvKhoM08CHKgAnMkeGFMnq7vLu8sAg6sAsm9
/e65JiJUdvKvtlHxwU4/n5a+4o5+1F/8/G2XCWWUMRktVlGHLvbgeFigET8Fo4WY
20SetGWa5n/0sWXzXXgNe3W12oMpeFf7nbdhSVTVel/d1yHv2EWt9PLIWHlksLht
5aG2/WnrQ8AbA4biSfIv4i4dE7P1Gud28VQ/JRez2pn/1oJHBJ+qMd2WWgh6KjaM
8LS43M0nTuXPTRthBcumuAIPeMKHYK5fTo4pKX5Dsc08EpZSw3XApoJRBneafxo3
ytcCV3RXVPH3rLiZCcsqepiwWEg4T0wB09Lq+lBnORPSTl6ieIEg6cg/iMfUxb0g
Eivecd5fH8nvz/4Dm5rCMeMAfOS+8PbugP3BSCBdKZi11uAN13UO3PQc3IgprIkH
kqhIxyJvsiHmssxQGDjZOaPYbR3w7qUqG0Rv7XDIsghkZqEPe8QDMTm/Yd8KeRRX
a+Pb0alb1uDhscISMtNWCSJrv951hllvC3v5+ey8s7vQuxOL8ZzLa2+kNUofe/CO
GFyZmGmqmuN8SmNx94jLsrwOQksBALkj9ij7SPfi9loB2d44bWKBk1QBUF0qUUJP
UrZg8PY4sBErG79xnCv1B+xTO6wI8NvlRRFk4yurfHnPaC6FNTXZ7nVDNRTqJrRS
n/AJQOuwOIl5cMe+ttap7cfskCCbeOqx5loBFSzeqJy5Drt+m/V/paAyRAv32AAB
jXUWOZOxD39QA+BPOLHrOozb0ol/hD1EYR+U14YD2DsHGOeEU/zyNQ8PM6QOJoe/
QG9X0jwWAwms/boKNLEml/jBkusVKyqh0bqxFYj0xRakMR55M7Kwllkjg1qFx6Mh
eScUk5lDwfcyRyrzN0ykoYujPRC+t9UDGQmxquX2LN5oOx7C0PTOlUdVrhR6FZ8e
kff8DKSiy4x8fiJ/kr5UxCnCOTwGqesdZn3jETMK8SdhvFeF7onkXJeucDkBGTfr
VF8ITzcaUapTpDY4P1IuNZ64VpPMGkWzh89TX+7jqGd44reCZqMvUu7vS4Qhsy8b
yIBlLYzgvDt5fl5DBqeEUaaP1YWtEekHxYAUX6Ri9CjBH3xMKLfivIhcywI0AChL
YWItblPnJ8fAbJ0OjqRgmA9HHmBcATYSLU6OwKadHfa5uB2KXqG64FISdaPdGSmt
UFfhS/sdRibEm0owrbNmSqYnid4w3sRFFq39J9iKAkJ0CcwwjD1ba0qxP9CCNrIP
Cq0yr3Ls2mGEhmjs+kBvDV2aIe9aifDaX7uz4NDRT8fQB2TrzYnmrAck63r6+56m
BWqilmb0APheAIlNIDPZ7bfjNEo0xMyMDTpgGTN8mzeIc0AKyZNTOkczzBlM+qgB
y25y7B4UPEHHCjdfsHWEhX3sDp+6vSowNIO+RAgVfoh2bwGO5QHrlrBCCq8SmnYm
hl4XuFnl06majOmI/sl4pLhNhoLjrkhrk11pjNz1EjhMWFu+OcRanUhko5S4Gheb
SNKSaCJZ+lr1sU7Sa2tzUmNtdJdiIsv/dVTNaNn7Oe2XfRELXofu5m7qdWR2rDiS
PST7YqaVUCChzlXR3fx2R3iT1LKifPh6oGbY9WqIYZvQ1tuDUCKaXxzds7fg4g9Z
/cahIJ7WMs0yeWBxiZ2G4RZuPc2i89vwGYrFlBIB8Dih9SqY2unDYHEhCESzbFz3
oDI5M/nGYEFWGpdAo2/3aH7Knu36VmCGshPy4AC8jt2OBItLlxZHBR07DXp8aLBl
NmwM7wGsRMFaGQh2lqaI/t66Tuq838soLCjfiHFpAuXea0dmbMbR6a4lUblm130b
VPksWfzacVfXV8mhBPOYmQ8bTx540Q9HjbWdqeAxn4HZ1fifgZXrfUg13feDTVkp
SvReDmwdV0RY29IZ+wZeh7QVbSspfUT0yRp1GndPhTIaITsijsDtTLdsHY4I7gIJ
N/mMhMEj3HMuKj+Z/DsdHe7PSlB45xi/hZosoKkZqdF1ND4VDoSPTFE9Whx7IHNF
4LOwDaehnh5Kgsryfx3eUOhXhJC4KmXff6ZugULGZBCBcGhpne9/GVHL11kPV0Ju
x+F/6Iep4PNfo/JFTkRZwNoWRvLV5Wc0rozvFeIQ9lDw2xulhZVhhaianLxgR+Q+
QrCNrySaGcthS/EqsaYqTC+rdq9Xm6utRBZPVsAY24LcD3Luj7WbffXD7Yd3JKcU
LxV5EUdG3yRqHfz5Fl7SPhOxRteB6OZkJta5nkMlliN2mF8Sv0xS3eVX3k5ZL33v
kUqAN6L2raj3f3x7zpKYxG2XohuZROlEddIy/ZEPOZD4LBI/as7lhE0v+v7ssCUP
zZFc8UW8FS39ZU9bCeXKWL2susZ3XcifEQgiWCc9SV1MGk/ImP9xQO81tNaZ4K7n
Rxal6Al0+eCBXMXMjTvq3WRB63vKavEf3QJnosdgB5q5WkSesRbqWNc+oCdL9Gen
krYq2LODFLlShvvMfuNdHMw9bq8yEVtgoPVVRdnc8oXBvMItTNWLWkPvCrD3xhZ6
s/O2EUk0vfkAjaDLMGc+PiP61ydab8Vo9vRr4EPa36ARwBFUgaYvBA6BUtNO/m3v
JIDXWv2H3lA4q10tC3Qki1S/wMA9n4SKsn1YRaDE5ihw3G8/7soCqHLsX45dQjx8
jBO3RIpl6qVpY7xlU+eS1XqNy+FlgZooTpumnlRTHhzX8Hc6W2me0gzmXu1l4XRv
/RHFwvHqMB9l1F1iAx4rOMzpGWIEUfdD337vOJRNjFgBhCP14H7yfJbPZwb2GvzG
HTQTZI1v3Se0a1i9iDa8l4sjQM9CwnJWVI9Ql+frUBkjVrfpFDtgsjmZ7YzEo9Cv
Kdaq0E2y3WXhH/GnorDzvczRgrWpAks6cBDC4wkKzL2HbUOpJMqzC8iQThPK5QNU
8KSx7XhLHIJEFmO88aDsFbZAHJGUcDHt645tjau2pjy6hXaVPJQyxn7dwXu0ZD3j
6jl5DC/tSVuEaNriTR6J5tTbtANsyaVE/+x2wctouUNtrJImu32xJmcHFN72MfFQ
wsrg59WQDUdMRqgJcUbvT5BP2Nm5NL6U2Wz1JxpGa7VC4d7RzbUUOU6F8i1fzfBH
r3Jrl9195yPitkX38CmShgsLN7wpXwBSYRWKcJf8G4zrPiD3BMOLobvKpyhFX/tS
8mIdTQMdLbGLrrxSJuczbF8swH/lYOkiwF1v8UbmYlNpeK/EqlQO1cypbFbUOGBm
bIWMeASRjHfPaVvHbQvxb1dIevYJFsfunR6eEI4YzeRIwbX/AvYbNyabTERKeuMQ
Ic2mnRBTAohTavQEXBZ/CPoGQouEfxkvSGaNcTXSzkGv4obRKOKVlrHzWctZJbsa
RSDWKZQkd+iuwgUQRhF6Rb9z1ykEa7edbaONDFVqZgHQqrqZ1Rxon3kHS+p8+Mc1
amxxlKRgIqnHcQ4kYYhPXEveL8aaQsSyYIwBGbWNQ7WyYI1ND2cO+lxgfkQxHhZ1
9m0/KV9zvUCcxpMtEJWlktXD/w1C/frvJaWWpE/Mme+bFnPnz52cVRyHOskg8H3X
iO9aeQ6BMUsPzGTUUGshYPM9GZGcLQKrsRSht9wphabN0bF7e8yyOktEnsGXUkRa
JqxR7ir+Gi4HLGzeAZW+xdTK8tUEJ95blr3DEyk76BDdl1sy03zUn7XQUXzSSm13
7LbqPN/8/Nou25Dcq4D1m6YiTR7a5mqj0VrswwRiniOvdG5byPdEdghljo1TBBzP
en/c4s0hvC/NVc0uqKDUSMfKy5WcD8gLaP4mWFw4LrDY+JAOTmDc3p8dM8Sb9WcA
8sgmYrfnAnffJUVXixz5fMl6rjIrHpdGrHth0vPxibA/ODcR9ZWX5QZos4Zf9jAa
Iaa8+xhwK3a7VdQpEyZozKgu83oYaG2xTXiuOoAi5Xtv97xgtqaC30H4y2UgTUay
0LkigJLdg/NcvP4CEuINUHKrej9XMBrF0DtzR+MsRd9lj9ZQ6gtf29cf2BZrOknN
jYy4ihUpjsuHDD0zJVZIM+9aEZ3LVbbt5VqvBCDAl6lGgbFSDsUmGyNiLRKMDwW3
qp9y8SflfzuU9cxqXdttBMtob//CUWNARssi2d9UgWkfBFbdpfzaOYrz9YS3Qt+7
KYNVyRYRKAvIsgwdOS6WhLNqyKhfs4NZwXhT6QvkZlhj+tJ7WIXqkMVaA9O+ZNti
wonW89ZKxg6irW0c9zC78b/6WZXaTYobgf/JfS5ll7IJ23rIlXy4OUryyDNFSy3D
LOIPuW5X+Dc38kkpuMgiQGJ4USd1UmHDqekKE2ee7UKgFSkx7Kchqy4WkC8S8e1T
Kd7h39/7+nypyFmMNcvN69QIEv1AvKLvoex5HSrXdQCynlxa/ZiTOj6rc6pJp8Y1
Uou9/HoZHTJDvQ4kuxr2nDNGIlb/AKmIH9EFSNqhrQ9hlt8610ZGNkiCl1yw8zQn
XyzVnq8GbiPsEQMfDnDkThrqdzlyw9Om2UUKLAUQ09+Ic8JKQtgg06l8T/Lyqi6r
mMasNHs5qH77JVLjoMTtcBsZal7JipQj4hDuW0iPgYz6n0apTc2IdRlCnO8dB+55
aa71SIlK4hWVG8FVkncz0Zg6FuUtPPYNyvqIJASfN8UsfhoVGWztDsd/vWClrOz2
HN6WMz8hwrB/IG1YP9ONCeUjHi9ylYvmHs5cCnI6FWozsO+jPC+AIj1R2SHC3jF8
+tq41Lbniag0JwYdF0SVCkLaAY6EWNb3XQ+CQlJ0/Wyf2vsk/qg5WBFZ0qNUdZJf
z5fS2ghxermXRvQ679pM3N/2bXQHFGWQm1vJAYH6hgDq2agVwTeZKtBWeefxGv4T
UdIPwvIDKYp9N527c3uzgcHY2ZfxsKozEBT46RdwONNm4monHRbAOaASKbNFAbBV
va82oEeJbC5+V6F9/J/BW7+sAVVvip78fJdUOdILvM1rBmy/39yj6y6Q6AweXqyd
9jS/LpuCPbyQKixBEzgy3Fav3+cy4DGIab+4KG8kiLzUPc2AXNUrdN4cW28TgjFR
08ZO1EIa322Yc3annuoSLb+VGjW1PmNQbfsBPvC39Js/Lmi13RwdPUb8Vq2Xe/2C
dJhZgaLG0BY+RDka6n4QLgFUnBM6VSuHWnh04xQ5r/doUy7umnYnVzanRm6BEn9O
A9qbIpWImS1N42Jrwd4TE7lr5noilIvBwUHFl2mYVrsBpZS89T66wJnziSb/HGsA
Byb5EDmsuG50S4MtYBaUBLXUywAPKCxN9Vp0b+4d+N0xB43VS7rxnwoy5BNSE/Z7
6uprplq1nm68zPJmJlW9b0tfH7UP1D+u0F2mD/WLvKPmzoJQUBBudrv4/ae5cwSK
xw8LWD+br4kw23FnSzRWNuyVaY4IwUf/xqayUhFs756s1BAwMf/KCujKzjFPyqbE
HXk4UyiG7V2q6b8p5TuR15J/beZQnOsWmmvvVh9DUcgKupwQ9sL59KlpLRSrU5vI
r6UXwBLgLUY4EDy+EErlti40F6IWCIJpNqpXKTsv5cyQycdXEcxYQzvsweEaebVb
Yupm/pkfzW/ks9XrS5ac3TdQJg5uomInMaVvN8hjhGnMogpm1AjyswsqblGRWgMo
EGcmfTh65vsDeQUjcQSujpY207Y/2ooltnq/vBf25mSswJHJ39Zi7pUpGZ3v7auI
DUjmQD3+cxEqGopbi+ILA3RiEIPGrfbyEBQKRPgp+2/adPWRw3THbrU0uXTXLaG8
wNQlLAMbgHApWs78j7Mq/V36DYpzkjmeasB9QsiY1nbKNPaIZSUDwMogEgZSswYz
IQ6ZhbiOo9pSjEan/qr/4P+mPu7ucD6MpdBHBSGTCvKw7usKOwyoGVQdqpAHapnQ
gW9l7MlCbjaVqjOPPREck1h5h2MugjRqq+jwVVchX26YRHGCunrnqV5GBqrfgVWm
MwuUqEDaXt1VuodJLHNo+so6TvwYP4I6zTAgzPMFoKqEptzaeaMSvQSHQljb8P6z
FecstPKM9pxtchignIiukg7sGmzufu36fKJhBlQdPm63NK+1r0VRGsfJGnR8dX+S
SqW0YeXjVoJiCyuYany/JJp9iCN2gZs+KWNA/mXFLqAJoYKFJ6ZvSCJP2sS/Y6/W
vyjDrna+nTTL5BW8rnpFU+VYBEFx50grFjhLQVAkkqNG+YfKwruZsZoVFxLKGEns
BQjUOgnmeZxJlCbNJE39KZLhC6w4uImwzznrpenaGvphFBKMeeu2pG2o0NrAud4j
Ke8shNMFwEZjUJD+GTdaOI1YW3R8YtFEyO1KLp+dJN2lWcXXxPTWP40SQpx2/4A/
v0xj3fV2vl2USPosCq2QCIdh43UGy3awegCX8w6z29L7xkrPVwHNrolCklJj5Ake
ArESH6XiZJeShNMfTCKjdtjT7qcQZZ0jDbmVUfYducgu3FA97QMUFBWQ1WT9d2yl
p6QhVuO5LFx7x7/FGrEBsL9ixGwV3NKO7jhEjCcTCQR8XLKYOS+m5NR+BjuU+JAH
Lm6rKE0bNwWU1QI/NZBPc0q373FHg/mG+Dd6JqyBVTWrRBn49CipypwBbsttR2We
45iR0A63awcffKrm1KMGNXES+ufChj+qr2CXFAUsvun1eFvEu6Xpfvi7GSOLpOBA
UzkMR86ceDpMRL4aRp3uyZNV9kko8KZGz9MbsOlDAlH/nxTFyZUvcPYQEKwbxwoq
cTv2juKdqUzF9FTWDIeVgM2M5Q9GefZYyITpWrc2gg1Ij1uDi2lQ/PtWBqmb3RmJ
H/BFQOd2hCsrcuCrAD0bxSpUAjEaSKXbUDKxfhcE3ob+wk27WeNIKN6ygrMoJXW9
SMF+ed97YVaQ+Ari90HpeJwuPt6DaomfO2H/LDiCzwl0clU/uAlmhM/0a0z5vc3Y
DKm0lv9LcurxV33y/v3k96kJMwKSngTgihxf+WR0x2b5uXLh1/7SsS7jtZgBFHh7
ECXQmNoz39TGK+ke8iwE3uNbQ69VrPMmj7pKXyZuvQ0pR/rVqbbg++V5ysTs6ya7
74/q8Erjkbj/ktPqppZxw2QZ7hdBPCbfDwBtQM/o8kJ+CzsOM1s44ZpQHXuN83tk
7HDQjhhwERDmK534q5JX3zhQAjekLqywrq0fEMU/x+3F8JtsRQ+FUlDCL6Et+n3t
wfanPGDVuB6HtvqGlPngXNFmFl9bjgITI7w59VtMCjpA62a77z51UOGiuLkN/Lag
xmkND0eE2ccBLaQJ7WPxEK8ODgk7P8RV9ubAkX8xClDAt8zcEwbDdpDso65cqjTM
FNvFx1mA/KCSqpOmg1AlT+6b9s9AGkeA63CWEviYBQP8ZzgLyAPzmRQXDnVbaVHC
LFUGdoz0G/x3ylw0eAGhX86kU50rX3xkM7Gtp1Vwc6DN86o7ZrLMqmSwZDp1RrRm
nCGmMxewJjn3O8SF2B3zKwg/svi6H4VaL7G/ItdYrcLaoLv4LOfozRMAMZ6QFYzV
ilRXYTiyl3S5MX6b8eOiYi6s9wU3rwwBzN4Zbmqy5phPXH6EpsgRrqTsAVON51FF
sOoflVEP3vW3SMHVcNmyUsfUV+6Pkj2oAPNGrXzHEGNVQabkqeCRxMICndtn1m6l
FbNngVEq/j2EMC8RCjUItinEnsoTONR57JJU01Ks4SHvB05Qx1yLnnoSYqRY6Q79
VN7+e/JyP+9AY6BkkbTzyG7D7MTLXoDFV5eR3TDq3/eU9Qvd/ivVAI+wbSlwRAAc
HqJzjuf726WgnCwTl+yK7uSsB2gn1yIed8+dJRNlat8iNNMPiVnIfaFCu7ObaeKq
ffrj3W11X6lX64jbCgoueOGbyD7rhQZ8YV+5aVlEROgrIkjtyLJGYCmXHnDLBbCb
PT2E421ICsPuc8Vo6eq1r4qMmjr3L0noWFCQh8emZYd+dGzKoxvBE/a9IOIbmm5J
/+WEHbVoecV7B7szrS/MlQEUhtLdzF3Ni7XrSDgteqnzEc3HACufhGVFNNf/1LSi
lNW+AOcpyHvFm0x51bDtwdw4n2dldn6uTYjbeAI0oTigvrgKzSzFocSZE6LGz7Wc
IDFMvfb+/TLUH9Zwe4EoGg6UF9vFdKglfBG74JpryVcj3HOqHWKewMN4vbaqScnU
owUzogl1oqJB/pkBEVTv+63KuwTzWqSI2lrVt5LQu94rxjiBYcY+yZHLvMtW/N35
nt9UYkWUYJ0Ufqss5yIvZyS2y++6bUP0mUNs9aGEbTJvsx7ksXTTtb65tP/EI4Mi
zO2K2yCc4mNlhKyxNaXKeCMjNp01jCSX3H1TaXvTNBx5KKo0HYqvUjVgqguQ8ato
vNDhT/RwF9RV68D+4778/eRausGoWxu+yWG/GZOg7l+9AZvSj1jt8aZm/q8ms5yE
VAc+UkPT3OqtYBtpygtcBRWXimzYh4XcnfVQB+Zj+mR7ITvXsDb+XezfCE+PYuVq
j8zTVSmSkXTTHVstRLnImSrtFc4PreRisEjndzhHpvwHGHD0wzO9XHu6+boCkepX
M74NUclipn6I8SC3yITMrgj6pfPxFKCov/WWQ2merw8etuKnU4C6YGDYZHZ3YDRm
yi885KoIJKVdBckxyucxWspNNmo7rg9hmEFT3Bfg8FHXBkZLGTBh5SByHnHD1VA0
6TYzm7/DuMU8bSgfHV5vy93K0HoRnmlYIKjlNZ2bbtuTHRdUNPgRapAWtVKR4MGa
hTHzjF+B+dBGkAoqaSpE2M3AVwrL+YKv0qrrJaLOnsm3TBA1LNhgqRPHxVWGV0rI
xAGHPtCHjl8XxGpRh6NVIrnYygvTcTlT+AEEC2sF1YdNBTj6Ef13mSLdMdTmr55l
3+uzrssOrLZlJ+Kms9I+CSMLYr4shbcbamEnUk9ZtZddg3XGprABYrR1OqcJMVin
rnK2Ms/7YOtLPk7gQxD7eof6P/fq9FlKPhWHRLKot5Pc4BzRQf6MAWmVUA3mqoyz
JBEsr72N7wsg9ciD0z6m0Y/4gXYyHvj33hkiA25Q8v/jNcwWl8aG3JF0chSfwYcf
e040AZ2MiDYcvPkw4KcuaIf0fB1Hm48wlpvrUMLJIbQPGBl2vYIG8p9vTLAcCskc
Zt66niK6NjeCh8nmX3B1tNI6mUSTEXeXKqJVCa42NCe2weC++XlR28X+pZi2CSip
7dz78pz7aN6ZtAwAMpp5o4SMwQrmm7zd76gEyrJJein5/e60OBwBi4MkBJy4OW01
A1PKy9CeEN+OBuwf359Y6FB2KzAaqYRyfRh2sdfkia2eL4MckK9kOi+pfq61HGBT
OZLCwvPbFA/uv2zWmP6TPKkdZ6VBdmmni9K+SayUfhaeen++7opEscSirQ9zCKZF
sC+hLzD8ne95wYW64mEyfejnEj4cIRZRvwRulc6v7+4a0FRKLYdQCNRC+eEgeQoE
8y3sK3EGEMy8YHR7x9xm4KubpNckiBBF2AB2QfB99yaYX2AHBDPgLgKeNmussiN8
3zXGifOMKMveU6FDC/eF2lHo5ynmotcmLezqHfVRg8cUfaVtjqdbWGAamZz6Xy1K
JEIzz0KZpiIClvT0O1iMZ4HpbTmzHDvph0nsJR685sr9sh5fw+uq2gW5XGZ+iWxA
zmc/0gPoZi3xxc15i1TAuJ24woQkIqzhXYwJc86NiNsAzOs8zZN79VyPNeKqo9jD
pLnVDr/WsnURjMJ+wAv+tkT9Nb767Y8DlZGd15V0m5uIeAmyygjjKMRsUPi44vt+
CKqF3eIHYGFzyTprAysZbVSConmbYuNBgrjy/425Tsw/iP9K7UsECrUfDYl5z1yL
JkTknQ/YRj4YLz5ni54vyNVjg2kTmyiBuVjNCLTbe0JmTIQV+1cgXyuHBmnLqt+D
Ot2KStxzJgbYsyTKovaWgGTFzSLmoOfAEPBwDCAXuhExWSWYL+0BnDZd1bIqeQwC
/tJOM3GDaI7G9RygHS+NnkxcGwjqL+IAvTu+3jfAmOtHtKl0NHiJQjVcUHSbASgf
W4m4ZO/QC2thuVDdbU2OPQm7zG13xNA+rxCFGR7p3PMGZKjiqPs/UcdIJ5YZrf8T
H7IWoJ0nmPDXZSBnAlEUdZbPwbggAuOIqh3gHvOd7f5/pv0wjZOqWecPAADS4u2m
VLr025japBIQKM8P9aNsY85B3lECGbCBmaMZmvKtLUDEbYqt5cBNJnJ3U70abpBo
2Z4TbR/hRa1p0do963D6rMoIhfe0pJHRbxrpC4x+OFHruLLlWLYE+LShPd76V0mt
KCwAl8+3+JQ+FAJ+fKSES4vCNxEy963BjPmCOQPYJuqyFYpgU82MI8bLAaehPDZU
0xrg3bHbNMI2as/JVoCxsWVva4ZXz2WeG3kh63koPLgpe99rWyagi5acbJ4zr8s0
1tikEilLapmVkUxdPbcyPfOHCpZbWYGC4blI3R9CFmVo1eVXTQFCgfqgv4hp6JQG
7mlmMnXdwBsRdL1ODZ22Vlo8AnoVULo2QAt8/AZXOzTs7ovXeDv6ibmWiDzJK+xN
9NzifttsDOabOF/drGlLHHL4/m5jLBM2IdW8qWmHLdB/TNadVfUJV+aVl5Sir6Bs
wSyVI7zfKXT2KPkYT6Vp7eLu5mzso2IPxjkgOAHYinT/c8tr9HepriBoYPA2R3Fj
pLSAXIRb7u2HexZ68kkrC2EEM8jkmPteCPu0KqJs02xu5f0z1tpwIYoe5EmMR0AG
mQuSTkVpMx1APV8oVxujiSYvCvTjm8Pk/PBySl1BSJuxK0zraoK1rJs6nFXYa9aD
3mELYJnkb/BKl11P1fGB/u4rkn3ur1I4qOCnYVW2gxQyVsE+yLP/TGZmsr079WmY
9s09WKjeg+8AD6MeQuAuclPdTZwazl4YoO6IkOepb7UThazYwEZ+KE6pmYfo+vo4
uaIqa7pks7EFRhQbDowIRtSXEW4GnRnkmJSA3U1uStDQ6f0LCBGheI14VfNzSqzT
gFNQhX6T2YgjvxR2xM+486UYf7tKHkvxvmpxeTfFpPG9hxWfzfSt4btLYQvRdxxB
7ORWrKJFdhpzaXsBfzbX9Qx7TclCXoRO7+B5uc8H3cwBhGGm/k+kTDSeMIB0lYcF
57lSg1PGZyGnvAWc8m79AIcR67IeeLF+0ATjXIUFulp/PrylvsUaeLtXddlx6yRP
l/6EXk1sTHukiN+H/GcuspUOT2+hbYWojDwzCT+1ZQICBUDylD4YE6WR+epe3qi7
QjLqrZt8Wdx/MIjZCny6q2NY9B62kPZmRTg5AfnkGKRGm1Mo+jHAQ3Ew8rLK4a+V
kio+1fE11f8uHEVYzuGqqrjeOu1o3/fxavp+bcYg/QtDMP7AziVAYLAOA1p1oP4a
nx94sQDlcm5//bhl+NsHnwkg5uvpTMF7GiHLbu9RPbmyVM3dk1m6Fo/PGXr7+p++
p1zjSpW8e2pG5lUhP8TfMg9wAhNR70qFvIfsZBjkmNl/BZmivY6lMRj+3tNJDPyw
5aicCnEXqRV+ZT4/sSLwqlOhHZbVaNJCnsn2PwIe1lp6sCautonctKJOvANj9DQJ
tUzKyJm3IApZL5q9BBu5dfxbqUJ7tkraPeEy66piTZAWsN4Y+eprVon/NxsqRTel
k2taidcG0RS3iOpzY0Zu0/Q0Fveb4UN0WcHMbirZEpM71UYLClS/udXnPVHVqrmX
bbBSasUGKNJc7wk5Z0IX60Jo8XMMrdqj0thVXaylleigXTlzgpRipDtZJe4lgwUX
r95XqG4q0ffE/vXSsp0A9vUgfvnmmehN9XAGo8sfexK7A8AaGzKPns+I6Hq0dVGQ
DTKwWx7HNW5O+xHlEzqdvuCMYxrsQa7pcvJM6yslJMLZnpEWD0F5JY0hsq+Dnmiw
aSn7824E0WdZEWxo5y0w4NcTf5plfJKxvCFOZbmQdBH6JPtJJ1UkpeCT6RbOYwlx
6WEB8hJ873xjEEBLDe0X5FqR3QSwio7KkqT7Wyfg7cKk7tszY7iPLZv2XVwd6821
RZvxrHtDOEL7m/qwqGfoG4vgH9mE4IyTN8pVDky67gFE+5RmUzkP+tmNCcL/m0LX
trGj47kmivVd4Al6aQ8KpkKCgtNoD3qIAl6WKWi2vd1qh/ThYz00520YDrGGktKK
gtCbT1qI2Jax8NJnyW51/HGI95hO8x+BtqGX+01PqWRSj6+Y2fQB8dRQwpxpcsk3
kKeVhOJR6zJy5HOmTYZCVvxX1Pa3ce1jz13rS7oxaXCDZcjrghD87yBy/Vy3L0QL
/WUUBxpyEqejTywWGtDB3dGOQYPxBj98NakWh2SVH8xCaaFrlV+reJXyxJE/1f3x
aNDMUyGH6OKEQrip8RD+sPrAq+jtyI5OfgH0IrP8ZntSAhVDD6w8xoUiOzG962gQ
9aYNIaUtWCY/kLNPmpNMmrAf3qCCS92de66Q9ua55vNBOwLtiTD/VbqTJCszl21K
dCJcx1iFnq9uo/4v1W0AvvoeUONe6cQ5o0Ex0xaomNdUH+sh7iMcr+DqnWkDUR3d
+TMdK6CAK/du7o9CeDfZlKpORoJhIACeJTQjUaPf3izAjRH61pSTgOnZmV4N9BsJ
aWpJYk/pXPW3j9mNbltFMB7PX99jvXvLAQidxsVQKxSL/Pvh5RU1JSF1rKUqmY+j
IxtbCzCZcRk6NzdAQ80I6lruZZn1ITxaviSuqKT1QIwlLuqLZB67eHSs375nQvgp
PZPertMg/PrWggmZzTlh5G4xtytsIExSTF3dT/x54hVA+cHYuptUl9anneRVrPKa
xOn23heI5us4zxo2STAruFOpg01hgyGRbnAdJ3OkaUagv+bTiiyj0D1rQPfHU7Ht
r2+dHKx/vqnaEEMFeWFLGfbC7M6ZBXku11Np1BVkjlaERVPzlp9JKcJqRSBkN+84
+w40ovvywlgkIAz2J1F4cT6jY8Rpw1OX82sWEfloUvU7dzBZTC8M5gnv0fgaE4sE
JhH0zD2ejeuCo/BGV+ofAwue+07stkSohcwHi6MMUtzxEDMkg1fTr5/AUW/7YWuI
yXTJN5f0K5T5WyKis58fy0FVTJxz5M0vqZMWjfchUnJr67ImmiK7+HjssjSx+0PB
WlHjf5iGsmAXjSH8mh/jrWq1aLeIJjYadImk2wG3KW1zVtUpzluC6bjCql8O2Mqv
INcnHyXP8EHbpLJl+ku6d4ItBjw6wsHKZi10N9IgLoYLn1UDu9lQ887BieNKVCNE
raswrkgJi/vAschC8tN5/NqhE8GUcc751zqGg5ULRBT4iPh1VUS+1cR5JNPe2gXC
EybjiKRJKO2WcemjNPSqFpy4C964aYQsrrRIIL4Ms+TQY0CZsFvUrutAbZF/gH0Z
Dx04DVdVCcgjS4TRv4TesIqCyJfyfi3O6FzoZs6gaMlNWWNiDstn9PgvBC7iCven
ZOS2iygT733JN9y11joRQ2amc0FI28DILI4tSvc+KGmyFNER0PS9AbdlrUo8cIIh
scxnFekY4psxYAUHcO0Fqsm8OS5K28U0f7Bok8xOug723Nca3pIOw4/4FUOlzcng
UhTovXrEHkuypWou3j63s3hXZQvnukiUBB8FQQBqohJQmZ4Ak7OFejQgT0ILsbAu
FyaHhojz4oRhNsh8ZMc4RJWXh6GUdRrXHS8GrNwaKhEWdXyJLbFCi90pJP+PtnJm
x+V87unFmcyOs1rbW5BlZDE4SqGYHh9zPpgBNsMxQr4Fy86vJz0AC5yppHlOcAvI
S2hRMmgTUjehhcDQz4lRyBlFFyi3wk/P6rgaeGU+U8XvYW5XHrS2gwyfQZqhr51g
CYnaJc1ijrid2wyrt75wdmai9Jvuk/BvYuBc4ZbxWxX7nxasfrvdPipsqfl4Zy1Y
PDEvRbGM33pziGr9OMV04SUlG775DmtoaGBbCKRGC9ZeaxDMkAGilTt46RI5ND3W
5UZXIP6cYu6pkauR3dlo4TlDlv9Dhl6NhFftBhRAd0hvP6dfW0H7QrXj1TG1fU85
FRjJGhUhyLjZZ+h8GizUsLGlrHcnWKzU7/IqHCKvd+M3W8vAaWmfmqEoy41FLQh7
96e9qxnbynN7t7RoIpg5Trxa1hNIPtSExmip4Pze7n27N0oOYOBMqnZtNiJ+MfmG
vRl/ZlPB2dwaNnSw+TWqQL5NnYfQQY3PeujZlntwnUnbauj64wD7yPQz04MRiSlQ
s8/wa0/PWdtdbmuXLi9xTwmJWu/V79ZEQa3799/voEV/vbudnG1E1S6f+A+04jFc
EjmzLhzO9AnB6kBVxPqn1vTQU2RTSLbllypVkfXP94VAM+DxQm0ZBy/ZfOtvvssv
24Ql5Hqt0gdIRiZDCEvbZXvT/I0fR67i9Sv63LM0AXe2/0llrslAn0fjsQ1T2mMF
7rkRBG5ThKnPuQn/p2qUNJDzzkMrdUXKAeCLTGCGmGF/8LJ0gRnfwynRlxafFULt
RC4IoG1I78W4dTsqt3DHGJhi842YXkVVhtKGsd61Dh9OWBHcZF8QTo7BN6EJN6or
2gGh0r57eVqlLnfXw5OM1yuj2szG1sDwhibFLlfV2lhrZ1ww1wJdVkeVrrZpBuQO
7tky54GKGg/V03+EAWfIC8ErI5j0iwjuFM+sKaGCp1Y9RuzkFtl1xsu7JIJU1qcb
0OI2M9/rx+QJbnC64eDn7O+hg+LHH9/GtT5gj4X1JtV1mXgb2peuOyOmx3nj2Kf7
Yt4DaKHxj9ebo/GkqDqfO4+vQ0j7R/afh6aOHKwwsK/P/8VlFbXOF+9ETO6bW2Tl
B1e85rSivbcIbBJppXa9zfJCGz5RGJ9W5UH2Uuj9h5rPi60ioFsV5YOr6OdpC+xi
SPQh8Iq942XmomSroUHtRwyHRqz/Rlxe4ulo83MYdfRbUpzOOAJM1ktw230hC6NX
U0c2myc2I+21ippHEzqP6h85zS13cLVs0VCU6tSPmwWUNXQ9pZ87eKYXAzR2ssHU
fpQrXtT6Z+tGvxlUw2bITEowKLTF037smNcAPXM75eGDekw4IahGGU+7eSF0ZGrm
QQyh4dh7w57cwA1NcDCF+F4TfcTtnvQrnbZvNWPOb4fcN141VBTlxZJJUupLeBlI
ZMtiCAHymZViGxUJCp/5lUyTVCuhMT5zFP8MZZtyqfnEM5EOY4/KtLpMGARQfElP
OkqGitr/62l0WiVV5kO3ncDBpTZcYWZvWhHx8GqtDvkG/fNogPlMrmYFu/+Da7jp
Wj0SxAB8+7OPVYVquFx3oOjw07h75dEv8N+3KNbT9DNSh4qLbI8NHHGbnx7IlUC6
yylnZ1VAUt8+FbVqDRXO85ebKihUK3AcrKK9NkeOgEyI1yfzxF82Xd6A0oGi9kCq
M4grS8555ifsar7v2TNeCg5pGJcaA6oJuaa+gPW/Zl7dr5NrAeMIasQFfOpe+AQj
ILgG5+sAC1B49+w7dGKBJlNEPg0I05Zp2pff4qSD+fjVPHfrp3E/uz1akust7C//
TuKpph32+HWnBZB7uns2zOnAgCsODxeoRmv/bepBHoTu05yb8qvxyH6WkQ+lBLPk
0gox+noJepW+afWcpea3B3ozzRmqVdSoI7qkmT8m6TX0Y52/IFiQ103q1ZUSFDB8
1kQm1ujdPjki4afsdjicHtmvzarqqRvMSN+j2P0Tt8wdUhvL3fvCT7nu7LGluNDp
2x1CLa3TuZnekIkzqL25h6OqMGGvm6dZuGOubeaiJ+EbWRvUuuOybz6dh4NMkobu
JGEsnSToF4zXBDG7kFXPLIQsHPFC/8dnq19WShF8wt/5HyYGsrZ54znm8kVtutaU
8f1TKOoIMI17iTZGqSSgK6iLczgNYsxOQYM+YGcN8gyAgv6OTGmRfwLl9RsNK69r
aurssxxmgjmeoK0GNbbKgIAPuHZ8sW9BQz8CWIPCNDndiwvSJiXqIHZSnmQN5l/P
l+fw7dLE02mD+74WUkKteKAiF5Xnb3D68TL1tOgSbghSuhPjh56ZJY4HBpA7jB86
E7OOkdbopYb6aGvTyD2UQGwbDWuClPtuBGhqOSwjTy68/KI8jE0dNo5nqtjaOBqq
LgLQfaeJXfICvqf1VvSloOJkY1EQbmnqeTR/BAvDboMix8pxk+ZZh6p29lMq+i90
VEB/ne3+/8r/elj6e8IihdKGtTg9E2mw6TcB8uo6w4lNxtaFV41D2KU9Qng6ABR4
vbq8Z1DSdBmbn76dxgRufSnSS5gBwgGJpSeNFAm4YllHlGFCfF0JTwfiKAyjLgVU
w+ODcrne5+WbnWCN5e03EgJZON4Lkbrz/1b5jq+Wm3uABfnkH+/rrmui6cOUlQuh
Ijhw0wslV4KKoLBZoYx064x9RTq1eIqSsyvPQR3xZW7ZBuXLZ0+cmVvHQpo/AfrN
gs7BqQ6mdr3e9fY4xFPAMsjA11OUXMaVCC8YZMPxzwrlhroA9YJ1hiuj/d42RtD2
kNqBd3vyZWLm1RhFHgNOfkCUSQenf5NBNwM/saDgGLMWt13Hp+GK+Ka41WS1L+M/
NNudAypn3NeJrEB2Pt11yd0UokwWmcvBbR6S766Wln4OWzQ7ikMQ0Vv6ph0TIfAh
8/p7znQHwbsp4jKXQ8YGqoOQV0/OrUyBRXUrwVWQqfga11X/auk7UIJvf/gWgkLM
orB7GMSufet6Qba/018Fvj7RxdXnGFdblhrjXVvybvULB4yeWHvBaj1aFTvQe3qW
5vby6W5bLOSY79PTJDsvj/EH0SrZta/uzS72nIkG7tL8JffHeiteeGrbWKFexpix
B7c2IeCRkc+AK1NzNBPi0dMsrau3PpZ+LrkP3G2DNUE8TaGXw5d/8dT8E/KSCz94
rq25bSJtNa1U3oeJ2U6Hnyi1fNXBmll4DIcje7e9zpsOJSrhY7PLDEKSBLwdUet9
7t0zfP23iP5zdJ+Di5M4Z561SEZ6HrDfv+hBgGyBgjSUg5ZRueAR0Ybgyi9qxeS0
a4MHC7FRfvOZncccH0MISIHvX+M4+jOAFqQoYsyutZuHRJHNGTNsf8JwEhT0YyFl
aLd5u01ORroNnUTYP5bLfspKCf50UJWbnzQdl9GWeWLHNhp93fnR/Q95Zj0qmg7o
UUIZZex8m6Snz4GtQ9ZCSE0x6xPIN3IO7W+gePFWvyDcCmbcohETIdFUHfwEiYgg
azz6HVQmEEHmWsm0wLTufQnnwx99dyPM/aGPcdqo77suK3ldIEDeI5UpmqW+xND/
2777lvjPkPBWVFYas/E+oY6Pxvf7BkA1jsNdF6QU2l7kN9hQIi5Bo9EQhEuCs2cy
8ccVzxebJxOjFFxiusqz5zSJddBdXMfDV/0IKYk+LMqD8ORpYDcAw94jqoyJYfMf
VTjSdMWjHe18xUA6HnpR4S+bUSw2QAu5Zs6J9neqjhQ42bY4UNvzhDanTIz/RA9C
v8SJvpv6dAiwa2cOxgooy8XOq3/6ax6gduLq3Xp0IkYFb+1RvwDconI288dG443T
KuU7WjkTnu4+pHC7ys0FnclQy6oDeG0luJ4JbCU8W+PNMN344BJIUrKEGNeKlIk3
TUc2nzo+cRL60TUmtxVwco2vngI/HZxDtnf+sD4TtnDYMyfCkoqtunyZ3tihzL0V
hJw1NHD8mcwc4l+8wENJcHwqWr/pFjVu4HrxHKJQqvyCIuh5klzSF8MFusaHItbb
PV6p1UyvxioYwEBGD/PUpumQAiIK3NNxT8MtanAbd1zTaqulJFgredz17755athK
xcjiGGkw60wttZ6cQ0eXhXM4tfai3810D5bUaN+NoBK7dUboVmS+kiTxGT7gcDrG
fy6UFq2a0L8XvPKEHXSx94nPVGoEX6x9e2SGNpAjPlBgN+YCivCtBqrQw4YfeB/3
rSXCwWMvvOo1WBf63WRETs6dusT0OE8QMr6eSofycBOOxAswfSCmLYsj2oalFGtJ
kuF/eArmgZY/JPjuEYtEiOzBbq8lO0mq1pgg/PXN1n4qjg4slfDnZ4eAC3EWfxBI
mMQcrm7DGbllu1DawdvIDf3cp40nwN6/ziKJpjSVsQoe7sD2VroUDmXpd2NpEUUg
Z6UqF2Qrhxa4XKFEv/Pn7jRCOaXPSlJWydpg5JAj9lKQJzCm6Qr4g9BqWYvY7trV
wjd7ecgBvH21vXWJXUxcvDISOiTSkm0PdsYodwPLHRexPL0Ixhp/yjYtmXxYrlJt
7xPx/iN8DekA4smnaHWKljkDQON+1DbTs6zEalUbNS/88o+2m2bNqAYeYtoj+gi/
Ppd9LTPm+MU98g0VUJotwo2AGoLRZdDJhzYy5vDgzzBQqAaEq5pDmvopW/ZkO+II
ksVeYJgY61nLECGk/jfBoBpiapwuMU2o68fKfwze/4RaOsf3z+NgU1yOYJGJjHpC
5/QBn+xYXpKVZj0KSbjdDOisSBH/ZTgx6ZIA41It2l4ANULigZEzZ1qVgumXWiZB
Brl0NcHq4/f8MA3eUdfuKrGIzWum9Y3ROXWTOwRh8XI=
`protect end_protected