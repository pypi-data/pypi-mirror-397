`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
zZSxD+gXg/oJR5jdsH5AQ5SDhL3kRNjCCzaK6/Ky5pRKOo+y3tMZh3xoDCuVd0Yv
H6STfAdEGRF1vKQlSbvbcvI4WtpH77Shk6p54ZLcfZaS8pVj0f77QPzzsJpL52+8
34xYH82nQRIynsBYCYYS62tbaDTbz42WY2HEEKVcPYBrYyEsgVrzqHAIjrE0jd1X
iJ8HWR42JUtDD9zG9TT0+BKFLp4Ow8218ahD8pr4smbNwi+j9KHl5zCOv9SoHwA0
q/AkjnVLH3VMW2YkiVURGTbuvoPge05beEVTRfM8tlLK84OcW53t7+9joSJY4ldR
3QDDZrPbIA4GMewIzBUD43MyPzYFBVPplWFgVfIBr3xlySGRfgkUHwp+5+n1Shhs
dIQ6SV9zI2An0aPOCTJbJ/NCYbkW0u2SRNkk70iGrGRAbh0J+mbH6B8M0NKilL4x
EnJjbAw0mFCYvZcuNOCzcFHt/WLAo8YgBU6PEPYcGokMO7qQpKzSuSYFgryVgNDq
6Uj+vqPsiy9ZnCjsGCPxLgXwJp4qSbLPPW7C+Iou19m4QAu2o4bUH2hsCFFHjfQn
TWyOg0FlyiiksEZBU+gNU91nPVkmNsSgs0LeNwbHrtS8Q00190rjrvCUs+kvWR5C
dRF6g96SdWir+lgKgxaNQ/NafYCk3wpXSwL9dkmO21kk4HSfux4ygDEbnuEEeMnm
KCkNk1Ie1dGSmR37Q/LuMWH+qQPAn5TrpvpfKTOpw+r7YavQsquTK6B89rMAjYyS
rI9f/9pnJT5JWItd6Xb9OK8j6GxZY+mqNz2KeGMmDJpQTs1pSK7VeiUvK1khwR8k
Db/cref3Ge39NT8AofqAGgxMkD5mCo7FgQcPGTret/SSgXT0oBCVfqw/YheIQRJv
4nsvZ2gGIIlTVF6/S7zpzV89eq5oR4rOaZQtLvTSwFKAlyYFsn5cOcOIg3kiHple
2OmfeLpX02i6h6LuaQ6UX+l0UYmMCq70BFpJwjYJa2kNE8BhymsHogGmf3Br5EXG
7EymvT5h//dKN9mjjLcpAYr0zypKNqNkzIceZRga06N5ZAZ9uu0LK4PqUVPZquT+
hKEm97Pju/aYr04rGoiYKlAQpVZP0yXKt3IPiyYuTPJnBNbe0gyIIrQFIgBUFsL/
D46dNA0LjvTfuvymBZpttBvxUboYR3nCoVN0BJCn4nHHuUTSlssh3+I/5C4KCIMZ
tQ6YW9PAyse565ojYcnxciedWmXeVrSW17zxB2CVkm6mE5clNcCHPdvLqTefBzsE
c4k/xfNbfkGKx9Q5WeX6V0mvbNfCAdcsO/bHnZDYnuXH4Yt/WI3Wo6HY3cig7jCB
uiP7BGaviSw0SYaa2bjxrlBJaWS+BooCLR7Umam/f9CVyaU58GeNhzu3O5wjhVM4
dM1fNuIFJX+sAQK1OZcPkCOsKNwLIH0jkA6k78BjhHFAG2GpH492QL/vNa6dhE/W
nrUkpHm9GC04bzyz7G6YZ/fPRTT7zf3aSuVL8+QXzJLPGdW5YTn6UoDyHbSlHnTM
EufajgiyWWthxboojXSUuGci76L7Zec6/AZi1sYs6we63SPcy9j1n5DdQYCPZ65K
BfePce9IRbrwFN/cQorTi0rNTCHtdebEXF+RkkBJ2612ptf1uMYo9i1D+xeJwzQ4
vM3HmhQRpenNGpfs6scpQIlZhsi/XQ9//VhomtPOrNFX6EdTlMSrFzFzU0OTP0qe
CdhyELf0f4TdSMqCLESYdSQc16A7yLKgHt2O7ULIbT0jeVygOR8dcHemz+88+Rke
pogYSvCcveMCbTLATLgVTEszQkAVsf/90bYE9O21FRjFCsaU3B6+VGouGfYC5eiN
GGsquf8NuehFTREkqzECFIlciB+OyI05U37g48uhszOMOp53UUzdgHYhmfDcg4MN
MDfBLzGMNXhpjo9/lexTfHgtTbxiu2hc+RcGpXg82AiZ+HspM3ewggdhMOkOpFXm
A6cspgEpFVOfUahIhjzMN447nC8fcTYempAEQ0NnzsxtBZhecomlYWwfmJ1gm+HW
6VdT2PuDulNoZ8o2GupnoPbtIKu1/HYcfRHUaUZSAdO0w6PdL6Gd+DVi0QdiCJfw
/6cvWmi+Rw+2PM8DKi21Mg2tX/CbcmowYSRuRSY7Q/ycTdgQIE0ao4CN3IrWYe48
4Rsvb9pDYky8j8rFbX1lF2hEbgZ79IrbBaNmVr3408ymLwbTuQKpU3IckA+eparw
h0s4Ep+R4yUv5UvjPfylueJh8CUYSLe1eIZYUYRyKsOL6wVo7caHLfwKgTWxXcCQ
NWVG3nqRAnPA+IN0e9OxXFPBy6SvDWX0TBEl1dJzgkXAf9MZuIZ4Vt/foKJLwLGD
7lvd9qQoyOrm8Bwqe6qIRtkSJcB3wjNGqknoqCADJaAVI5us57GErrBvcuc5mEY0
fPMStWqj0SmfeAmDwyZgu1Soq/cI3S/pipYnsKYltEsnNuwrBT0mV5LX7D8NRaGN
iDVbqWr/xYbpdozrTXPvugIAZ47n8vr9/WZBhNLOLap4x/JpQQpJZ7EJRBVIr0fk
DlNKYQw8pkle5x3TI0Y3r0uy0A1w8UVvtS2c7dJoSBKte3j27t+jkgj06vgcvbk0
TWRpxf1aBXHGbWVInJ8pPLbNX5eOuvjFO2wdrXD9CItjNx+rgEwplrrSdKFkttr4
ZUbjpQGBlq6rWqbYz1YhyslRU1nLpPfkzWbVnEX3bVffX8TJLuROTrwuUUHtx8u6
wXwjFsiE2R5c+XcySXfeU35yNEdgvJiczGsVlhUMr+e71y2ctk2BLr/onq0Niovy
WWuS/vTcv6Xh1ZXf3mKR7GiuVrmdQO1o5dRaIrbi57DbSdkVicdnraoYmdFGGObf
DsePXfs+oq5D01JxrbtwwtyzBQWQXfX9NFtsDeReFZs1iUd3ivqYPoqPhTmyOmyZ
Np/tTHbKtE4J7I0qsIOl/bobf5RDyryIGm3yMd4T6JKnSUFQyEezDJtC/+RVncJv
UuJbkQlqTQLeRQRxJyUR0wCzNRwT4GPJyzFZsiwaVmkv2ZStqp8xIyC/A8sokNzU
lyeJzy5ghnTRgKGanAnibvoBo5x9p7qnwWOzhUQeW5Kmtv+oEfhwvCduvSfV6RpD
JmfXydmVnLiJr4bsZldwDmfUntkpGtTmog332sWPKw9jx7N3R9HgkafTBv+T8kMF
tupoIcTKst3tgUiGWvyZeMY8zVLAXnpcreyuPBBJ5GAodpAUiar/ciUUHqUJlCKt
QJy3R5i6jXUWqO0EnIZ2lOOfFaDDq4qAEB5QP68/AtF9967uaseP6XA8ktSjUfWP
8KLkhMlilM6qv1ZINibmykCRfy4tEeB7r9m4h5xNASvXfQdnsMArrDY2aBWIIV9E
dDvuhTs1U1MckWVZHEA1VD6EScnax9p/6RsEXos1zpLf84AMr2URUgFDR/jknD7R
05QAi9o1PQN86wXcDkU6KVCEIDrgypKT1fPmy4OJQGkkH9/+Xmo/FW+TfFj6g7+C
R8riD+SU96JV1tLskb29av1wV2eepb/U+lUdV9oppxpAOlhQ+JvIE4X0j/xEdpQf
yR7nxvKr50uj4ozN15EThVS0gMGzyxWoGHYUYLB/AVkp6BBU7+DdqpuniGcD9SEB
bhxF+XA2zbyLphPt6sScJn8Nq6Ih2XAUr4hRdTfDXGaMYFe7++WHHPuJJCIYtScv
wLzKzjDmCdxcISjh8SsnvmiTB+HZ18vpF7e1A2365cO2+XXH9/QWWzQinr/VhAMy
YmV8MEGSAsZLBKBcCTgWjXJgFG6ZQCAlhYaujohU6DdJd/HIVnmv2T71SXobRkVi
ZDg3UVFC1rFxdfWAJTt4TbRZVkW4Pz9R1CjCwknIv5ZpoIufr/oNQRzJbCpZcW0n
6Lsw23Ud4MaQnEaR9UmJXirW/J7SdIrd0zZsTbIxzNWzenpm8ec6XJw5ZfN6cQfo
M4nLI+7OVvvFfi7hMdjtUp+jEac//bNjGcVeDr09TFNcylZ7vAYlhIw1bctYL8w/
+Mh8LYm5r+CrPPzQmjWnom6UvIIJ5zi2TqlY+89ZWeyGtYLQ+n4Ho7yUIg2XOIZo
oLP+AKN5d789RYly9atnZNWObAqQjxhuwNaachZX6bAeGBnDqUoMQDeCRI3e4FcW
kuqnQDFP4NuFmYeM73BYcuxVAPl6fllvcVgmBypiLKCbXWNIqQxXiN1E+tjXEzXA
gcNuLVCVcaTjIrlAhV76buDn84N3l1+/dwmYynvkmv0GVByi4ntAIUyuMc7w4Nt0
0jlPizJ/gmQsv0wMyxEOSELfYWxU73dsPCfHB3gKBw49ZqcMMYorl1ppl5zJgazd
+34IeRz7VlEW30s+Wt9DJYWnMJ8tWpQ3eKctmv8fXqYiIldeuwb420XOItjJA0m2
ufPdDrRGcAh7hz64JaOqf9dZheSZwbwpKHSajtW+qrVRdxPnRZmf+PtjyDVrAxpH
gd4HjcT6GSkBVF5tclGwntXb9FpHFLZ98/dzTS95hcTSCTFNBT5034wna3KXwdgh
JBVEgfYQeL0oDvx9K6j1p99g472ZySp26gFrrkXuWRJIRIeFdiRuQzph+rxcfNpS
pnRzRXtNtSHqDJXVWondTrFGy5w0Cna+D4RawKq5yn7z0ekfSJ1sEROKjnOuaUWH
Sm5NxjEtaU23vm+100DkI7wEl/pPPyIhnyfJ4WbK/CVXt7T1gtjOP/RAmFElG0J7
tl6cfevyaKwM8049EKCu+Mfl6REuSBREN8I6JS/c/BkspJfPAB4MY8k0thRMylkJ
OdoVOZk7/q0N9MryeDwdRzwAcfOkz1kVEryikqNiGx6962jxkJRVNVbuMRm5pc99
kTY6F3NvuAreLEU9t0QBKrtO+qo917DSL4bLQQWy6UPu1VPXQxZHr567DB+L3y/d
uLbvLq2cRXpUwJJ271f7/hwTYCfHjUY86jg8ORvJbphoY5GQnC67EQM5DinuJCUb
8y3HWa+fjoPMb6/3PfRLkHl+spxFs53bE6J8RtsayOPFx6mpkA7AjsJ0l2FVNj50
IEdpiK2wLbpn8RrU+hKr0cuDpIMK6kGwmB4LqH9ePyfpVOqgV0cRGT43x44w3m9N
DgBAWO5fUxVZIiFmB3Ryb6tGVOEOt8yZp6QIro3wiqpsiae0jKc2Fv41OtI8v3h7
9iZHM6IBChyIA7OHTRwACyBFuyBxz6NSp7eB4usRW3Uqng+1W7Y9or5DDP3fsdgG
D1xPCycBY8Soaxeq7jhBCBEy0db3Is2n+sA9L02H0RmqmEyzORMXB/boz4gBtHDa
hg7s2ch2qLHJDmR8n6nqU7P64S4PaTKlLOoOHIq/muP9RWId96ag/qSyAFyAVWRR
LgDl29BZIgMlA8fVetrSETtegQUuakSQHXmU7K8a/VaqD9k2ZREsKTAP19JCeb+p
A+JzsgwSTkP1HeU/+Nd9eH4ogtHCnY7UIsu05QiM5AmuPKOHePPJtg3xjKeM3yoS
fLw9aeZ7AsI/0EHiq4AlX7RwXRu/r9kadxdB7GQsekk44SGCcyL3xFC9kAb7Z+9Q
ljGQTbCRTWlsqGnvbYs325Y+Nm5mpURXe7uT0v5+nQNTH1+71Iz4N/x4TYw9QP2U
6NcvOpTy3bzukE5O21BpqsQVoSDoXkSpPMs/U9sd2pP1707hUJOvinNzxUwCLLXW
J/eWDMrl0rAQRzLeroLpYN/BgCHLN3HxMkbAbI4QidPJ/KEnNT3CfMDCOVREHkgB
wEF26/zlucFCeokVEhSGiXqYocbBQkPaHDoQBVc+/J8aIntEV0uudYEci3+vZRaV
sjNbCHT3WIOPah0NeJzQr6nCVBkURg0PgHBxjpm/YnG/H7JRGvVR+4JWqcPk8AXg
kOvQbcNCzjyJ0RqqzBGaTD/fOET6meaAYu01O8WXLVVpuzGgcVVPUHPCG5x6pZ/g
3YPsVAFRBfSjKBauZ4KR5G8bvVGoddWLi9FAB225bJ1luJMDZ8makHLeybTeRXW5
+p2qGq1PXOspmZ7NGaS9OGMAv0lSuXIrPixUl4vwCDRlGYAi+ym3NB99m+uuL1ON
86OVX3AUSoXTFIyVJjjSlTqlphg9h/pn1SpvSyICaFf7AGRJMmP0J86gtm/0wMaW
M4tqHmrRoCIcde5mb6MIbc8qdIMEZ/yXaxoLTClJ/K0Ee3jF1H17KDnvCRUcigvV
cZBmTlztZ4EHSzmCzSet7spKgHe2lDvMQ7iv2F1B6DCvddI4w9e6+ejszyMMyIiP
xBJP+dJVIo/Azn9vTvTET5szmMUDmk5usnoYwY+jGXX3Wt6RN95Z9EwWsjr127az
Zr5qyqdzNMg233uutanW0bvgj4AjEpr+0PjgC2BQljUMjfh0eLuxkd5WMEfo+RR1
PcfKrkGHemBr0yrEuh6pgAiMinxZrz3THhPC/5BCHkZS5g16PNQ3iGPckjTCyAN8
uDnLk82m3+Edd48/9M133IC2u5RZkOisTpbPBQ7fj/hG+PNwVZ69ElMj369X98WI
Tx60nRD9LzRzl8TLij/+By0GyF/pEZK8colE4Bo6zHnHFDAz8hXVhy1HQ45Fqi2b
indWFoxcADlROCnS6OLGk6SAPpQ/xJIIrZ+iz9ws/WE72GbjsiDobz8wTIsfpGBu
TIrrghsnMioRLEPEyz5Rgi2GpJJquK3MZykUBraiJP7hHMtiNPNFoRePZQMxlNID
s5bMXfPM3oQm0lbHdaW1cC0962ix3vNnrvmw0RjeXDailH/7RhKhY3b+PxY3BkGy
Uw6pEyYCaMGP9E05vzr/ob35s4v/71qeNtFrW+6UslUbkrJg+7gAsP+cVx8LA4mS
+qCU/Eo4nljSTaSvTqb2YUw8MuIuJUEd81obtF/5EqHm03oTFmd697gY3owX35md
oDYy7EvWSPk0CU6pMjcbIO62vdGLktXKximRU6p1luvmTFssphUKJw85iJR/EzeR
YgdclZyo+Bxr+ljBeO6GLmvlKX4elKSDHoCxb/MJ+jMiYPKZg2YO/kXf6co2ql31
Ombbcv/T/QBqg+EXhfkXI/4zyFPvmkXgklsjAmTgBOBaiPeVU2IuCK2WCtET4aJg
4ShULGRQcVFHGQ1EZNAGRfKozQ86kD8JEs/v4/uG7Jo40V3/16KeGusUtGxHIRzb
P7q5fkG6TnHXOdL7bEQ4zVtrkZUREVj87gTAOvSlP5hwQmVmoNxTtT9F5DpVZYxK
wxjwyFnFs/7EwZgYZAQWndnkPMfUUSzw29E4nZ2v0Sc6QkfT7vIqViYxCIt398zt
jO9OHh9raWza7JGWeAuZJe3thykXieuHBnWDG/GBZr8abw5FHf7fhvtcwcUd2Fzd
9dcI0wkv35KPCOd+dOzX96fapk2naIIUJgVeMTFVCwp6S4B4eL/UzPw9RiSvhkwF
kKbJ7YvRjhOniK/QJ32VIVJD9TlR1XVJbPyGu7pkSIzxFeSW8iByhxXNIvH5hsbF
O9h6sP6gadLYfcisz+b/LF0TRnDhQZhTglnOq16PohtNR+4Eh3cyTF/2hGZgcSxp
wQoLflMJvQLzWPqy87BRS4mZ+ouvQr3edHTEEbc0JqJ0grGzrLYyhv3Nvvs9oCGI
nY0ZPiHZMP/8MpABKegbgj3FiTflcjlDaacnQb7S/9nzxKN1HOqNQj2/ADaql9Sc
1Jke5naTN2BPLCBjKr4U1j8iGPfcAvsoS9erRr0debYvEGKXs+MtTBFreALf9zeS
tf1Nw80K8lv31Ko27BtmIiUefrWCFlYgUvRn3EzoQETxr/HAet1Zc7YJMICCzHb3
BjwT32gXoCNsyHlHyWYLJlw0+AOT2YzUyShQVvjMJ/bvneEJ3Vaw4vAtgOmmZ4T1
enQFyf58jgYyc5huW9EcpdskZX4SYSfqQh7wZy6klSWiCeLp1ov75ip90lsWM9De
4yJZj0ImMghDbgw7DCXqGBbe8bft06LFeN7enL0IPAncqRmzN5yvLFtsocDByJgB
HbJOc70m+iH/tGmlMWDZq8TXsuc4bbCSQl5Om2KrxcXeahfVsMc9o35sItPwjSos
Ti1IqN2exyonAUDG+8tkBHMSexnXtBzlW0tNH3dl3lGmUUxMOLnfmXhygCJHROXg
MMu8YPl+GQAY1zJqXNtnbs3w1id7aUXfAtRNg0XiAaHWPypwSMJdb9X2JqK6rIad
BmS7/qZdwfP2oCMJWBPYxiqwwRNVcEr+MCOviBzOT/HlJoQvYfjWbmGK8t/KnTBt
L9vGTSEuNWyXzmnrHdNTQtHjexQjLyJwqRP23W8Fgfj3jzUFCjZU4KSDPQUIGsh4
ktCDW5IIAEcqf3SJxC/Gpw4CqR+bU2ZjV82v4d/bjvHyOpGDLQxDGoMDJZU1UOr4
wDarNFfXwBTLdVDQvRUlgsUzEp/th2u5cvjv24tlAiw5dko4hZZ6kQsY2z15CsIv
kqUrNu3AKM8Lb2bZNu1AHcuLvGf9sndP/Y7bES/+sALfYlcQ1qLydO69WBcmmtnk
smdTuSfFUcKXCQYx6vskiekiMaSb+GRy5up0q6GPXz5ac3Suci8803gPnM8kruAg
yCATD5EQS+ZycyVe1rlhjooLIARp56qLq+IhzJ/Us+RReDC+zyeqIIVnJxXhxE+U
T1MeUhJeIJdqwDoO7K/RQupk0qnM/KbU3v5sbdKxnCR/ibzWgOF7YJP8UesBFh2h
5ROsgE1MEN14cbq2iU33jYr/PeV8QhCDnFvdBUTCaUFde7hwaB9s8I6frDr15z4g
ha+HZPVNkqF1aKtNHHwJUi3zZb62PTph+7dm2D6wnTRWwubw+OsGfmErbwmpXfP6
NF9L3I0tkDNOvO73tsHg1d/sFXA39gZ6m87WOpvmQWi2IJCT4+B5pRRhtsexiUYX
9JAcIK3zeLTCR1NAVUXYEDUK6aFdT8g/zNn1NTAESuJf/YuNzQza2M5PTaJzk66f
5oFSMtuqmRlDwITId1mioMdbb8XOtUQXPDnDm7KB/lpFAacnO8Q71KkC6s6qvJ8K
TqMYE9e/TIp85QwnHcIxEmaTSXs1A4R2fn3MF1kSUp4GMFcooVARazqiFK6p2oaE
fPVGM9o3zMWyZjMWTMY+52Lqf7qAhOQUubLTtVQfUfs2IjLqRMl7G+ro7JOTVQFR
jgBd8Joe6DmDUt2rJi5vycQXI0v7Psrp3LayyWqxDuR09Po+iprvSXPVOWCOWSyd
5w/XXxQ/n0rhQWiK6RjOfR0GC33wGKQ+kj6dww2k7v1tAHYh47WEaQ4BChzmGXvl
4RXW9+6ft8EeFtoIvRNzolSvThcnKxPxO4+1t48U+oB8gyLkzMJXLHnJek4t97xZ
CnwKlR7bc0+gQT2A3c4egheahzYGObh/RwsB1b81UOMpCai4CW24gH4pHi4qV1Dr
y9RdA6/PwDHQOaKRpkqt+ba4ETgxdtMLj75y5g39AymwML6DwwA8hmUWdhfqr+Qo
FmkvlJtNyZ+xmFVjUX5TaYRTWr9eiEAva9zOhLg7OQjAdWyvs6paGstm2A/w63DM
nNb23oxTe+kZ72m7faAxOH2rLDUBhydtUKcCeHzcOT0xtxOzeqvpqcccOf9JsAZ4
uXpF41Ld65W/CzAxbVY7ck+KuB7CtnMX6Dg0/BExwwDBOaZijF0uhke1aFhig9ex
sr8kkFOdczhIvj311g/ZUVn491EUo/FzyaSASNHemfDLm6lu1tEXPxl5tot3gLGU
Niy/gfLqkCdebN9Udqr8s2O0Z9/YaLiMPmTG+INnFbl1xmgKS70z6fy74M0em8mk
5rVsKJakZ97T6mYFW7CbDuzURmHuFfY+eYTJpz5fPsdoLmmeZeNR+RZkvS0IGQoF
O+aNv6rCLv+GhvQ6ibcwmMRexhNVDU3EMB+PvAB5W0p0b3b39JdXZ/xQtnXESicg
sPG9z0leu+cGlHJoCkYcSGEHnwyMC1mLpiJ1Jn47zgSt1VXmao4beBzddHDZDTFa
X75oPTAAG6+fFZugTnqC7fU78I4ugGUYizpWcBPnl6vunlYioH9MtotiNL3HGuND
/x4PXEcITwDE2A+xst1cS07pyGbh3OLtbv1hvp/Gzj+r6UEaRfjE+vbKgk1b14UB
+BeDSA6pSv7lrwtcB5fvEjh6iCeHxYrTQWMBx2oTRG/A4Q1Ct+wB9IiFSlOnwtj5
/loo8SsQDuw2x9lEfUqamTr7hIHS1wZSca3ATd9FZT3J9tsk1giPkvk/40VHnqJE
QNxKDjVr2KvsSSlk4PLYWXkhvoiJdRy+GSWtmp3BywG+X2SCCtCsG+mDpO0RlpnW
zu6tKQ/hqUy7WU4vvu+eXmV27quo2d/KM3L6J8zKMYayYHFHN//lTGWWCVYMF7EQ
cjHA6zxOWfs+PropvrvmmpQTrk6+Pb3zu+4byr2IlwY3e9xrbUwwTt76C+tsor4w
F3/Je2WlJ9WJh11Dg37NSr3/QoYM2UsBLoe+r92x6OjSSCC47ajG9ve5/NY/f64l
UN+OuA+IWYx82y2WA9oNuUSdG/uGXo4ht/UQPLI4pkbmKXECOsmOCh22i4C2Nene
MXj3vKZS7r7BBlIt41mgyVPBRPX/VM6msiZPGOmtjYTKJ+LmYssO4XJXHt3oiJX9
llY5CsFP1fUDw2hYNN/aDZ+RBUSH8ojrvj3BYSVgE52pqAWxHx3N0z1IEqZGnrFW
JdBr+T77ujNpEybbQaFA3EuftuD0W0AuKPU1BU8zaB8GieBrF1uQD+BkysqEieRg
lCXHGY3yQji0iIhH0hibCIa00NiCTv/idjVqbPoxDQtLT8ZSs31YHfg19ImC5WFU
E4FJH3gag/eRDnkk+34W9dahTVsBE7RuSryawvqkX2EznCbFfTzTd8xxlEZi1U8K
Hf29hySyWpcvuQKbrn9eMa0WFdyS/xw3BN8hUKa6bqSz/1SJ/SoWb+Q/ICdNMJb9
Ynyt51pRJ3//nOUZjuBw1ECpl10Yu28mcnkZyY/bXnevrQ8C5qkWrIh638G7Z0GN
HXsRCYQF7qHw40A7nObtVAZTJiXSIv+BTz+qy+IaMVmucwb2BMOXBENC/Yt2MVFs
RqUJ3Mcslxzym794F7cPAGdpzKXQB1+jFgiVqinOMGsehHWGKDYukX0Sx1hLer3Z
KTLNZJ7cah76LMXBntI+I0UGcb27wKETqH9qxoNMwFrMXvEjVmnGHG/qp94fmqU2
1yqz9YlCk8NIxT9wLP6EQA9YT+hhhNtjgFcZyyH2SMdcJNVBc1k2UrUxHcxCEyS7
CzYekuRap/sZ7tHrgqO/6xsazQGMkB9CoW42Xa+uVBN+TzkqdJ75NWARN7u3Gtp2
q6bBfWYfp5OkE3XASnf8gBLL3m2hITLPKabo/CpVzwpPTgTy7phrTQya5+iVaqcT
k2l845o4QfIQW/kLl6jGlH0Af2ueU1uZEnsR0IpYKO68kF1eXIHpYuLHVX16EfAP
AEjN4HAtXdADyOWM8AACVQUm8USqzW2H03Q3GolARLMIlTuHkzeissFPHED5TmuB
CSntu61XWHsPBikpLd9vkXVCla01qedwFRYLgGm5imYZaEbBW23nEdZ3LDkY8/qU
/8Ms0x/lcjNMns/Z+s1kHCf0c/rhCXPuKPZ+YDEXNZSqQshRZlXyqsHYX04E0Ksz
iinKxqrvu0xquuR0ctSYeI1nPhyIumqrc3/y0Gn/TrV15+6ZjRKjqbZFPDefh0h6
KxDzx0nWeSm5LZRO5vXjLhkZGp5YiraBtm9UOeFUBZlWELdbaeroS3XxMFjklm2K
dF5+FkoTPiMuNPcKcOIuCuBOWJVcX7zzO8vD7ljrNHrHuDXkBKboc1GVkKQ3jng6
AhKmGtzQTvJEpk3VdW9nR52XIHbvqoixMk7KfbcU6ZINtElz3Ljl7CXvEnI6xAuX
wFWT1X64GI+wd6Mk0/mXjscw4Dn5LWqzEvIGYUoDm/xqmrDzIu6l3PuRcshHaslX
H4/knN0q069HBzZ8mCfv9iyFHFou8h7jG+Nx+PxOF5WLebNVJCyWNV1Wg9EDcYIQ
FOG+qKq9BJ+xHsXuBL/k73s0T9UZvAOFz0SsHJ/8flpkq1hY12CibC+9GwhUqvki
GvwtmqLT1H1xoQHXAViWCArODc5TusCsN4SeNszvUchoov1ZhNCxU8IIBRrhRMGR
2Up2vIhQpXfCv2KiBZYUHxhlgiAwPscGJKzNWu8juSRizVeA1CjuIY6v9qd00E0w
QpnClxP6fX4lyufzd6nY2SLVuCbVHT9Lo6SdaqXXUQa9z/t3JJ/Axp8e5Lv0hfR9
xFJQOYz5isrVvoYmb0J6uQqJD4fc2Coy5rHun81nkFRXgtvoJN+rcu3MHfudVTIq
zC8LnnBiBDQ1FY9srFLTeoa4RyrcWAiOgFnvyvZto4NtX3n7UWtB2UEY/4B1u+hd
/+Hzjz3F5wRRzL1pc6i+RbmHH2DdWUym7GVYJL0YWxEncTW+7p/I+eWMJC8ZJiQz
HgO6lqWv2+Z4Ox9hjK8p/qaVecpUs0mpIh5xylPcA09irO0kwZgvOKKLKRdmABzT
kbjr0yfoQ7NDSNTrV1Uj6cZOzCBl2AH06M6gCSkCUrfsoGgrcRkiwHZStEJVsZNl
32r8nwKXPOSUHcH5YkCN1MNNZobbZkNZF5TbiFmx1QCVkU5Ei7rs9rJlEbp3lcOK
ggnJTH9Dv/TJufXyoA0nrB6YQJuYiy4YZGApp2uNGDe5vvpwljuFbuWWu7kPn3s7
MponIHfGIYz1Rw18T/cEYaW1XphhTxZgYNkp9CgykhhDgyoqf2uHzP6811nyOPSE
kiOumIKIJzDwt1dSCGx3N0aOU0iWdR4F4Rb5L4O2IUNtvWwrTWbpPBA6UaRxy3lh
4AkY6144gLp0x49FLuwX1/i1jsifQCEb4+vglp0OPPWzATe8T4KkfhUZzMwKjC8x
vtXvuRWtRb+twnRZ05nCNpQCbYYSvB1JxSF64OE+d+TimvJCOAWIpN+mvxmXR1Mz
r5BZBeG2DzMEiD4+/82L+AYUXDuYMCmnYp13iKdL0GNNMFBYQB0X5SUCMkGk1zK1
HpKOJ22hgvLypLOPSi2UcFV316TLGvir9Cov1I74+4ofeUSZ9n9RHOt81id/ZLzY
OR/QsND6KyBUhLho7GJ5qRVSGhlaoyfIFWulZOjlqv9Z9muIv884VG50OybRhGtL
ZfWlw9Po4C2E3Hc+SJK9zMzKOWJFWowJUFNOOUOXavRXpm0/pC+1UkXay98c9awI
mK86969/MvapRzfoXiU6ztcZGgDge/MvQheMBUlRVdrYZmlz1x78uHP9n1UoquAq
Wv64KraCROGireAFP2aiJU51Z0fzE74afUNNYiW+8d0faQOKkuo6sRUDRgEnBvoR
TOVxHbo6a9CzOBFWnqfcaXRAakrQ77lg8bFWqDVJ5I4TFjp0UhBlL4ApQmeBZPu/
2EnjAqxOPqI9Rj9DXGJF3IZ9nY5ZJPTPzN6EumpJdXeqXqSxAAyWuey7+JDQGo8Y
BTxhBrIn+vXzpjWWbwzR2KbQLsfxjudo+jRY7iFjEIf4J59A6b0vXwIX60IrjvUP
p//NfC/DS7KAzAYNAHUo53pw+xn9QQnc3gH2TYAdC2K5pMq9gp5zzVF5QlrtM+ZR
jUcUQGSugNmdBvALUC6sT1frYlyZAw0+otHHjxjWbLel0FdUEk/qo+93r7FW7j4w
9W9geqJd62muSHooza3WdAAy2BOlA1awfV6zLO+sAbjesMmLQYUoWlIc37Jeb3gp
UB+MX28aZ4RmK6RLEeZPbYSS9H4sPLHPN5SEp4bK2BUWCVWH62UBhGPYkLF0yl7T
FPqisY98UYIy4uw6kdqwUqCRBjlu9oXRLQrhgf/yGvl8xUfIERzebzFvcDmbqSNd
aQDbVI4C5AH83tedIMlSkOId4pdmpPPwQJ242LDmzt9tUpSNeGpncoDMjPuT6R9T
ptjxC6Dmi07J84RstZz4pfA2/bxoLg2PintaBXzUzb55uywR+KXZ/YrEN3nJ4MFY
JRFrfg2poUN2HDTrIapKbA6oDXQsvZMKJihNVcxo8tWXqNXoan1evJw7SH8DEOmR
PpeZaWSnHEaUYUvW4qO5+Bgu957SbmfhRtMeBOLdKBg3/D756LgIZxd8CEgVqE32
kRJOXW/iMe4AzXDVOZllb24OMKsUmsqj/5kjpq0DJJpwXIZJ/lkajlOkB47QL4Vw
3tGxwG/keUl24IxxEIXKIyMV1DcueTsqJ+sGbGzJLMhJHv0IPxXBztKS/X/1yDuc
50VUhdG9EnVWkJPIV2Ken9sIlZkcnXMxCH2myr25vyPeQzybX4qMlbCcYdB6aD2L
fFL6J/c235HO0r85PO4sFo3FzhW0T6AilLSeSwhnDVwyHQww3eFRZHA9IFDL5a+L
AEZjc6h3GIK5e6ASPGC45dQmJQp8eFLBqNraWxtr8R0V7i9HlgVY/OoR0jd3LSSy
9xUYRL8P6x65lZ5gvBs7VIX94YgEgW+asAOf/91XFRAkoBiuO1eOHkuejsxlzK/H
diF7IiqHMRVZ89ZqpxIkJcQvSuVVeJYlsf5hb6dh4P9LMkDFGXxUM118tJQGijfn
1UrbB6Jze51eJmRfuiBKOyhOih4g7cujrAxZc3JN9E6P1hfznpDEBT8UEFe2jj5N
nWR1gKGssCGtKQXtHCjllUR8O2KJQcEHniM2nJ2/Gie4cBOpsyWrGwvHM3zOgoBG
voR75LTcJ8SpoFxILR3xSRU6W78RJz05Fl5X4Zkhq9cJu774PokoiRlIXL4PfvxP
10LdDBe3mHqyx9qp7bSY2lRGDbnTKdQS2QlCzBMzrszlQqrO2AbgP03NzGFR6Zfo
o9djXyYly3WlPamdeUyj+jRgxfsRhbwASNTAebAxDpbL1kyz6GYjeY2cAJvLIHjY
KJxahJfkEKGxE7eECAyF3/QvouA1dGqs7lkUIhUH5pPNIr2UZm873kxNk/kZUZlx
9Ddc63TRYRNPDm7nsJ7vG1Dvr5Vi6xafxY8OOL2oMVgVnhORoj6Ys6caDXP75ci5
8z8V+nLueRMiBRbe52OtcGKvcsdnsbXw3Bir0Jt6KOTOzv+IKBbiW9csj1dYlFC9
kOcgNmebkfDn6fCgtgo231OxWDGTg3gt2z8mLFpXfHWPOUIgKPjgaB7B8SJ1Daaw
KMWl8WeXXTHZUHbWTCMlog==
`protect end_protected