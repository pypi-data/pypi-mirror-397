`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
tmR8SrUqlxuDWoa/WotRNFPDa0Fh7ixcpFWPDlyF87WJPrWX83/0M5NCQ1FeuBvJ
2XjybhJLhN9hIIq7bk8OJxbrON0DL7BkD3U/bNfUesuXs6OMt7/AvJPLi4xNBBKd
ofiCP3wNiRFofb4o4E1emk/6JexWbFh5kyYr3MrJyGQoJhO1Ak1kqeu3uPWNBUWR
Enj6ENXf8QA/NVo8yWiQNQhXoOoYUdvuHb9W2nmDBGMhk65X8OsAGjLyJuZ7I4h3
wR5s2Fumk44o1Ad/OFtwP5Dfx/zU88LX3JKhQnXDPwrewBdFj0KBvAQ6WP0Bl5BJ
7Q4k/ncgTWGNvGiHYYkfWZeqt7ZOSsIEIhhyLkojIp46pIb049Mob+69wnoPon0m
38lh0BG/DnY7filsMDnCYecdQg3WeXREY5NRPujpFpWZuakGBvAYOs6qPE+oTJLB
jAp9GUy/7rRaF/18hiM54fKbXVlbbg2MVdZLtgTFNtncmIDxvDC/aUXm4cfyWJLU
eP2Nx5A+uhTBrJCcU+O5cdqOe6qI2s+bneiQ+8bzkjSMQg4qKygaFxl1ZjoEvysZ
WnZWfJSN0gmiUx6IQdGMEkWEpJxzN1t/B6Wr5yP8JZLsdxMBeZ3JUXMn6LG9gMbz
G2yj1DvOZz4vCIKvZ3Zp/PkwhXulVnCx+slt+JbwEhA24aQ0woeo+84diG1447K5
j9/wmh6c7sHDJrjKO2FLpmUI14L5hxuhZnLOVmzPST/cMxH6QVGDuhJOYtPoPngs
cHElJTapiFLamjEk2xmgNZxAwKbKbzIWTG5Eg7ugTgLFNDkYjQbDG9jO4te3P8pk
7VuKS0BEYakZgryYA2TFB+6YE2d14CAp0hVYwcZiKEW+7JfCrFNMXJ2PMA9uIZii
QiZvgf/dgGjN3EVSCqrOhN6yGMuWOx9aKBu1Im5BaKvmNglzMKDpOjrAgsDZ9kth
5Z+lpdyWCJKKDa4b6NQf/n3ksz3YnzO5nv058r6LbLaZ6VaI+T4cVsKCHjA/j5+2
C/V26Msico6Vg00kUnccsbKTFcSB1Rm+1TUmOw+b1oO80T60zp2195gEeSbQnxKv
OueXYPdTN7gZiXHWP1MzgMhUKo24BQ8sml6MncfQOmglqpzzR56jkoB73J5wXFxS
AhHhnbI/FWT+bYX+28ZiwqLHr0VENL3gv9S+2Iqzctd114mHOVvOMGAB5eXSeWuC
H6QiYtW55Lpe7S5enzbTI0w2IXMMZTBUa9FKWUZeTzckXP4i0kW6pjLZVB0z+kCU
b2EH3IvDSP/EpZpRfAGVZl5AFkqJotkN9ZJ1+ANu37D9+8uZ5YuBp+t99ihUCmMh
m0dgrZ8b8DrXldVn2BvTt0TUOUAIbBV5RjOYqQHcUCjx28idiY0VLGAAHhK819So
eBZDptW1j+TqBFrniwf22RW1pADEPFyXg2xH0wv12X+sDP5iZpki7Nh+laUa+4kq
NnIrvsTDMEjjiYOLv1w0OEfWWlygOdqbT+Ghn6W69SHuspqKawdsZhZwjFB4OaIj
/cHnSc9OfYN+MrTgVWLkAarFg6lG0FE5/u+yEji0EYmPgZ7rRtg1SifrRXuhfoXU
3ujpBAA08OYqFBAit5Rd4lQwjtdSXnD8SRt7TZRStQewfJmV2qRwCJ6mALZgsYA1
TYNCla56wcSDLCraOKdLgzLR4B2BjqNAizLZE3v+Xc1TrtABJq+9z3WSWMw2LTqX
IT9NUWK+LohS8gbC8ey4xY5YDWc4PaGFOM7RIAmqen2z8UqzXSXB6GVBjY8304No
dNMiDlOKeN/+XmD7WdzgLqWRFlzIO9MS4W2P4m4+/Rhue5emXDDf7KPBJRi03cg3
qMbEhTJkNyI/bazOV678noUuqM8okGCFjnkSbJbQ2h1iY9KtJSoGqgXKSXG964/A
l0+SlnlI9gtt0NKWy5nQ6Bk5LXJMxqENjiFUR7Yn9fy73rKTj7GVeaFoznbKMTLK
q96arzXb3jb6A/gEC9rfe5uxHdo2mFg/DpBTA81gkUAa4H+iMIuSizGEAG0FMycC
xrnqIy0qEIKJnhr9nUYJY45/JWJJfQEBxPJKc3zkFizEjh7GpswnP0ix/0Z9h1pl
+uDZgUVRYuppnCOBz40rCpLo4QaWpbV5aNJ1HqFSoHBJX4J4HsBWsf6ngek8YBhD
v5cv2t5V2serjfcVv7BKbAcqNMZVC2rJNIS6jNjY1Z3VODJyy+Te45NEtDLsml/m
xXjAZ8uUkgFPkzhLIdcQR1SgANqU3QiT6Fhq40baxw8ZYnqD4CCEuw776sUIggXU
zhZ/ckE9R+YDuqMOq1wai/Zs+AWRIxXIlUvI/vQQ/sViJFkrmQRgzochGTCJ3uwj
FMrZlLMc3v2Ikv1sMQsCHSbbtFMMgVb3MqaVCuVSsKWdgS9hhEYpeAmGyFRB26jg
qnJ5ptZiJZ11OX0Pmb7hdfUnkxuMmV1UDgkTNw/mNQF2FKeZ4WEAau8v5RSOPDXK
T9qmPC4iQvbSN64kC62mE3cGSZcddqXe9+0AmD3I52v5Og+I43x3X1XfYGkAwuwl
q/00zghI1Fg4sx1WNxMuAzbABdQgwoBtkWnauLwRV2Jt7Q1fTnsm7mlgZtnkO8gf
sYIhXLl1KBji2Wp1TpEUMc+sqqzO/yzEbghMLO++dvYFZ8gxGQA1z/xAx3K4N2ve
OIheUkIta6Wn+MlD+mqw4MpxVAtTBqvbeOnxznBVh3l+1CMf+70H2iUN45JAjaKM
wWYW4P6KhxIVgm4PEVtSJx8U6y39uu6pJPX9bRVCmSbRkzlndhyGR1uqhTrrLzHO
yXZBeWnT3h0xWL2PIe8X6NZJSAL+QhTusLZknQWGX2ksadLYAqCZP3WKOyerXYWu
3c/nC5ya8l//pVL8Eip5l1m6qWfrWCUs1QhtKUyQSzM9MOKl+THDuTiRk3ueQJvT
3E+jvuEpas4yfTaOXS7gCQivjxWJ+P/oDrAKz/re+HqeDROkkBRgBGhYdgR792HJ
99ZwpMlUuqtGii2sdUOEjxepg27A9Qskq7TVkgVDR8P+Q+rBCcbuGn+DzXngYZWD
WdCRnVvMMNA2kDiFHp0bbZId+XClDjINAnSuLyQbJI5cjf9zqOMamcL8sylN5Kz3
1RmrpPfu1mZdujpN3nTi7ohtYFxTYmaaH84HRL66/z1Fp85l0VQS8slwmWm7tOVv
u9aqqd0bhlbTk6PZI3xcDUmbSyoDYS0Aph/hGOFuaE/jjod0FfPkxsE4JheiuGu8
fWHs6rJJGa85cDhit1FwVcdYb0/2BSlqm5Rrop8HVcxSMDTg5HvVBcXy7pbmdt1P
479LmJdt6LYATO3z8ml/XoVCv8WvB7VHF5fFn6fl154BLT8FAjdKkG+H5cKqpI3x
iijy7D4HxGGfgjK7Fl/tkssAXhsCUwRl0+k8l7Xx0OZs5G7PziDtamWmt0jR8C7W
/kJjbXhls4rrqgwlDCYcz8YqhMvzIsbEt/K4TMMJL9KfDx137yGi2fDgAW/o6y9p
l6Jj45JtTKixR0jUc/babbXa9Rmf4b8QlnTapczx1kifgBN/ZX8FwNDI+LKySdCI
2LJ2jjpohpxKLrBcLdbYZsf8sQkoGmQrHb/ly+ca1Dkiv9tgZkxSxBpSsNSWpRGw
F4TwDY0V7sPQ2hbzToNqEUF+J93R832uDhi7xyQ2pCTaQUF9pYONQ4IYQP2t24/8
DE1kLkOI5Uo3PrslMIwSbGktrmc55PwElqrrEJ43rTYRDBVCUfyxfsZ6Pb91kLG5
DNY28o43gtJHt/8+fXO4GnUY/vKWXdYNkYwJ17zU6GmWMQKMQ/5Vb1PHUywC36Oc
xR5+EtZK67ckx1j12f6Xj573pm+60wr8ETM+iOvKJImLngwPQ28bkaDyl3ILoaZ7
DjfOj+HsuYoyGPICY64Bv+D/K3AjThWW/2J2I7w/0BDCgjq42grptBxZPE1i+EEz
a5EM6HDmck3HIzNwmo7WUWYaP759zFd7BJHDRHK3VQMkuUZr2R0x9bvn5z7Ok4Uf
uFdClxcBK/VQ63wDcS8BJxxi3w1pWcw7vJxJ/OX4JP2wtDfm7WiX49DMhEWSJw6z
Dsd+Zw01sfzGLeHeZUWb1h7kr2B31UFwDK0vaM79hHJHp4/T7f975eRBABZ67eR0
j4zIhSYfHeDk6o70Va4n+/G40RLWwhkImiXOe8qssRpt/AKVXABnb7J7a8mwpLCe
VvEr1qXLZKJCIReD5zy57GfnCV40pl6JwopNfz0YuK5VyVRG7S8weLQWjdUsS1F8
MWM9/9/CZb9eerE+yvB48Hziw46QeJ2aYE75NDTokYmtfSD2t/WOtmVC6SEZsUOa
kAusTiEeCakB2GkVPJzAXXZi+6tdl9tsvHSnr7AC5+nNLbjV/KrzulzXPxDgChzM
lcl7BFVMaEyCjUH2gPtnBGoKA8YcJdVJ4Lkyn1SC0cR2xGZuT1KhSN4S9HQm2b4q
sgaSWZPcGW3kjxRh2x14rczV9WUoQdCNjFIFWdnZbNxRaFZjIK5YNsSWEXEIjZ7L
Pu0w8WlHtUD1F2UPRFn05ET7riCP4lvGRcGpJzrKzNluffAMKhXu24V+fALkweCR
N7OQSqHPElKAGmYuKABQrcsVrgnXoS+4C3+KSOkIHVNSzEv0Vn6C3faopu6d0EyF
iIQnVDvpdXpVn5hUuNeOmzfez7kvpZpAerM7z3/4q9nntlPnuEmDlFVDWccxm7Rk
DXRA6FBK2Rja1AqjTsKUEJdziI8fs//XJGeqG/xbtOiiY6JsczP9lMDBins6uCd3
4O4zC/1j3++lg6rCTiCCeZlasn72oXdiQfUG2xeNuk4HWo2pJRDYmiD4fnwiTkDI
AVNrYQQOjWLyyDBFDshBD0QtgG9njj9ulZnuL24Ec3ZVVFNjl6ztFYU6QDGx+7+R
tGGfNq7D3ojtzoTB9h9TnzIsQEvyKgkOz3wnL0g40q0n6DW93N7UnJGF+qN9OBxK
rhnIzkv4nXeJgD/4UbrKbloteAZSLPvalVlSRu7p2QxOHLyp0yq8NvkFVEziSGRp
28bc7hx/CzJHWVfmFfaD9JdUc5Q+Zc8qf0dAG8brfjsKeGIgyvNHjkvhFIDIPAEt
T5KBiJzfn1vD8X8RpkpdzqsG2mLIjF7+P8pY1VXx0aK59mIriPTgZ9gYsmh1XYHb
gxt/8XNIVCcPEyh72UKDr76t58Z6Z6kJAf18jexoSlnBSZBSfDUwdovfaT8tkroq
NqpNJEz2VdIN4H8cl96ckzy8Lb7aYXUkoJATRtmQRwb6C1eUbJVYgqrEA60bkOIS
DqnWy2T2l90K89KMDi3psGiSDp1RuS04gg27GNLQZrjeisW7XjL5ijrldBM7vRbT
`protect end_protected