`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQCG67q1aRaKD5brUrzbLqYGpSDl/s4luQ5FdSbrQgdTN
qjowphLCmcv8EkG5rYvaAZsTlSCTo7dGYwbs/hnIT56VwEo7fRWfZZAHXrShwJaQ
k/2xy7zfHMprupm3yD0M6cxW607a5NUHK128dM3MNd9aDb6duuMDz1Z+817goCLU
vX5/sZqJSBiE9uHyHw3kjM8ZbNnfE68tf+9DR7STKhKGDW4hZNo4gH314Spd7Y60
C5Zs7XrMxs/eyuj1L5kNFdRcplvdi1ffZZeUsG7CWwE/KJOyFe/h6Gc9HQPnhV7f
uHua7ECqIWJ9MjElAdyjlXJv0flnrlF5P2gQDDsDg7iY9P1fv1dRtZhvFWF6nCUS
GprYiM5ZmKKOby9ZWg46ElW0Z07IKJq/yxDKzNVr3mvHAOX5P655wU7RSKaCPQD0
NnH8K/O/XWdZAnWOosncqpRSqNYn86BoaYcquzDZKIbON7E2cvXW6t6AQmsEPhMI
R4dX8oETxyZxc1vMMfYi0lLeoJY7SiAJTE5ybQ8j92af8ikkYLOzsuI39OyqxNwz
xBVaIk/+0sc5/qTh5CDmIRIUZYBf7PFbuzjSmipgpbUg9mYUZj1vuxGVfRTRU2jJ
EUOIPBwfkrxBr11B4VRlPFHzgtC1qwGnYO3EOSCkQnbn4c3rYaEvH6Hlxdta1Nau
xDm8ZAp2wVlKIMwv6NHtsJHJZCgywQ9nf4B8E2CYk2PSOy78t8mtz9AR/53mRUyy
wHsbdUTzDcw27/3fJmV1Pp72XDcMsbzBQqJ8tbjSfznTWqPFn3LoaURVkzPBNvOe
JLQj9X6PCOU0wS4xsUfgYyYrwL71sgzfI4F1tPBODLkQYexb/DvjtKJhMqgWKXYX
XhCkbuqPl67eL8AxdqTBR4uW3+42+b0tgS/gIbpfpCVfM3oL7JoJOZi6gtYXr9xA
K+Y7fUeyQycRF1sBAy/IbEM+qihAzPsTY7cNV+dr9BnMKmCzrAOEKe+lyTEP/zDC
5l0fgRwiBd8QTyKKLNe59UkPkfu9wYDdBs/u5QkNtrsCdLF1uXTOANOMAQYamveV
hsSf1KInjm3/I3xiHlSv9Q/SbA0M7zAjtCyjT9FEiDSqJ+eb7yKqaVFDqBNZXolG
36JQ9gARqkDzs3Yiux4Z76eFzFvqI0F3YDx7VfQsI3GduVDyYXTse6vvyJyL2IPN
F0s8hjZy+e/UE5QfNcG7KwW3RRHewEjBJ57op7RwJbEzbh8o1APclwvkmhb0q3Ef
yQmkcwUTOzJDnoMQKKlGWtdocNgaiIwv3an1IYPfxEA5L3YE//kUUeBk25x3v/4E
aX4VyUHw14qrzdQTEDUSsaKWhh5XxLFCKqHmaq0MPy6Zq0dVuHAAN8VjcrzYOZGF
UdaY7EUDz5/y3zLdBp5XHtIc3zov0IeLtHrnopuS/SLuk0w7wlE8XMv/9/5K1h3c
UnzoFvOhWVYi6Ol9ktNe7bWNdVWmvZ5hNN2VzCS4dUnwKGwUiYP52QY6Axm/EYOt
w8b4DaJ+GNJaJndMceW2YmjIc1buDDtX6iQy5MV8KqFfitygOL2xiPJ/HIlnkvq2
FUhGbV3Guqxn6IySv3tnm0gIfiLB9ANguneGp9taKNYhRlATzNxCmNz5Y2Ju6T26
e3stW7mzYS6E2NIdT3bh5f7UfGmEWmq8pc8Q2WBKZ8EvgnxKSabGNw2Uqk5Dfr0R
CvCvVmst2QCB51et+BpJYhePm3Ls5OvmVCjIaoVEd4Cxl86lpJjgs1KsxS+bta1h
5DUhv6Vu4X9PrVFvEcLBsRpNr0igRGAMqJnoduQlehEy504TjNuvgQ403fHoHQZm
TaQyq+BgSFtwVHhA2IUDbUoQKsTddzAuQ0JGsTHg6GSrDN3e2Tb3NiMb7iDPS0H8
vgBPor0y//Pp2f9UEQ4IGaQXN8Z47LX1WBRADkSLse+EIAQjERrnsKOTz8gMbLFV
CT1Z5so2XU4/8L58XaDdNO+jy8Om5ElhZePplwHu+LYgjHgSduGmbaNg8HVTbbZm
IxLPOeyXZnLQ78+Q2/0tDhxbIziZA3JVFpk2gjDMt/eKlF7Q8I+aCDOyCRJxZmRc
f5Dx1hjO8JDklNVN4JljBohERmIt9GZJaANWl4t0q3TVocdI416W0339erSmiQWg
NdkjeTZe+rojqZo864fp152Q8CmZrTHFgq0HPZtzg0oeD2zGmRtdqpUt5PvjRz+9
NB3MOdSsXPuK4ibQJ5/V6g9YEfbxiBddOLGwNvyKpHGN+0IjlLoG1OxYNWgoUTbu
/xNvziEIxiJnk1q+q+cDW8jaCvKhHlG6CKJHLgLqMwTMDfaZDBzrmlIVyTPXAYvS
qKRbFHqiMZ0eEJRtAlqIyibwalBbsZNvAUh9H4M3bJchNpShzI6+nDSQC9UWyO6U
lslKYRYTey+h2eV/WxqlIAzmjx4d2sUCkrkHhNBgHcO9h5wOhrLk58adijlI25Lx
P+MdcV7u0xzID0V3f2ub4IkZlQNt78H7HvFI3O/B7OMcwVEdUWYmhX62YGNhLOkZ
9wTkHX623yTX0eHAS/866N/tpKg0GLKYcuGuKG3/z2ENdLB0s3F0YjxNPogo4CzS
RGWHQ857HOqwDJW1RG7zhfMOLV6XGc5sKa9J3Nw0gShH/9NzNYfo7nVojZ/p4MdS
YWdkmbPuRsZzOfyto7oQIrumZT8p4tNi6gCiLOpb+Etj/1DhnOvYyit7AcgtNKDi
2L8P3qgA5DJ7usEVGWcEUx4AARuEQ2CjEiPz8fTe1RL/p6xxCFT3mCOUVlTS0cfk
pbQPnnpLsNXvGwj7jWIHwfzAN/kzkYweQPEhU5ucEMxwtDw2O3bXOtJw74770JLs
S+Yuyr+owcywdlMRV56vcUb1lFa2ip82ctV+HF8btzllCJBAvtoze3nUYJrSAtKM
9o0tNKXunZvgtBOmucmvSfScWFy9kE3Qg8MnH38mRJCPrbtlEWeLl6fD9QRaJOsl
gzpzwHK+dmLNbl868RXJOWai9jUW/depsZyJKInieLYFq/q1w76PyWJldYxx+75J
Tb3LgrHE9JZsSAH8fysvwuNZNUC6qmZm+xaiKizzljINh5DrZhpOza3/nIGXAoNF
oZJLoCzLFlnrfLOIiA+dC8AdM7HdK+3yR196+V+uGzX/jr3HpvHl0nfYjXZStl9B
UlM5vBOg6NQ4neUUuBqL4mUzLfSBUmYtIgh9Xi2Q3X9nOm2/5qJOEwhG8sc2FC1J
oBo6qLO4Zdc3RNWjL64zw9bKB4cVmWtistt/xeOsAblFS5SFJ0YrJxB5ZFZrMjmJ
TV9d4JIDT2hbCkV/5NzGqKrZ/9aaFsBEYiCn9J5zqd5KoejCPrrndAATUB+hB6Ec
6KGf97hgdumJWYAKvdNu/4dger7jHOEA01XWRnCJf7i0JsorpOM1musWAVitJrK2
sl+YMkCpNZC037UxUzkfUnpVFkIA17m7Bq5JEaC7uGOQJmG9GONpUsqUq2iK/p4F
rodW0a0x/51HqSWmaqOP+Qe20P2NmPZdb7+ptmIaPEWWt72R0FDtS5JINCJmDh6m
WyQDWGMwnIUqdlfCO24s31DrLPTd/MqQv/bl/+D/JtrcWjKG8H9Bv/n1g6XbOgCY
A4Wd4/vZhysUoKP4Din9qFydtp6K+J8zenGXF/dTalYzHiAX5R7zlulJAvdZT2Ux
muCxO/qsTZ4XsCp3n1X0pFoBJkZPKWdgHkTgdjj+T4Djonpt13PWnnCjXcmhAVPg
7lJkEXMG00JKB+NMd6COSEvGBNEYGQgzntmOslIdFMfYnk3V7fnmMoluMW000amN
4VDFWvMefzs06aoO4wtlXq1IeN/Z522ryFhJuwlu3fBklWMefO0Z66GFZdYMqyRA
orHbwl2schchQTsv+aCdw83gyhbntK9G/7zkuV2B9SahPzwwumosgXhQGXVB7f4E
iPUESviFDjUdQRPNlfCaJu75+VzcRiAd1F0k9q9wCarFYTL/P9QqejjOPnYMLRZk
BGy7aLRb8XiFJR5s8d9l1MhRpEaOPKxzYJAdv8Wz6ICsCYH9+Bk/ADbRk9FxQb4o
YzoM+NqKE02Q+VOxThUVJzOGtG9a8UnewqM+4InORv8FBFXbDKjRovvfF1TInr4g
9y1ZOQaytevKWaNZOjPpgMWx8lrSDs9COIJZ2qGbfvK0vrXwt1dm/cQuorvERArs
hYFVwKsCPqe1oc7vujUEkm24YRZ5PuT4Wr/TYAryg90Bftw0RQiIy97LfSxIhwBf
nrE5PZYNiEjb0WBdj559lE9oautOLsGQDsDjtsDStejHxBuRnQtSXJujRyKUl3bv
cO5obK5Af6DWIsuwcO1MDxLEe6VMs2Q+HwYeR6qbFNMRxpeB0VSSMR2+/6grnRQd
89YEc92EgZs7O6PJBSApk29Kh6Rmbn8wmV5BaDyqjPfeq4eu6KG72WPmlRThQPaj
Ys58u/55Qygp7oiFASUWC5QKE6b+JxRGA/2YTe2kdv51ZK6yUDAIVhUztGicNskq
rA5znOI4Eal1ZiQWV5iE6o5N147XeS8fJBK9Wh//uhrzj0x0IdLq6y0dQpFL0Xxk
poDirrOlMuIlstoZjjnjUZydjcznxGxcAAPvSbh1BJ94nuZk+X6m6aUSvosxT9aj
8ZPVbsOHc65MomD5J4X6XM8qhKY/KKz0ojSma3wM7BhQURzwS5iY1mZvOSdt1N2O
LJ1jFByG66M8zBILmAelKl98AEIhLjuyG8FIWAfh0jOra0jAjaSoZHBZngNzALVb
H0dq4wwGJNzSL3j0lgyAKAVMX72ltW5MmhB1JfoCzxzfmN6BsHHwqaaJxjv2YVnr
sFMXTtalyDi6WG0f2J01P+akhIVY7lkxtKmepckBCqN9atIMXAXvtW20Mzbhb1or
KrivTfOyf/N/dIGGPcsT7q15yg7qX0btwVWM4rKavC/XTeDjY0VgKvbPXzZHMYog
wKngt0QM1rrGUi2gweGWk2M3DTxFm5gTIFquZBgtmjZnJeiiRFspUpBWit6B5Rld
LMy4W94tIIMZGhUPhx85eiG8Zssg8ptcQdJZyELExl0r9CK5G8Sfm2dMv8Q1VArO
cVTQy3opILKYv7AWyx6d6YEdyl+OmZUlytGy7nHGwbTzIq3gvXJtuMNkmNY2Z8Tm
G88YGL2eF1VhOxTQ7jG39mILgmeZGugt/yJPufec/nlPGZYpE+cHPG+hPel7t3kt
bF3rLjZwyDswpvd8LCVXkf0YEfDyDC+e3mPxdMAQlV6mubK37rDEX3iqtVUqqpGq
k7IuvVT1dstG/Qz9iGulORg02xq5k4EbyDI6tmi2jEDezS3D49cn0UIAKwa7AoqR
XKjcc8I9z0FMQQNwBdW4VQnymDwNQIvtpQXrsbKtwBBpbfZXDsYWhnIkRdN9gQaY
pPG3JzCvi5zFu+u1E8GNKt+j0ZXpdY8VlKNLr9X9mcdPMWUmLfe1LiqsKgzReS4Q
XLQ6PzFDPxSlvv2M3WkpY2cYGigue8KMhKMY7spv9dNTKTvWbFcJOoovib9+C8ny
zNBE9LltEu7ldCvx8hGpsMJ/3nVynJEmpKu3Wk1Atm1YXeTYnTUZppurUZjndoWf
5ZdxjCxPJNloLZbIGAAJqeQ9m8iSzS4rrxizS9ItxeFb5XZ3iuWzUG5Tw0CpzNUb
dNEGjBVd36/10G7Ou+d/meDk7AKGLAdcOlbVI7aqEOeWZO4iK19s2odl0tebtzzh
af+6co+O78h9KUUEv4acoJkUNFFR/r2uo6AQSqsJGAC6jLRwNDjT/7wTvdng+2Zj
AN5XnvCeitdIncUIo6dlyPlmcGV6afseNDaOWek7kwk9Z+T29pDKggcfSi7rx7Ov
HrSBxvSn31mS7MsNAmHetuOPewrpy1ANW1CkV2DObH+aemZafVxK0c+sLRdoKKML
7OWrQ5w0JPVG+up/O9C3apXeIFqe15JNxp02w+wNt7lUjb4hFpbVmmPYq9Elitqv
E1jskFNMVPjfvs2QaD826xfGQDmimG5yLBnoJMOE8qroOl7wBCX2eKPz49yRa8Xq
xGa+GczDyK+1lnmqkIJomTPgPECG2tw8pleFip5vy/SQTUJH9+CtubE4RAnl5y/V
1ypZkpiIqtunltB8kY66hu19/WyKn6ZggYI9F4vdgsu38d/W43rEAUwzLF+gfPrg
rzC+Wf7bOfK3lCfFoLcg1vIBV2ckZ7Lok7r+KTRApVBLEh1Q3/CiMuwsodR7QxSz
KHo7q+jRsBEzAfbUcO3QX+tpaZRZ7GE+GF/9zMipZWcnPesK3GckAfZAQSAZ6gv5
YKKdaFqurPe0E4MfFz5o7aFx2jJxUQTeTqexJlmyzq7HmhgjMk8G+g2gOsJh2nYm
tMxTC1FCLcrzu9YUgZXfUeAH/ZFHnd0FI38ahBs8Rl/X41emBcBiCEGTXf5pchE4
tT6YkdKNKTTLkKexGDEY93zu/nWF6tayw8Nny7mi0jukx/VAFKrNak/wrh7uRzHc
EHd2/QYehfjtcESHcEPEHoYWwMNRUfSVYTtdTX/HwbqVm7DC64ekIWx7tEobiUxr
aNELHA448B0UXa6VgVrwkuIm6AKhBjlE67nYWsht9+VCUYbs7Mhw3QbM82wRZWF/
MFcZUAtfmT1B8QaOWHAoCZBgPOIyaDvjeooxcAYnDxaWwErQDoKf3pen2UKaV2Ge
9yBoB+7KDeoJu1b+0i+ErlK0Z02+VIV70A1JXWosyGn7kkeuVW/b8XmRIpHf05qo
OlOIuHZ59SwRrDG4OLPoMgz+Ymxr6LY3+vUUOpz3TEjsj4r5IOR8ebv1+26kaCZI
pdikS1Hv/XWBic54wSwlxN/QAjzov3YSmvuRiog6NTUGvaKqt2kItoV/5C1RjvRz
kWnB+asWyNch3i8sSGkn877MRNWbyepiNB+y5/c8KQIUl5muM4afIb1P0qh/ZF5E
en0oiQAARdRiwbbtEZYrxJYMj8N4JNk10WthbOV2OavCEBkhlyhabbzuW663eucr
lUY5FFJt2KSwoT70Yv4R2LDnRiBOkAsrg3d4ZT7cqGL2NmmmnVsh3aY5Ajc0aVIS
djpCvsKCBzy8F7/dFNV7ju24ck42uJhTqdSf9ALhaCO4LMqAikoFv7ckyXxluCDZ
AbCZ/68JS+IzCnhsoU9eXlKo9XxyeXKoIslOYeLlbKURJs5jYLdYbpJlsXcjhZ87
JksdF77axTLr874Xb4UkIj1te8JFUfGHMeRFemy903g1jGDlfN2Qrd/+BcWKg95+
TLa+P5ZxPlpDPTqEZgqBk2ye9B3fXFdv/3wX1TlX/NFcpcOd6LKCGbUOTqZS9BTT
+xt0KuEOT7Q1I2HYH+4R4GRGpoXjMpLucicoL8gpjGYNC/l+nr04RLdz/m1YQq7V
+6QeoBzbOLWw0iotyOzgen2jr+cy8iLnigM4uxlwH94hltK4kwlaH9ah/QlETQJy
5jmA0tfpmFVCPcYBYOkPdYPrPSfsO99lEYbyzx1NjGSDUDTC5JGt0aAZ7WAQOSoF
nrmg1yOS2SeR0tG5rS6OxQ0MWnNjtlQQIg1Aw2sYK2Cf3LJVaP/rd2OvhyQ667mU
zGzuGGd6oL1gJTiUD0FOl2S+7NC6m/XCoIocgGVOqsYfy9G/zWVc2xqZJnefuQ4j
FteRhGHNkwbKlIRHQVjOuT8f8QP+jBxaqWyFXF4NSJb0Nww0//jLn4F+sYnuAIki
terbMRK+WIISQZYELlsFhH1SFTPtJ6uk8wBasctky50ebwufWX7ckaMutUGyOj4W
1OoBxi3knn0ZFPdOnZ0rVnvUiBc7R6AJZL13HEA3drDpmzmBXHtS4EMoyeGUBnCz
BSsjBMJBHZ0UlHaxRXSOrk1+BdNZe9cM6tlA9lyatdPscrbtzmgAFsH8UYRa6uBE
W0rwPJD4MI5Ac5rqloHevIf61m6BIXqRX0+gyh4VQpVl2WJN6nmj1+y2PaTHybrG
7VSqNItTkhwobSFp8WyUFBBbcND5577aF3PeuRcPKrDBfmlowowVleCx+pVyFZEz
5LWBhY4dZiNJRys5hvQasvsZwpF7lNtMFUN3LhbCLB/mDN6LUr9bpFX/4Rx+QNwP
V48UlKf0H5zYLzHfOINXytr8DnS4fJcDwt1/FBWRRgImo3+1QcoW8t0y1iUigLlg
3O5jD4zU4/b1wq0MjUlu8IW9Dyo1jkQEl3J8zSelaplv1PDqvLq/vp52g7xz9dKY
sFfQvTV1EZ4zxucPkkQtNCSBbbyu+P0zcXPzkJigCpmDqiw5mS9oZU0c5wvndmJc
g2NI7PGlE3qqoxW7bJf4EDsPfW0UT4SqTnIQAwcBNAL1Vkia8Qb5FA70rtAp35dV
dbo5cP3N32vVuwMebV/Rjd0Djx/rV0SFjZP1dJTnuO1uQ77XKmh3pNwt5tJBK/ZO
cNs43V5OkdKvHJvlWZqrQLz5p9sBYJUEvL3Dubo3tfusf06hSKfOnt05Hoh9Xqmr
jzLBsPSfenzg4Zd15BnJxlE5N5JUF1uFTnFvrrMXVawAUrLth4ctjUNjxhPk3glJ
5poCSJ4bOJpTKqxZ4ro8HzUWCOw+Q2Tgkl3NxQPZEVU/yN3fPp7h5mMr9RsNr9B4
KF9N9E6icyJotTz3/uRI47wKjSiVP83UlC9KA1EL3odnHG7V7YTYaU/T3HZxMmYa
fNzfT6whf6DtpTGsroW6Y0d0E2Ytp8J5DI1U4UVqip4sHsY/BoKoWbAx0szk1Td6
tNwSc62QHwcwAMBf/Azx575x29bQ6rn9TV5ymavF7jFEM6vDKKd+tg8bsmqTdFCG
WOkYmlPJjH3OAFQKPfealyYe/FzEbhDWtRmIqMLmd2rLaW283d0d3dKGkORVhoro
MP3xNY4JTJ8eLE/3Q9grvLfOD0adRCz7m+1KtXRYGrW+kNyVDSnF+Uvn7K/eACWi
Tlce47oyN2bCB2nYIl64Z0K7Iy0uVlUMqb+NlzDYZhVjiArYie9qT9mgDVxZwdxh
aNSSbFsZsHK60AOKCRyYCK+cEy+MWk21wf40EGMT5ocb2XCU2QL/aRV3Zp8mmc+A
+nqskuJdKdpJ6dmEtWXQv4DBK/1Tqvs6hHj8VGE8UyvgIGoYchvDznLrux8M2qqt
0DPfmwaSOKPEW7TCe3NYdIPEISZm8l1B6UQ3tenjJZ5gcZJjCd95dhwtnH/WoOPs
XYsTUDGcKH4GZiu2ovf804OCwEakXH5rtfLE7E9NVXMTl5Fb2WC/pROWYJFlyn2w
PwTOgoJqvnJYBTK+fcuig/hYMB18mwSlbk6tlGkuvAbHQMFrUf13k+cmGCYxaQC3
oXQjv1ssIsJwEONshd9/lTNJJ1iu7NDMyKQdD7U/JrV8CT89oX9o3kefvbNtZGHj
tQNJd9uM7sXJ0fEtrFLCXq3YoGFVS0j2AkVaIEX6tPx3oApO2ubhBkIIKo6jeo8c
4rp1zOn7BPxjDG4+t1Qon7DpYmp/vRGgkeuD8iHk9cMhifssiukAdnU1SY8DDfIF
MSTFByKBBlIwkbly3vxU8w5j2DtHpYMbj2DPHsGTDe5g6SROH5hDAvLMchI6k+tq
lEZHYKU0C76MuNEPxG0ANybcJiyNDvDWfhHYk+zFveAu/jIe0tjZv4m97xAU5zYw
h6FD1RAcRQ0s1rsvUqFy0eF3dWq+lU4TmO+B0x7CNxYVW00fGndAxNZE4DmAYsCB
sIk5LRPxa1I3W2E8/aHvlpuaECn1f3jg9ivKHJNs855zmrzTQv/QrsFzomNHrsW2
cPptcccHjtNYQPFFRG3fGo7SvgUNLcDam/RERy7Eg1oG8kDkbqWyf5MO7IZFfcEo
l4ZZQ3grv7A5gBiFr6+4DF9o9LvBy2p6pFEEFFBGTdrtl7D3Ppe6xtTdG6s+d/GF
IjlZTSQVJKYO902W9yAS1hfXqmMAnvhymE9awngSMrAX3sfobXAl+dpGLghicvT6
8K0YEqUUcSr86kVMwnVyLZ/xrUWrlqL4zp5RT1S7Vl4iLdqe/1o94lM1gNX3rpk0
xw6VyzhkhTWVCFu6MZaJWIAt848CzIkUATN0FeseG1uXSyDegSsSNDdit1ewO/lo
YsPHxlzBPlxlW2N073zJ6aWPvNgyQc3KHthM6aMa2iSXuy9aAqTuO98XUzHOklxm
Z/JojprDqZoAEBTh9EudfKlAUaLlLCC3dfqw1/kg+/R1uBf6cPEfRdCa01xNpO0d
vDZs1KBi3qHXKsWAoARYze4lmtS8M/Qrx4X7q383671GAsIoj0Ew682UVXF86xJu
Ws5BSGI4TmLU6aBLTxmYIXNGqy7z9caO+5L25iOH/H9gTFxTsHWFHbeqJ3x2WqrJ
m0lhZUR4oQUBlX7xtp/OEu/4ahluuyNADy4aqCcsuEBWQYwikfdjByJBGfmaD+5K
5/LuYj0TidMJlOIea4UuBI4EjhfUiSDS85YyRt9UUXmuMT3HqMo3LvmyIIM2Se7U
3qivrVqhdyMltL4MVpUPxdgK3RF2hxsZZ76uVDZ2SHpzUPp3n1zSI3Jb4yPhrqZN
YDeOIQI2eGjVP6jbDU6UFHxMbBezBdXjpYu78R6o+WYfbj6KgiVzYS5vNrH/JdLm
yOIc4NvvKydUYnS7gtZ2iZMNuwuHUJ9vqLYr8+eqq+oeqB3/oDeS+XwsBo7YELL1
MrBX4NWK7aWyf9u7o2n6foHiLje+L+SOqC+we0RghCbZRt5Y2W2yXduxR1e2ZSnh
7a5qp6uaARPMu8zphWMRM6csYUc5j9PfJPIiXFDrFa1Pvwulds5YhqU9FlOGNlNq
YDF7G2snWKfMUmLhE26CAfkE9ijh1XKSa5agOLtuaQ2v6nSgwWMI0EBAlmlyAVhV
DtLG+WLW+OLFhcAWj9QSmo64rnHreCsXfuMSSVeO+5Wok8JnseQSt4+Fl/UVeZLU
rmh1Nxx/P50QPye1I6lPQ2Grv2dxfs0gf+9L6QnJ9+oYLC/Zqg4f7Xx4OMslOYtA
0HMLz4x/w6MywyYPkT0Y4Rb8eR6ZLPXTop7iuSMrayyFijKn0/fIBCjeImr6p7M8
5mcWibMusISPPvuqAm16AuDJVJ0R4YxyHyOogfvWuHTpZeuHJc+qO958dG4MOFqC
mHIwAmPg5Pf82WVni4wtJLl4N2l//FPDkv5KMeWlQVTJJj42KU/5KUDtERaXy22x
jxTay1oxr1F3oi6PC+jU8zavVUKNM+9dEa+fEIedtboaYPcCUc47h6Q5p9HnYS2J
mXJZJea5MScNffWSlyQmvwVbq8xHFMO8+gyinJFGItpN7RaB8VOeXmcBAHGBP0xf
HCjvoCGMuu4Di2BlpSacC3KEAcEz9pnq5vD9YhRid/W/9+95vNdU+cp9mamTe8Dm
Un01TA/wxB3nKS3rr3NMp90KLwgFUaUTSgsbExnhm3D5eid5Z28elTh+Imu8uScq
FyvP/ErAGJiI0fov2Br+wfVP4l3uWsFCcK+7zUsUYBTcYcnnwyW+q9dvLA1yVpgL
Cc4UPQASIk1AOqCTiTJgPyHBj4HsYZa5dve3VsCHLmGQgVXubmMOXaj4cUk/GCa/
Utdk+kwilGXBaVrrzNyvoLEHdR7dQe4A3e+gdP8ljIwwee1cKBRJosatKcAjqS2t
chIU20GvntwpvKyKMmj2lsAU51VU1CyAdV2sxJypLX5qJn96lAt3qWdFdCappLsf
CH0MaWyY8xlrGTPd6PrpfbRYgU4KmhF4xPdidrDCNtsqaHKSSankNnc3qD96edLm
hXHxNmrABz0nSDpHjx2qLiYsm+1Y6qmmWw9SZEc/kwBQ+piBquK/EnhW9v1/Vatu
K4UH/nyqZx6l16mptpsTMCSopnCjt4+2aSmTYh8VuacTRGGLYrA1b2I0BECFyQUy
TfICxJbbZ5Kp1qOJdJARfCL4WuD7bee3yYyZ2e/6WtT+Ams70rgjQdSWwQl66epb
qRKzaSUGmOCV3OH+xG/Q6Aq8fMfS+hfs4InlGI7689/pgOQIQwNzHVyZ2CGXKbFC
VPQSLOOBHNRAF9901w/GgKeym59MsuV/ZAOJhfWInOt6BZRjb4X3UpUHCs2R2ixX
mgMmQ03/+F0kh30Gb9aJRAfpM+NIqFGWGtWwo8C7ruLeZj/u8BijAsKdgbhlInNU
l/B4nLJ8Rvml3i3LNGTOWSM0vlmr+GGpeJQULBeRQf2C+c7zxcgJr3Xuqm4BlQvc
D5Krba2Bb4hBoouyBgOYYIuDDzl5SnlT0nEYV0dVAnCeZ8jxZAJXYAdoNnbno8ZT
04b6Zx/f0zHUN1hKuhKcxpGtxDq3G6GfcRm9O4BHWQFSX9mwKU0YSMK77Vv+ZeoX
agkWpMPyta5DlGmPB+RV8w4695twBecpjxgZCvLJTNn35n5SO4PpOJ9mI82CI0YL
mDFrxWIK4OXcJlYZTIQaPmtycUbLePMdI0qEu4FiVHNjgTiwBTZB05vr2W/+4B0w
D3duv7MRMsX375aa4M3oQA+3UmmHnplSPGHAebFcPkKdDYESNVyV259BJj8c/3Ay
TRVkH2QBngYpIk1Mh7rxrxZq0JTXX81dSyEQBZAbwjeHjJTJiYZS8Z1FADpn6c6C
KyBz0tIr6EP5MEWMvlWttMv7xCXtAwwgIyE7liy3yav/EhzNYzJvQpL78aesyxkv
+D2/YZGfP5fWjE1yGUymlHwMY8f+x7F+0WDbAZlI3IMAn0PFWdmaVn2GZngCpMZH
aOAz3a0s3AD1rivO+HI3GC4k2bSoMlkdrgO2yELeO3mGzGlxzzd8E0ZfeX0liSP7
c1bPdthcy1u+yG25FIG4CR4wXkmEE33xZHX1XF053IkZddI5b7G8p+FYkeBZNw1G
m9iN7U7afVS+yv+kb7+7vDVG1Vd6QRE/eOs6gy1XOjXSUW+Y1p9v9dbsyUpTkBV+
dztG9J+B+QU6MjX1W+LrXhAg6ZHxYPC7uOPr0/A2DZrcDa+YAJq/5srow13cKsbD
+gGjEwM7veacTeu7SSdWW/fuEud1b3w85Fy88uydtFuoxugTdsW75hKiWb0K9h8i
N/TB33hVo46k907z8/N62St5TScDplKYx5sJ3uNq8wZ35cH8/C6BVFfK7GbvDAzB
m/w47wzFNjH+UFBJgvCtEowonxMQTFVeDYZudGGvN19nHt0453VSwi6C+56tV0H6
X16N7eMtqSn0cJrAGDlVAT0CB9fw+9NE2VJJigNC9QOX4vhd9zCbG54Ja53howYr
f5862YJxcZ20YUPcpbVdiL31hsWjII1lvJO55HF5PWRDS7D4TnMlyaFe8CKs7cPG
Zumtp78DJL1bQ57o5kgoLhmMs/RKRiOJrw19Jdu5Q7sgZzXF4ckSstqqmxOcf0yP
axWDjs2wRCrQXdjIO3+sZsw3hr9g5WC8qb4p7R1bgZQB76/GJUJH8rpHprE1GO1h
rhHx4SmOkEHGKumCfyYrPxCakPLh4edaAibN3XJg+imciuE7Ou4JkNyefMdpMT/1
ndqJk39FT196vD5/Ic/gwapSTri1eUs833hgPwYJb8r7IUmVfpIceqDhvhXrq+kA
0bxKHOhCKMLf4Q+6uWP5xwVp3CSh3pz622/jEEfLLbudVL4T+1S4QnrzFhOLFQ/k
5nRawJkid7TXxPfnLFmbpz3MFlo0k6P5zGCL7JIfiNWa9sk00ChREZwW0A/Mkn6b
NPLbsQZJkPFuumKNIhj9fXg6wXX380Qk9S2SI0ntLKUwdyPUgFs2BRs6kfhnCWfX
CoOVzPKrQV/ATcQX41Tg5dcKEoP6r9e0wlLJ/gB0l/W6q8YEv13Cfrw33X1t6GWP
m//5Kn1TJPMTkAkjEwZh2W7pheAgfJAEP5az4F7Tb4IOq1eFglHUpKctCz18Q2bs
etX/QjcekrjACN0Rh5JMA7KMR42L5IEKDFT1WHr2Z+fi+4vJAkk43UQJ+S8Wnh4Y
VAA+iq5tIVKf5hYubmLzR3IiJY5Hn4K0a/MJ/lP79SVfjiHmu0Upx/Mt2bKGvtmt
gNHwED133vRs5nEgM3If0fAu7WtoU16oERYSmzzl4lqA65EbcllqjLCsWcPNQ3WM
Pbz09isYoObHO36wl6Vy9LV6rXZgfJU7yTdTa+AfiAKwk2FLnw+Ki07+tHGNdx7K
ZniQTuLSd3GTplOn/9n6E/k2Z8ARwXqf29mFtdNO1AHWLEjW78XCO5ZpV2slAGaB
Zf9BG5Hgey59EhoLe2Va6AbZvSDjdYpXg/AVj6D5BCGst8p4CG/aBKOW+4AYoTMV
F0EQuFd6RoXV71PgcGwtP7wwDh24Eqgb2kHyBVf45YuZzEueroM68ti1e6s710sP
bs03S8OeUFU05dvdwLW0CH98O/YKgKrdX/Rjkri9EJ4mCoMA6vYGy9FovJQ3in5b
UDADa+VY/rTAG8CVaQOyJxM56e9mT57cezeiabX6/sKPEGgSMArb4SVLI9jmqh+e
Nq/RNGuPpZhKvmyrn4H6CSVKF7ZQ444b4iYbc5b5XaDikxt1u5aeyv4rpweaikWY
aQCt/L9TWPXB4j+m5XjlzQA3NSWEGE9sqGnlSiL3Hp7/BFRpQlgI/DXuIo+o25qU
SjamvUOD6MJkW0DxmOLiYvpaWI/RoHpDRHobi1JESpnlNrMzEhzJ+Gkqj16xgYqO
vuPFldn/L8yvx8kks2qfygNOQjnYg7sbMpHgv4nJKZNRITsuCjKSazgNJS0owZan
gtbFq0QRV5J3SHzUkM4+BAlSVbVh0Gz+7s5hn1yAAb1gKAIC7S2+nta+XdEskm7w
uAzfc7nMnS+aeemS2obs4slIk+Lh1J+4GYXcKUng/iHVpADdKWRw7AoMLDbfMt6N
UD4HNTM/ibNS09v6/KM9oFbLdyEHJoBANww34aYyY7JsWISBrBy74OzGN0vRBf0U
BcipU3pWPEyIsGfNBexacJ0KsQphZs6LRXL4fYG1ZPM6UexCQtfKBhWrc6lev3gm
`protect end_protected