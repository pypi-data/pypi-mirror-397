`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzY2+EFIYXUoRGNXzJ9ubqwYWTSK67T3WPH3VcXrcvwHL
hGBB/qCkNnuJvFDccVepOl7v0GjpJ8H/iJSwbXWRcVA+AnDNH1T1TFn3VZyEx8v5
FPN+/xnwyRy2klFbPuCBGwyCb2ac4WaIR+m43LDgPxyTPn/Bupj8iERd0xyf1rdS
wVuP/7iX1ogR+5+6JaXOTIuza1vhbyZCfkyVVvMLttVBHvxEdadznHEtIG6Tr9CT
9HOx947jZN/TnAFudxPjRzh8fBihaZ4YGZbv7VMlFIvholEBQiMMxAAAejS64gny
i50gq5yWbT6zmUnnz8QL/ZvmzEyiPQhhZjEN5Ffa82XgrDZ12mrGELGws+/Ef0sn
9XnypqjJGHKULgbfyUK9Q1+/R2lv/0SPdb17TUzzn/FXHPpbXXOq5+4QXSwnaKjk
DXqcg1KgE/XOVNuibtTt3Ok4VP31z6UcrXvzvYcH42NiyTKd1S22ywcy7KU9/S2M
auNYjuanySkI3/3dP59Bf9n8N/cJNoDO6MVho3mV2MWHCjGcUzuCkGztMS2wvL6d
ZSaeiSerVCR6uey7aNWesRR+pQkfVSf6zxw2uqp52Amb8qaM1gIl4MeJOR0L7UO5
KhQZQ0Si3e8yD1fxA9NYCGMFiSxaIw54PQyil0j+cYp7x8f6BanFCnyCKhIH6oI9
Rrj9MgMBkc7kquSB44g5SZ8U1C7mDwPbvUKqeRkSBffy8HzMfCAqhas1gJmRvYIJ
WBUZzFz51j0AxXc8dCXwNs7b1+NayMVui0Y869JA5a7PmtowlYUHRaJd3s1EGdWI
zA+fhbUdeSJisr51kCFO7yx82wzBZZDKX2VsC11Ns/WXYwPlln/uZfWALhyftZMT
5euVNVZ8vEUgd+P/gAz+uAhZku8pOiChCfRAWTTPcXju65lIwBQUd8okClJX1xK5
x8okH7b0fkDi9kWeej5kPulYRjkIsXJTx+GNzaHOhiLD8G5T3lmxTd9CAGxCYGG4
AiIRawp8WJ/8EvkjEDELTPwrUm0SdTQmlkwpnUEsmqCoX/5huWYWJd4nsBwZqvNl
c6DEzjy8s5e2SeCwcXVLZCuUWST5eI06Or0pmByEBUxpkyyov0GGXJ8AMwOW1f4o
CNQ3+nikYdVdj/zf+o5P5wBf2VLhi0Z4CzVkcwzZBv/GqDpXiaFQPrE/LZDP0giX
glSW8ig+rNQWd7EePbAepsf1BCSZqLSECWoKayWoU9klgTKu93jLwnCgYPifYn+Q
oY0uYlIRtjrCfEOoQNVDPTkT7EJ8hd5WKWin+BaT8kV+K8WLDdr5wDWHqYHeulpz
usE6nt8udB/8UmHJ/g7IZdjc2SIH5Ku7BA6Qf3l6+uW8f6/4UJy6iGI++87X9loT
3MM8O6Zj3eZInKaw0Jwc6nfqS1jkn5gs1m0+4BCg5nJYzSvX260AHCuQgBFFTysV
1TYDDkROdJ+u6UUUpJF21qFWvgQfldPRO0eogfZYjZtFYbEyxCSZJSxA6TcbDLJV
STdv2CGfvG0NhXakOV2UFdcS89fGDT+ii30/SbnPpFYKSaTAWBr6x8c7OKw51dRq
4GeEGKvVYKw5rZRm7XmODfl37IkINPq7SQINdDuXmImFUwT+CKrjNi9VNareO9Rq
eYnkldOjR2/eAiumoxreBiodmkRo/+P5hk5wdq1zq2C+MPsPuQxuMV+UYXcWTApA
fMg6J+ug+sWND4aR5ibtufHsFRcVaUbQA5JSJEtNgFbH3skmZgn9hwNiWklSLxAn
LjLfiLBHdtWLYpHlrAeKsGIQ/zRK8gJVviuUgxZBrvVkWKFE5BI2EdqunAdbM5nS
U2O68Mpj8nZlqSPv2cVD8ReFriOSvi3qbSbHFhoKQ6RYuOcggNd75CKXRakmJrnR
oVXxk4p5xOsrQnK4aCXw1Vehf/O0pHuzDiE7R6WEUY5UYjmTlTScLbIKF8f3R6f4
TFqFAvXYJd2Z7cUSlLBwnWWHJ7RbT2nhvKUOP8R4ADbHlPFbHEz90saDwPjdCFpb
7uZgLmNumjyb0ZxLjCMa4BlPBwyILErz1R0WX9zmazy6qMVa8sJOY8fNNTHlxHjo
PMPlzFdFwJYsi/Bdqdtzh4ezlh6kD7JKKtKR6rjFNAZWGMKE9vbe2nJR7QRwqNqE
gIadA1vWLG5aWDoAuo+NetrIOrEls8Xdyq3cI7zOczX62UEWcAGDarLt2VHRa3ac
jNAxapFjHL/YsRhfBTuorRuNZgku3qRpjKchUDLkwFHP8WosAlD2DsvbYFy8HUVl
ws8IoNku/wE6XX3DkzDa/5g2Q+3i1iymE1qMmsfkOexFss4unopvymPqG+ug7OFu
iKYMvAs4cE6w55DapIpnTgPTPKvjAz+b11tFfG45UN3RQEiH2+CnlODWvuPA2xs+
WIlyj31n5tCeHDbsK/lIvA01pImqOXPOMgtJhQG5MO6LkeHNVtDnrfV0BJi3Gj2I
yPAWQ5KDk/bULbIIvqxzZQAXrd8EOJTYMjy9Ji8eWpivXfBXPLwco0bg5S0rTdG4
pgZA8PL39yD7HaL1YXVBpXwjKmK+aqsTxp63DmMwEuwMd3uNMYRJl0EQPhUq4Euv
fDN5vT+HjTUNveU2VmtfL7ADJ7g5K5P3eptXfkKKuWlCqBz/vAcB8vIHRJvXDa5L
tWvE+SfjjOpAnSRlL36u6kI6VyUl9rVsKfUV1KncPwr2xeP/w2LewGPxnwr2F9oR
BeoHbprwi/vdJUCAzlPDhH6qTy7BfGyrgMe0vtu01l6tewgFQaW5iQExLtDrYkxr
J+G+3wfmX9b+q9fxtOwOPUxuORGylNeF/W0vt289dkMADagl1BWRoZhAHH/2wpq/
eDW3pQj++aV33/iwzA/GKgVi2qycR/2gedI4LINevVZqAsnmnS80fNBF8aDe/3qm
KoLgkMm+4Dw6feoqr1t5/yXoRRBjinV43m65NvpucOWV2QWPQLejyHg0QHdzTH7q
o0UXHnOIOy4QZgcehekCByOyAojyvjNlb7A3Vjk3FTaVVhOFn2XirX2meJWLwo4e
h20mSn2jfmY/OJGnFDLHpTXTOrslNbNWXUaf31eNW6zxF2hZ/MbbrA23uVFYsd0p
dkg8msUjVwaH9fqqcdy9ThqflrBs46eDjmcc3NxQLOo2RwZTmuhZX9xCU+nTcVmy
DVcKz+/RbC+0cvghMBfGUWlQeOhCDf96EBsU78Ym0wA3hzAbk7/L09rMUogw+qQd
fXsk1fstzlJr6a1c9rkAUiJxMpAoWxRlGloXUyIMP5qBEHl88G70hnFVH/RurI3I
svsxMvE+Kd1ryH/MiXklZmZNxRXnlD/3RmKTJD87WZ2DOchp6zz53ACHIri8fuky
gXTcIvlujK1r4/xU1GDLH4GXAEPRtNUb1ZYqXxZOd7M75MdlHZtHGyAn+t3qYOXA
EZuslS8ukVF1NxAkqcilen7j/TIX4Oc5ZOJOIKJZg65c1urhAmbOiG4ACzAvLm9F
cmzcbUD5AaMoxIiCFATggQK9Zse1q02cEMvG4u/4gh/Kveql3ZroCXXGkFHXOpBS
+/UUJ6rcy7x4jfIUMQS3NT+cDW7HIJiKw4dC73Y05WJ6TFnKtbqM6JVvmXlwbsPr
W5/Ies28q8UgG4VnWgoD23q7HFoilCwOEIH4RQTTCuenVhHhtZDpw6LsZCtweuAc
YbHvDvm6GyOe5+gFdfBI3IWt00FCBqbv+vtee4/Ui2ZABVuR35K3Lk3XQEJU3HAp
UzeUKkhg9tMthbviYSVdvgqS6zJPvfVtXA1Hi0P/B5Yd/RjwjtDesH9tj8k2QBIA
FA6zEpw7BnfMhmBJT6hhZ8JXot0mxEoCyvTgGR4rbyxi56/u0HdFKOdl1dDtlFv3
85nBORE+eKqWfRehdgH+dLDp2u+7rzJl9odcdLji6Q7XBy08kEa8xE8BXk+zYbJN
4Ht7aA40Gkf0blPYZD2gqM8E63j6SfYWfpkV/ntgwtCCJ75nKy0KXd0HyZwyzK1V
2/T3B3I//wSTHpTULVxfzWsegNXNTtvy5OO+CV+zprWnSC7WUdP778UHXMnQ08CN
vsmjzpMnEjNzVFJC0CuKis0dW0IgRdGw+UvkiY3EmB0Thu1Bdqh7GfMyJH0vvwZK
/3I7kIXGuNHpo34RHUNHJSpym3HLLLQanM2NIWzodLqlqbipxGSgSfx34mbEp8yf
RPf8/ktutCgQIXyUp5fG6Tsknwtd8XffeIBcwKlEmAmtAC5FtoOQc6s26fhSTCs+
veCa4pYpzCeGnf/qbbj/LP31bH1EHrlpa8idKqL1lNnMxlwPurCWZDrU9gVhzNab
mV5ZU88D842mnWl+ZIy+yZPI1IgoErc0LrmoLv8sWtgeRjfoNHkOZGas0uhSp/qk
Z3X16M5HfduEstmEX4a9c4rln40OtYMi6bTQhM53XuFvVgF/hG7c7wlQYpx3Gugm
Jrlcfye1c0+Tci5lqDBfwxxTWhX+YlbE4tcnJHCpMkDuwjs1t8jWgPR/QofDCDBU
PLZMaPBM/4ZwSONJL1vqPgyjIZZdSBZXAXpcydzyjEeiwnWV2jKWFbi7h3V827T7
zgtIqoBVUsG3pTChNJNDPM0CsP11me1gZZ3zykQH3YDf52ltCfVZNfM5yoWbFf5G
62ofeZMhjwnonHsL4HFQu55KLHgma1l4V1RAAe3eZvVmIpP3iZUOvgYSDPci1svp
sWTg/ZM9xyrH28hHDNZQwK4SCUkgt7xlPc1rCnw4Fb6gduQrPz5CjkpWlOCUrdGM
dsOPmBGmsVBbZXMmEU+4kne90pOFvSQ7k5bTZByRVzP3idm+QBn00tbmKw6A08VS
5Zz8HB/a6oJeVm4iGnG125pxxrSJ6ycqkt+S2HLVLdQi7JW9GqllR3X9N2l8RDVS
Y5TuRnvx7SND0NnXQeJ2zUPc7elaEvuuFyj0tMO5Yo66jvbtgSMTFotpHD1/cewF
6z3SNZxG2Zeb128UKyGaHFITfGZRUXh3GqyUYipSQ3fcvLmljR8vX0aP3106QefB
2n5WJsfxPnLxuNG0FW93rPmNY1MuULPmiY36oUXPvYXSPwXE+brBlc9fuCWIV+d+
cM1jWegCyVtoyKhRS+IX7qxvmynSNlwD61N6qAHRoIvgrbBYLJOJao+0PPRM8oMq
iehmeFk6RDQmxIrihYK0RHQmra1/+cGr8pLO4VqNlvAydhTwRL4GcACmzWc58c6C
LarTohC4YZgBpv/QnhHlSq13DepAB3hqskyySYPFI/FDWDRacEbRZGJaW2KOqwE1
SrpqnwlLVU5nQ33oNzbfQk1Of+PSwgcdr965ZxHenOpSL9fCRNGs2Isz4L3t0fVF
yiUx+jh3NAchf3hyYsIsYDnTJbfcMN6cThbVCuwaGQJ9KrtINCGd9vpsY323RJEK
60ky4qPmAjAmEEtppCssNDpfHR0+R91sXaoI8BZ+lYI+sKbhs8M56pfXmqxsKAMv
f81vnxVOHjmfcy0lX1j/Ss0Pumv7mtiq0aW4qamtetTy9T9fEI3wKuJsqfhEzNsZ
87WFb9OOGm0O1qUNEhn8gVif+fmShjzKo6QsGD/iAhtm6xbY6hUrRY43yXdF5mXh
K2yM7eRds6G3AFFH/rHJBhJJB7hX+PUu3ahq6CDY6g51s0hU1w+0OLKRsrs8oxR4
+8arSsSlKgDzQ4vHKx2mBC4NFduXhUhBnM+4nLWy4tAU13mnB+L5AAZIkHFQEZ2C
TEXau8/KxA8CVwZwX/YjYa9Qu3U68X3l2bLl2mlpYn9GJw6eiubz4l6sQ2FDu8No
1RWPMv8lDHbwOuOenVOunTZumLcZA9fowxvLEE5+gcJ/GXrm8jTKdqV65SF6an3v
dS9KHIxHXo9AfBGMGyw7NTadF4M4WztS9MvRZtt0xciaXd78BasWbTcLonsceRyv
atPnmUaxTLrMxDn6qbFDKt+DS1Fe04XcS+GPG6PhqomRgdG+/uS3kHrF+PR3c3eh
tF0vCDk4Eksu5/Xg/IPjg5410H6c6Mz1EYothmnLNVHTew5YORAzu/uzzyJ7ClXZ
ZBQxiK0frBQPdXWq8h8ZqSLoZLnGGnSZTqh2hwgnHCVu607d6swfM9O6nINt4qqa
s1O9iJnhPIfCY4pbKSWvIegIVh3262eK117AD6DDurVBaqk0VhBaS72vVE8IKQ1N
qhRhOqnOpPWI/q3nSXXQs+Js0qMsUVF9mnP4APeADqyOfC23wDhvQoKNdcFmnJa8
0hErCqItVDfxGYFiRe++kheBXLHBh1hrS/2t07j4kIZIAfsxQ5VU/vvtSFUegBwz
EB9385nB20PLoxZ+NJd6fuDARaji9WI4As8YeFZ6H/JykCA0unVardB9QDo4umUP
DrP4VaqTOYNC643KDte29CzMB3OcoDSWPHcm1rFSzb4o+ZNXFrL3DWenM+PPDjIf
eBJBX/0Vb44BH66sxZXxwjnaSO79EI7eIsBVjFTNJhtNZZDWSN4+4+zMqPA0+loo
GqDsQOnApY6qe0SOtpJ6/Xku1TRsTZCLcstXZD1hBaFdC04CD8dANtXZ5AOzi2gL
wWp8FmqK64pL05B/PkBLZCFBYHH6RTzGT0Qabv0WTHZv3/c+dcHegUbiR2Uta6lu
Iqmipg5QRAzc9Oa9IU8AoNe4jCTJ047DsjyWeR3K8CYIBKN8SD1kSitrTbq9SgfY
syxg8s2mMCEU+vxSaPn9WyNPMrU9TWEhPyvOzmkvY43Fr5+SRZN9OkeZMtZ0l8/7
G4hTM7G+3+1f5jfuXwjIjkAsu2VO9E2YBpW4UZb62YBfmJN/BQLZWwj+qtKIxs34
ia+KlPTY1SdQ1rdVgRcf2TfUFSFOpuWGTTil8B8B10Xdl1KjLkshXXFfOR5GXrid
dViXvmYKVSQ/3OZtkw+PSwoCvh9XdyWSDgdWclKnnJUOoFrBNRC4pTtQAf05nE2W
HzJwPSnaK7LSmj+plxPVxSIuKiO6GtQUAWZWRWwzeV6PvYzc1Xwz3st23yPvB0sY
tKfQpIUdBnikTUYzPl+58JOkQr1aDIot+0CItuzAo8B+s/SqQBUC0CwwR+q2NVDs
pnAFpNHoDqeWZqMA+9vIU6PFx++oQVez93I3uD69aSuHNHUXtHWrgcE/pQwodz17
noBErYuXu4Ms03gYV2zbkTO6PXrrz+NeSqYQtX/Paw2XLWWfdwDVNSBk6yIvuf9P
SF8SpRABbdsz5Z8M8QeuqC04WiV64MqRH4geoCSS13c/BGghtruIWNEKyLeR/sXJ
MpLrk1QW9BqL8xTaG/Rz8FW9mgeSMglFo3Tt4Oygtnos+XYGchaIUV287tfXLMz0
lohyO4nCsJuK60oVQ/gz1ywZo8sL1eMRZ8a2Qofz2dJN+1cgyfQR14uBjcdpN4Kc
SE2VZZ+Dltugz4CpClPs95EAbE6VFGEOaSjysgQ6qV6DkfTNk2JqyAHBnFSdABiw
ttlK2tIRq7qCH2xLNunU3JtRrup2QValRDVsT36pOzJts2q+j6vg+v1Z4y2Ix+c8
mv0HJKkRH4v4YTdz9Hag54UqTxpe7pjslCry5syu19eprvLIBUQo44YEW1LERcuD
+O5yFkeHYB0jbai2Nl4h38I30Jpz7luYDnTCVXhI99F96AeUOSWG1ERG9txmtM4/
86HJI8TU0kioFvUWY7iEK6P0B09nxqOig4/WLfthHMXeoNYBYg+xXMj+13PVLFRX
LCfl2VZ6xNxskeJFzn2oAl7tzOGr8vSboQo58KY+s7YRRsAo0gZVMYKkAZGfg2Py
Ayb+2cDhkSxDeyWshGGs/Ey4ssEviMKfJLaCqjfIkFi06S2MPus/mxM/8tu4fMJ4
lYfSo4AIPQgozeFoaN1036A3OmCdRGYYRMuMMZL8zq5bHQnkBNett2L1CSErACn1
cm0eOwAGc4KlRooyLoaNvkZ1+k/7zBFnll8h16vTrr7ompAr7SuWWF5sE3lNhZGN
8iXt06BiZYJ1rHb3EcvxDXCWqOpeVk44/RuspcfFZDz3Jh9JLyEahUhwyYFpCcZQ
J5cqrGgraLBaJCFwi/r5s1ltBBRoEw2iAR3w1y8c+x8YxwXUZqyEjDMlegrWGutv
Y3xPfLuLNGYj6mCdpu6Gw7qKDF2q/ZurpkT9y3mxVwbqy+NVgyC2Zj7nNjXTLsPB
UCdH7bH/UvVRYSDDHiD5Q/girpt/0WM4nD5WLUhg4rAPeXmeUbCB/C8xq0fUOwrn
HeNXS5GeBXssvCqKdCfgHkk6gpGOQfFH3a6zxYA9MjXJ3xCx8cgCXLgHYw+kux9K
2yXlt8MUTQwAy8vkLCR64j8eIV9ePqbxhOSSAYOwgQ33Mezi5ixvJhK2Oyzo/Rxc
urY+R7cXd/H0AH70W0Fc/esC4e6yrtFcvLytMnX6yNC6cdYVYVBrZRUm195pNsv7
4eAn2S9RMBO+gdVey9wFnx/QsFnMm/l6T4LIBq5nFJtcYc4fYXOkOub8g+sZfXRX
kAdute+LRZKt4+Za7Bedm8VvITsL+K7u0/3OkqAPokeNza1Pzfw8G6nOl/fJIvFt
fRQn2/jGgSsgwa161Cp4rybjkYa+W/F0vMx9DipD50FyPVp26jdC+2i2cLEx2sdF
EBfKPJgbBB83x2O+LUIKSnxvO81NIaSzW6/+KOFY/cmbV2PNLHcKMh6XRKPqlgQ0
SokEF3a9lz10VAVv7tVSAl9zopUzWH3XVZpGiHQZpnhSFQeJSNevbZTySl33Qhag
5+HyFGTh3MWeZlzX1ZXEqfQROp8N66W/bPxcM7oG7H3pfnMEeoKcmNKy7L8DPb5F
Gf0umQFTOeTUuWiThJUUnrU8ZmeUNplmdndcBbZseVQyeun5q9ObaT3VJ/34seku
m3rTr1jI7UUMMFUNazmEtb35PjY2YQRoHN/QQDOixem0p37lv3T8hCO0V/YKxhd3
vxN0bMXFWuiBmBI6v+cw5KyXSoOFaF/F3ldHjPbsASWzHzi/8R1MqKPztKbNGOlk
BtPYKrfHTFmACjUrUQKCWomursulwJHJ7y416tA8yY1faDTcChcFqEm4OML/l69h
U8ZWGkNZYz4E79Ya4mT/VNwIS79QvWmihObJ+p1c6HiSkBvr0Kw87NR9t70pWUYZ
hFuwilPWW1Oiy2pH24MJMgFjW8Ri71KwG9C9/bIFI0SgBxz5B1voOT5hdjJ6Rfzj
NLqCwU7VEuXB7ZrWBf7UsYM2bHgmDwDy1ZkYhkkl2Cck7hH2RYyaI5/0kh5p+u43
W1f7Ny8aiBUn9XVUUotGEHCD9+AcVfLkDtUKm2sv2vGlpCqj1gXFVFuz5ylJIxTP
z4XDEn4MSABO+rMCutGxzp30ZE2S0o2M0s4PRvPbHMUe/8c7VmcghowXNMz85DuX
RcXt9sp4HpKPvjMZOiUMW8IrErZ7xSUUQoBPXiwS4iF461icbpaGsKHYHeEuGh2r
zvvAcKBiU5A1GFCLfqRXJC3ST8Br9Thl4oF57jnCgPLdW30pmHObLH9uI3cMTVnV
/a9nCCFgk4atA5nlhQc+q5EAtvs0ApMpXdhTNtynabpObl6F1812JOVBYPrWRiqB
GkKsOl2NihUPKGv5iREuwnHKNywT3fFxSLLkG1unA1hrs99xRwVYfRHOiLTu77/m
0PxWkPI+QOM05xk9fErihSE5fQ78+dlidFREBwiqF0jNdgZhnWbzjfuteCeo2SJT
bgRx3cs/jcLRcHyd3C1KpQMU0+GH2Fs8AYsHdYWEJJu/8jpaNYs5VA7C31eCAAqM
VeXIoP9NytJlq6718uf7KkF5nfznjNdsFRCY/TRAF77gEtlNDamhIIznCJNYaWeK
7V2mGKecuFCIn7I/SgD0XJrcSWlmOOyKAhP69+QwJe4M7zWQQrMBZh8lRBWUuBEs
lL42LwAH8XzZuhF5ZRx79B8kQA97drVPHLEVa+T0C2prAXsgvau2LLY1JIKRrOxr
n5O8LLsR8WP1tJu/OLHVChSGDdR83m6OS2lKxxzkHOzzdNxiCjvYmkd+9cMRih3A
rgFmGNAxYdiODwgv3nCABob8wu9AuSm1gAUtbaaljdQHXCm4Y7bUHDtrBgtTL8SL
u1x/54ioN+WKFgIULU1bFCQdPKklwdq51NqCb6uKM7Er0kFaaufB8yRZFRzAQNRD
Gh52Vh7z58V3O31uDne6uJAPJ3hAGCaI7RazmHj5h/zXhvdTaPDbAEzb2k9+wVW/
yCI+3eqdixaLxrS7sEET4n84AEkPdvRD0a6bVqki3j/Aqr9qosgIdcB1pL+I46sj
G8KfhhLLuQt3ZTRvP+OnvATcenE1yJDNd9rNFu/y0Z61hJexv30jEnM4r5d2LBbF
7mMbrhG1e4FMny4bklE2RBLamZJQStrv9mhl1tjOEZl7J4XfWLDCehepJbZWut0f
2VidI4xs1m6y4x5CAQs7NWGiHsU1jQnkNskirS8UbPk92J+xDSjqRziUFpg4KFxU
hRWykQ3v3nYBV+uEpc0ybCzNKlCb0jLmewTBWh6RHx2KzPjgZvENrSV7vZ8paPPr
Tj9HHraoFeWSjxmezRqKIrDAHiqfYwJwwSSqmaKaSyRiqt5qw+4IITdwLq6J6+na
URvG80HE/Vskx44Jjhgx+a1RkXFGyNedahzy3xfn9mtNpEVNgPD76LzLSmnWbm5K
08pchYWTpmID5dCBnn9FSAohwb7Y8Ir68IQWwfh+X4DtAfaierthAOOmfEMrwWBw
Ogo4LZo9I0C4mZH1H+R/Ob9MhvaWRUHEALAJ2ldA9PTesyc2AnTASFhFm3X0ZyNp
WOjjqbhzZTsMY5RM0rtMww6kzCp9Cs68jSdaaLQSNMSK8pDdwYj8Xmj+AsBCulDj
E6HAWxhX5bSKl080jprLGWYO6FRRITTGSSJTlhKyqc1uDj2dlBrKuIDLBC4aJmmo
jjM4yGWVB32q944vqXeF3PO/AhFyEh5+KOmpdlLeBT+6YigmJnpuNbgFv2OcesLX
At6RJ5PYu6Onv7hUKd7tr9DCql+9Dydqu2dB4dccXK4P7zQhZ1NK2lhqLNIXIc6X
saYFE7IDBGg2alcZdYrq/yTY+uJD3yduUes8WF9HcAx2FbvNkn+lxwRAPJe7+ZqF
ODiHPMbqbVjate03Dg7pWFKQir0oy4XcQnOnSqWUSY6RrLeiKsY0kUaikef2Vs6z
`protect end_protected