`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
Hm0rc5KfjNwPmEU/4qyz3Shjke+cIa/GCneKewEXB3n2bASaGijv9rfRnH3PBHb8
8KdJ8yt7qcQ30yDODGzaXnpDbFJ13UvhDClrJXbfQtKGvC+Um8ge7tkOyPrAgJuN
h7tF6whetxx+3SBG08B1XE6mDgX+Sux0C5lV9foZj6/WYH8vz+fdrphOzw5OyoDl
KknJeLMrK7HFwv+NRTZU3uyMqf6gILgsgh7ZGfvNSKt89EVRddaUKOyTdcUZ+X68
/D9Pfq4aa6m3r/dHwZe0boZera1v1IDvdxh14xErwEbeixbral0UpDhX8P8tkQTj
h416Jg2dVlprlNF2m7SRRgCDG9d0Q+vpThl9byxaabQGuz0JbSWP26laufPg3ZTR
DKZiCH54sKfFya4thMLigOOBQay1XgeNGHFGBbtfHkU9AkF5vC1MXqgWaB2MRpBm
p0BsvPidEABNqMS7EF3z8ch4RrzC+9XUUrNRGC8QlRYT3wcSuH1CvAov+UE8tlV3
JF1cGVetXHhqt09UGYBO65D+gwWc2lQDpTR2fn4CImnm6InUjdmPV8n2+U3ELKuc
Vc/M15T7oNQXI+K9m38buNo2rw9clPEK/R11nfU8Fe5gjQxS88jB0oOXGhRcQMHd
cHuHEGaGX4Zqd537P2h0JjyMZjZxaV/ir03JvaJOZCU60brZ7YSm8ocFKE+JB0wE
j4ENEj1jbwjwHRHFSqkGKIa052TZAnfKDmYkGgmVyqKqEPv3rznUS8b/HMleWHE/
05GDl+ILOOIelVJy9eFG/CDmzT74y7GY2CH11JX+n14IdtltWN8xeosIKj9u+z7X
alARSba6TV2BCsVQD70dbXrq0o2UK9B+LT62hDTRgMdV0dvP5PGq24+899HUkVLb
lkYFxJymfdqjheQjgopmhfP+PLzJtLLkZdYl2IGBvSVq9EL6YI8/G3jlcNkjl/z8
sCguJbDfOtKmKttK/qxu4MS4PLdheQ2oKBa0bPMGLvxFApu69exVCDC6W4A/sWc3
4v1//zNUzcUARE5C7ZKrFPbYwqX+uLps7g6Ac1joo7x2LsW1C3PdrVp4T0rUZ6+u
jsbEm9aIhcapvUj8lds/xoL+hsDDrus6wgOFOt4tVkTiHKuYdc1vJNYPX1ePjDxI
UOd4XMBB99o/tu2k2uHOYIBgZ6kSUxK+27cWtoaouKRuIVwIN0/k4rnSr/QcfndJ
mK3Of1wIMQEUNS9nxy2GBk3/ZXeBGECckW2ssp33S0NoenWB7BVcLUUSChvUOubB
46RmAlwBRzYuz+1VDhMWmHJsOmVqg/SCaECiYDR/A6PMF8KKyR49m9XYTkYI9mvU
lQXhZ8b34sFd7jxctRRwHvlV56d845CVQJgN7CMXnseFyxsYXnI6TQwvDeziRmYO
D+aiNUYPOkkR4OF7wAlXydJfvAK680jnPJxIJu8nAoI4aqG2hPFQ96ju4MyzGgVv
27ZwKdy+IAq8Yd3Ad6SnTSo2GzOpU3KttSA4FvSJUD3PEL0a3S8cnQZ2hRcA+ePF
cHzbpkgZWOI3tMfUtggqcLEAuV7a/IMR/+u/gYiLg9igA7M3rEXKhyxIb6Eo7mLu
iSKqwYPKlQz0UBft86ostTeuRiXyaApZvZweCJ85LiJWe1ZxGwOu+73xTPlI7zy4
EeIFHPoV/K4gpQx9DR+jyK68n9sfII9HEl9DpsLpiGTHOrbTKJpCf6fupOF/5X3d
1sK24Gt2gdwVr98n5EBLKh48xFdJP4+wk94Xl9DiKcNB6E+sPt35kfnFtAtUTLph
WABwrhLV+uFtOHdTz8Fi9g==
`protect end_protected