netcdf testoutput {
dimensions:
	latitude = 180 ;
	longitude = 360 ;
	vardim3 = 12 ;
	vardim4 = 9 ;
	vardim5 = 46 ;
	vardim6 = 18 ;
variables:
	double latitude(latitude) ;
		latitude:FillValue = -9999. ;
		latitude:units = "degrees_north" ;
	double longitude(longitude) ;
		longitude:FillValue = -9999. ;
		longitude:units = "degrees_east" ;

// global attributes:
		:description = "" ;
		:YAML_config = "grid_settings:\n  gridsize: 1\n  projection: conformal\n  lat_in: latitude\n  lon_in: longitude\n  fill_value: -9999\n\nvariable_settings:\n\n  - name_in: Cloud_Top_Height\n    name_out: Cloud_Top_Height_Day\n    attributes: \n    - name: long_name\n      value: Cloud Top Height for Daytime Scenes\n    - name: units\n      value: meters\n    - name: _FillValue\n      value: -9999.0\n    - name: valid_min\n      value: 0.0\n    - name: valid_max\n      value: 18000.0\n    - name: scale_factor\n      value: 1.0\n    - name: add_offset\n      value: 0.0\n    histograms: \n      edges: [0, 1000, 2000, 3000, 4000, 5000, 6000, 7000, 8000, 9000, 10000, 11000, 12000, 13000, 14000, 15000, 16000, 17000, 18000]\n    masks:\n    - Mask_Day\n\n  - name_in: Cloud_Top_Height\n    name_out: Cloud_Top_Height_Night\n    attributes: \n    - name: long_name\n      value: Cloud Top Height for Nighttime Scenes\n    - name: units\n      value: meters\n    - name: _FillValue\n      value: -9999.0\n    - name: valid_min\n      value: 0.0\n    - name: valid_max\n      value: 18000.0\n    - name: scale_factor\n      value: 1.0\n    - name: add_offset\n      value: 0.0\n    histograms: \n      edges: [0, 1000, 2000, 3000, 4000, 5000, 6000, 7000, 8000, 9000, 10000, 11000, 12000, 13000, 14000, 15000, 16000, 17000, 18000]\n    masks:\n    - Mask_Night\n\n  - name_in: Cloud_Optical_Thickness\n    name_out: Cloud_Optical_Thickness_Liquid\n    attributes: \n    - name: long_name\n      value: Cloud Optical Thickness for Liquid Water Clouds (Primary Retrieval for Cloudy Scenes)\n    - name: units\n      value: none\n    - name: _FillValue\n      value: -9999.0\n    - name: valid_min\n      value: 0.0\n    - name: valid_max\n      value: 150.0\n    - name: scale_factor\n      value: 1.0\n    - name: add_offset\n      value: 0.0\n    histograms: \n      edges: [0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 60, 70, 80, 90, 100, 150]\n    2D_histograms:\n    - name_out: JHisto_vs_Eff_Radius\n      primary_var:\n        edges: [0, 2, 4, 6, 8, 10, 15, 20, 30, 40, 50, 100, 150]\n      joint_var:\n        name_in: Cloud_Effective_Radius\n        edges: [4, 6, 8, 10, 12.5, 15, 17.5, 20, 25, 30]\n    masks:\n    - Mask_Liquid_Water_Phase_Clouds\n\n  - name_in: Cloud_Optical_Thickness\n    name_out: Cloud_Optical_Thickness_Ice\n    only_histograms:\n    attributes: \n    - name: long_name\n      value: Cloud Optical Thickness for Ice Clouds (Primary Retrieval for Cloudy Scenes)\n    - name: units\n      value: none\n    - name: _FillValue\n      value: -9999.0\n    - name: valid_min\n      value: 0.0\n    - name: valid_max\n      value: 150.0\n    - name: scale_factor\n      value: 1.0\n    - name: add_offset\n      value: 0.0\n    2D_histograms:\n    - name_out: JHisto_vs_Eff_Radius\n      primary_var:\n        edges: [0, 2, 4, 6, 8, 10, 15, 20, 30, 40, 50, 100, 150]\n      joint_var:\n        name_in: Cloud_Effective_Radius\n        edges: [4, 6, 8, 10, 12.5, 15, 17.5, 20, 25, 30]\n    masks:\n    - Mask_Ice_Phase_Clouds\n\n\n\n" ;
		:Yori_version = "1.3.5.dev0+g8cec38f.d20181204" ;
data:

 latitude = -89.5, -88.5, -87.5, -86.5, -85.5, -84.5, -83.5, -82.5, -81.5, 
    -80.5, -79.5, -78.5, -77.5, -76.5, -75.5, -74.5, -73.5, -72.5, -71.5, 
    -70.5, -69.5, -68.5, -67.5, -66.5, -65.5, -64.5, -63.5, -62.5, -61.5, 
    -60.5, -59.5, -58.5, -57.5, -56.5, -55.5, -54.5, -53.5, -52.5, -51.5, 
    -50.5, -49.5, -48.5, -47.5, -46.5, -45.5, -44.5, -43.5, -42.5, -41.5, 
    -40.5, -39.5, -38.5, -37.5, -36.5, -35.5, -34.5, -33.5, -32.5, -31.5, 
    -30.5, -29.5, -28.5, -27.5, -26.5, -25.5, -24.5, -23.5, -22.5, -21.5, 
    -20.5, -19.5, -18.5, -17.5, -16.5, -15.5, -14.5, -13.5, -12.5, -11.5, 
    -10.5, -9.5, -8.5, -7.5, -6.5, -5.5, -4.5, -3.5, -2.5, -1.5, -0.5, 0.5, 
    1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 13.5, 
    14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 25.5, 
    26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 37.5, 
    38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 49.5, 
    50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 61.5, 
    62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 73.5, 
    74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 85.5, 
    86.5, 87.5, 88.5, 89.5 ;

 longitude = -179.5, -178.5, -177.5, -176.5, -175.5, -174.5, -173.5, -172.5, 
    -171.5, -170.5, -169.5, -168.5, -167.5, -166.5, -165.5, -164.5, -163.5, 
    -162.5, -161.5, -160.5, -159.5, -158.5, -157.5, -156.5, -155.5, -154.5, 
    -153.5, -152.5, -151.5, -150.5, -149.5, -148.5, -147.5, -146.5, -145.5, 
    -144.5, -143.5, -142.5, -141.5, -140.5, -139.5, -138.5, -137.5, -136.5, 
    -135.5, -134.5, -133.5, -132.5, -131.5, -130.5, -129.5, -128.5, -127.5, 
    -126.5, -125.5, -124.5, -123.5, -122.5, -121.5, -120.5, -119.5, -118.5, 
    -117.5, -116.5, -115.5, -114.5, -113.5, -112.5, -111.5, -110.5, -109.5, 
    -108.5, -107.5, -106.5, -105.5, -104.5, -103.5, -102.5, -101.5, -100.5, 
    -99.5, -98.5, -97.5, -96.5, -95.5, -94.5, -93.5, -92.5, -91.5, -90.5, 
    -89.5, -88.5, -87.5, -86.5, -85.5, -84.5, -83.5, -82.5, -81.5, -80.5, 
    -79.5, -78.5, -77.5, -76.5, -75.5, -74.5, -73.5, -72.5, -71.5, -70.5, 
    -69.5, -68.5, -67.5, -66.5, -65.5, -64.5, -63.5, -62.5, -61.5, -60.5, 
    -59.5, -58.5, -57.5, -56.5, -55.5, -54.5, -53.5, -52.5, -51.5, -50.5, 
    -49.5, -48.5, -47.5, -46.5, -45.5, -44.5, -43.5, -42.5, -41.5, -40.5, 
    -39.5, -38.5, -37.5, -36.5, -35.5, -34.5, -33.5, -32.5, -31.5, -30.5, 
    -29.5, -28.5, -27.5, -26.5, -25.5, -24.5, -23.5, -22.5, -21.5, -20.5, 
    -19.5, -18.5, -17.5, -16.5, -15.5, -14.5, -13.5, -12.5, -11.5, -10.5, 
    -9.5, -8.5, -7.5, -6.5, -5.5, -4.5, -3.5, -2.5, -1.5, -0.5, 0.5, 1.5, 
    2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 13.5, 14.5, 
    15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 25.5, 26.5, 
    27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 37.5, 38.5, 
    39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 49.5, 50.5, 
    51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 61.5, 62.5, 
    63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 73.5, 74.5, 
    75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 85.5, 86.5, 
    87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 97.5, 98.5, 
    99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 108.5, 
    109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 118.5, 
    119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 128.5, 
    129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 138.5, 
    139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 148.5, 
    149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 158.5, 
    159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 168.5, 
    169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 178.5, 
    179.5 ;

group: Cloud_Top_Height_Day {
  variables:
  	int Pixel_Counts(longitude, latitude) ;
  		Pixel_Counts:FillValue = -9999 ;
  	double Standard_Deviation(longitude, latitude) ;
  		Standard_Deviation:FillValue = -9999. ;
  		Standard_Deviation:long_name = "Cloud Top Height for Daytime Scenes" ;
  		Standard_Deviation:units = "meters" ;
  	double Sum(longitude, latitude) ;
  		Sum:FillValue = -9999. ;
  	double Mean(longitude, latitude) ;
  		Mean:FillValue = -9999. ;
  		Mean:long_name = "Cloud Top Height for Daytime Scenes" ;
  		Mean:units = "meters" ;
  	int Histogram_Counts(longitude, latitude, vardim6) ;
  		Histogram_Counts:FillValue = -9999 ;
  		Histogram_Counts:Histogram_Bin_Boundaries = 0., 1000., 2000., 3000., 4000., 5000., 6000., 7000., 8000., 9000., 10000., 11000., 12000., 13000., 14000., 15000., 16000., 17000., 18000. ;
  	double Sum_Squares(longitude, latitude) ;
  		Sum_Squares:FillValue = -9999. ;

  // group attributes:
  		:long_name = "Cloud Top Height for Daytime Scenes" ;
  		:units = "meters" ;
  		:FillValue = -9999. ;
  		:valid_min = 0. ;
  		:valid_max = 18000. ;
  		:scale_factor = 1. ;
  		:add_offset = 0. ;
  data:
  } // group Cloud_Top_Height_Day

group: Cloud_Top_Height_Night {
  variables:
  	double Sum_Squares(longitude, latitude) ;
  		Sum_Squares:FillValue = -9999. ;
  	double Mean(longitude, latitude) ;
  		Mean:FillValue = -9999. ;
  		Mean:long_name = "Cloud Top Height for Nighttime Scenes" ;
  		Mean:units = "meters" ;
  	int Histogram_Counts(longitude, latitude, vardim6) ;
  		Histogram_Counts:FillValue = -9999 ;
  		Histogram_Counts:Histogram_Bin_Boundaries = 0., 1000., 2000., 3000., 4000., 5000., 6000., 7000., 8000., 9000., 10000., 11000., 12000., 13000., 14000., 15000., 16000., 17000., 18000. ;
  	double Sum(longitude, latitude) ;
  		Sum:FillValue = -9999. ;
  	double Standard_Deviation(longitude, latitude) ;
  		Standard_Deviation:FillValue = -9999. ;
  		Standard_Deviation:long_name = "Cloud Top Height for Nighttime Scenes" ;
  		Standard_Deviation:units = "meters" ;
  	int Pixel_Counts(longitude, latitude) ;
  		Pixel_Counts:FillValue = -9999 ;

  // group attributes:
  		:long_name = "Cloud Top Height for Nighttime Scenes" ;
  		:units = "meters" ;
  		:FillValue = -9999. ;
  		:valid_min = 0. ;
  		:valid_max = 18000. ;
  		:scale_factor = 1. ;
  		:add_offset = 0. ;
  data:
  } // group Cloud_Top_Height_Night

group: Cloud_Optical_Thickness_Liquid {
  variables:
  	double Sum_Squares(longitude, latitude) ;
  		Sum_Squares:FillValue = -9999. ;
  	double Sum(longitude, latitude) ;
  		Sum:FillValue = -9999. ;
  	int JHisto_vs_Eff_Radius(longitude, latitude, vardim3, vardim4) ;
  		JHisto_vs_Eff_Radius:FillValue = -9999 ;
  		JHisto_vs_Eff_Radius:JHisto_Bin_Boundaries = 0., 2., 4., 6., 8., 10., 15., 20., 30., 40., 50., 100., 150. ;
  		JHisto_vs_Eff_Radius:JHisto_Bin_Boundaries_Joint_Parameter = 4., 6., 8., 10., 12.5, 15., 17.5, 20., 25., 30. ;
  	int Histogram_Counts(longitude, latitude, vardim5) ;
  		Histogram_Counts:FillValue = -9999 ;
  		Histogram_Counts:Histogram_Bin_Boundaries = 0., 1., 2., 3., 4., 5., 6., 7., 8., 9., 10., 11., 12., 13., 14., 15., 16., 17., 18., 19., 20., 21., 22., 23., 24., 25., 26., 27., 28., 29., 30., 32., 34., 36., 38., 40., 42., 44., 46., 48., 50., 60., 70., 80., 90., 100., 150. ;
  	double Mean(longitude, latitude) ;
  		Mean:FillValue = -9999. ;
  		Mean:long_name = "Cloud Optical Thickness for Liquid Water Clouds (Primary Retrieval for Cloudy Scenes)" ;
  		Mean:units = "none" ;
  	int Pixel_Counts(longitude, latitude) ;
  		Pixel_Counts:FillValue = -9999 ;
  	double Standard_Deviation(longitude, latitude) ;
  		Standard_Deviation:FillValue = -9999. ;
  		Standard_Deviation:long_name = "Cloud Optical Thickness for Liquid Water Clouds (Primary Retrieval for Cloudy Scenes)" ;
  		Standard_Deviation:units = "none" ;

  // group attributes:
  		:long_name = "Cloud Optical Thickness for Liquid Water Clouds (Primary Retrieval for Cloudy Scenes)" ;
  		:units = "none" ;
  		:FillValue = -9999. ;
  		:valid_min = 0. ;
  		:valid_max = 150. ;
  		:scale_factor = 1. ;
  		:add_offset = 0. ;
  data:
  } // group Cloud_Optical_Thickness_Liquid

group: Cloud_Optical_Thickness_Ice {
  variables:
  	int JHisto_vs_Eff_Radius(longitude, latitude, vardim3, vardim4) ;
  		JHisto_vs_Eff_Radius:FillValue = -9999 ;
  		JHisto_vs_Eff_Radius:JHisto_Bin_Boundaries = 0., 2., 4., 6., 8., 10., 15., 20., 30., 40., 50., 100., 150. ;
  		JHisto_vs_Eff_Radius:JHisto_Bin_Boundaries_Joint_Parameter = 4., 6., 8., 10., 12.5, 15., 17.5, 20., 25., 30. ;

  // group attributes:
  		:long_name = "Cloud Optical Thickness for Ice Clouds (Primary Retrieval for Cloudy Scenes)" ;
  		:units = "none" ;
  		:FillValue = -9999. ;
  		:valid_min = 0. ;
  		:valid_max = 150. ;
  		:scale_factor = 1. ;
  		:add_offset = 0. ;
  data:
  } // group Cloud_Optical_Thickness_Ice
}
