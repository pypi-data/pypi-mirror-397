`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
dYVY1GBMsK1ODCn3ZUp8SoAWP8Fvt20jOclKciHf7Ysn2OlvHpNHbXI7BFbSBeZ8
c0HSNxtSIQSCmTTcVbiOe5bNYdnShY74EmVDlUagwaODhK9Urx30VHPfg7K0Q8Dj
u4EuL8LzGtWyNpPuuYUPfH/EWWJz8j2B3GlAugKl7fR1RciktYEXyNArDzj2i2Lo
icoQhkynNgC7v9DkMLR1BxAwtrFrckccZalCrbzlnjwD/DOLPtfjLaczesJPkKoa
xZJUnnMJHmZHdGCWDxS1eicDF7kXXzsE1BA2jAX7HQtg/mw+vmEQXKqvkKy9tRtW
yhUEHOXSIVFkC6gJ+buK9Q==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="SgR4h9hEc61j3UcDg7JP89NUc7gPf41F4aolx7zbZ/Y="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
PcTZf+e633x3tw5Pd+98Hvg8K8pEx1TP/UFyHup9OvIvZyp7VdJ/eQ7Czw0TCb/d
NGL0fQmqipTyP1VBR/CwCDPv8pUq9mWdoIhPzGBVMq1ZfAiLygNMWUwFu0/xPfyw
rAKvJfKF1tLDCsja4oREz1+w00FDmJ2gsQcbY/9d4Lw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="fB5pBzxyhRsqq3gFtq6qZ5Drx26WwP+GzJuJsgJq2oo="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 118752 )
`protect data_block
Pw0LuTSwA3gmWF21w7rVYBcj97hqvAcf4dxm1w8M8xOO9V5Zp53fD6281Uk66by2
V+2le3pjRQ4JkfVvu0vvltrqFdWvBln4SM9xPIyOvOgxR9dZ/mACNvSM4sNQA0B/
KMPlNGmabCnuPJDdj1MYqtQkNLpYyq06umUo9jVdvvnJOy67/Gjhoik3+mSGV8C5
qW4FQ314v4HwNtq8aZfcwC3wJzDc3Bzdt0tsBDNHZZTVaEuEyJEp1uVL/OLbkQ5E
Kn83gfApEDtwzYgEaGaSC6eNheLzx6v/8Vj1gMY3q/15+EJ0dZnUP2Zolo94SmBG
fsv0kf4b6yWk2DRIWGmieedicCQOTBuA1oJII06PKCjgJd4RSH33ii5qZoG6Xe+e
u9x+hgbPSsmH/LGAZteqHkfwEIeZ+Y6RUO1F2B5Mo9PeSCvLgNpAmJDGbYsI0y1G
Ueqyo65iNoA/d+LwnZiG4CMFvgNusfefFan1denzPdbdv3VIN5WZhLcF5iEMgJwY
47ZjmFYa3a0G30geTV7HqerxqIbjwjqysTWERMO6JxhiBo05R4Ya9Dvj0IAc66gr
zxGbQaViRkxabKiafhjPIo4J/Acqi2Fh9oG9iHB7ESuctAmUtiHMjnLFSjDbSyDP
Zzynr0XYwZUwBnxz11AKtz32/eI00yS3V4Ln3h4on+3V1WjQ4MLrVnX6sYJI1h9u
6HhabSBgjKhrKLN+nSC+DJ6qPkZJhHiyj6nPFCAtUSDigejcgAYD+Nubj78PPgqN
Bi33obRsmTMk5umEtzlfKxvHt3yt3zbLkiToQ0qo2ZYUaEIeoOmxFgabbVDOmogk
5FbgSj7+iK5yDeJo0c8BRV68H+TBO5iM0Zv2OfIqdOdFepKepqumGT7HIdXvji9i
cKia9kijITaoyHtOQzHXC+7ZL6HIu7IOougeFGzUE03/UJuVUBMv5d3rMNh7hwOa
AvHwmUnm0FiI7W19eZCQ8MVZXDBQY5BCBpxAa/Vh2FMZcce4NKCoL5aJ96GuS6pW
jS1ZqxF65OHW8S9DrH0kl318fJ1baU9UbU0Zrtq4gJNjYaqcz+rvak80b37N5piM
rvGGrWQaYkzOEE9VvHba+n/nlmn7XbeKOy9v3nqtP/RnlpO94HzCYFAXGVhDtZxe
xDXtGvKuavB1mecYMs1Yv43oM/Ht8WQbrBf2nUSdOu/GZFy8D0BOnCaIffvxN0VM
uWVYuBDnirzfJc02bkVcHQBg+8/jrZNNMEOXpRUL+wwT8iG9pwCeio2Yy5Pj1UeT
Bkln0Ujau0DAkrzsEnrtLTzIHjpNhaN2VAgfoG632PXCEYJ6J+pKu1Opy3x2gqWI
dLjuUpLIkl/U+O5lnTvo25GyeMzxGnwWkwMUNKVOiSPib3wb8ihNI6UTFHVw3TDe
pdDYvYoO8jOCSc0QUtx38HMaBSjlzCDLGxRtiFZ4wCYga53eZIhksKN27IGTjume
rpjV92rK44Mr+Vw/tzb+6EMUOWJxXOBfo57/i1LycOSxb1l9Ec/KBvTvnPgMLrrU
7yfLsBW6XgkYNjxTuaDfwLZvFEpvpkPZ4Y35uFWRc8EHScgAqx/eXRkte3zaQzt8
NX9n7DQsyv2l0M8PUnj/xQpYqS0FOQigX0lsPIvEcKpysZ4umd6SD4fD0S1vXSXt
famIGsMqbsNAQM9/n1uORCv+ie3Yy5NVxBk+pY+S8JVaFRYRXhaiw603TRB+K7J/
ud0jQzShTp+HZvIL9iV6mWW3LGucKKRfHd6bDlkI49mL8cX6QtncFB1A9T8peBqO
F44qAVWPZ3O2ZVYcZdFEoszo/3grbTVePYeMz/jDbYTIW7ctlwkWgHCPS59u8N+u
LY552nayRzHKBgzihgqQOgnkBwamtzbByYfArTU+FSWTrJqyXvKZXWpmsKlYtZ47
9UQCwag2s8ORSWL3HWfnwaulj1LuKcEkZ6ba25/s9dFBO5tyUN0MtJavqTRhBieG
qCUMeUDOLgVtQD5+wuDMQyX5WHoxORg1IcgLxrBxd/0EgKx+TtLmKmBcUHEfuwP3
9o8hjSFFL77UB0od64gJIU8+rpen2kfk5mPida/IBpxNf+Y37ExSYYpngFouNKuj
s3zO7pC8Ta3c/X2uTuS0p9VqP/7/NV9a0lXjv/DPVnlqvHzupcxveG2+qdx/qqkP
adPeeYDamn+QbzEZLM8Ol2f/zDsXEPi9O6xBVB0zYSUi5d67Gf1f0FkH3G9S8Ool
4xRB/V8LoOstur08a1ZybwjQ7lAxdsImeeMS4X/tv6m2vb6kwv3m5Gyh2kwkJwlD
c205ts2YZvOiPHuE372DWz63nqy3Jivdfw1wErd/fKUFkklyBlFJ8SkjlMKimX5c
VFUJpciXuoGxPKN/K3d6njKJFssk2BoSF0nA+zSp5GIPcEP86bREQAZWqv/T+Af2
BYZkXyFN4trrHzOBMGzqzUnsLNQ6FjWL1+q5aSFEYK8/Ec3UNPEmWaxUWBl5CFfV
9DhyfGdncOG3/pOKiotoJArX0Dd/S7xNHjg4LA66MrJm57jWIpuTa1EImEeO02Ig
+nBYQRgRlDQuLXInLzAu3aEUvplqOoP/qTmqSahOqOIzHB3vnD5ybi9RWuEeVWj0
mHnvFPcTE044BiBE186BAvg/0YoiC+QxQFrSy5TZ/myh7Luktk0eITxs8Sn2Nc1V
SqCOxnV2VBTkQeD+k0eswITVVobJcd/LW6iV8dhzKIdPGoaWKB33+s5zNYO1uL+3
Bq96P8sM3trOoPD8dWtBI1Rjp5BrHypMkD7md7slSYO+n/pxMTeGavary57V/8M2
HwUoVxclQMe5I94RMN8AjYp1bSUoBWkuMzRgOV46am+P9BqKfjyfLbJloxjXEtbe
6zwXhSLJ63mS3iQLUWysyjUP6fpdvxGWACXSluI5u9F2akPPsw7RiN+yCoyix3EK
C7uqXdoL60aHTRe4vYXJvlMYm72QAoNcyeCJFqdPMlZacZ2cQi262wGBc5u6gud1
CICaC09ui3J5O1kZACM9NPq60kmo0lxfi3c9BOzRTXASNXs8OeDOt5YqGgiZeHqa
8zvkDD3BO2zWe0J1nkpcQkNVlP4TtMy0MdHXemvQSB1SVNdyEOq/riqYQSizCwYp
jRMZ+scozbkO6CMG7fidEq9bitd6FqXXEU9PAAxob6hWrPlY73vWAmrlWUVY/1m0
1/YzubKLv9rdR4+YqMfW840edlNiwHM3p7EcxXy7QlZkbK32IHwAbKY/rUQkUuL0
yar7zOEQU8Z7i58JQD10cw0F9xgUZ+eZZJ3K6CDdeuA956Lfmu1qGG3rF9eZyU11
FeMHsvIbLICc5M48R7Bcd5PlV6thy711xzaaDA/+iSwyGNKlIuPOZxUUsR01hS7H
7wrty1uni44VKvY/rZjL2Opi5+xtAVc0kjVBbDtkrNHkeue0imv09p69XTOMBX4i
OJCCQrmX2cht4W8JRLj+zkfvcnCQt58edtCLGQnvpJxF1DgDGZnyXqdniSFj5MQ3
q94WDA15JAC32Kh+xYI7qtg0lDNth17PfxJzzG+hulLbvDgtggRqgQ8VDCYVIof0
q2+0OldCClelx+DT2JOyEuT1jvU+wfUReeMK4HLv3oiCxSWuawwdJWNP+IDCTFAa
mtkQ6YfISpZFj0+Bm7ZbMrRqpiQTwyIy0Cy2gtA8fJ3HKoorSVlKBmeVi1wNYmhI
Q9z9DRzzCioAHZ076P8ebgWexC87fi2JV54bOjJHsIVoxzOXRpb6/0FsbJMCAjiU
04KNwDDb/t9kJYmSUxMofb6axJ2z5Xghjp3quJZS7S0cv2lfSjIft1IPsEq65V0F
xwyPxK0ZtmizzFZ31N9iafaOCoD/OV6qQY+9zz4gqJNX8mwDRSQ7JJ+yGoKiP8Wu
SR2+EYGFqcZNi0IJHRJEIBRWHjSjzy0N24X0QwK7um2RtYW2EMNKkW0WKInvf1i/
T2niqwBu6v/RzbPBAOYDA0EXi146N8U9z8uk7iLpqbhzCbPC/jtmP3TjQlo5q1gq
2TH+eA2f9up+9Dg821Kd7NbmERuylzUK1eyv/itO4dp3aZpWiSWOMESgO7fp7nfd
HnkFsnmMuUiPDyfeqyVXmneNRsYQOn5asm55Eb+7VZuadB34iAxOWV8BHgPHnqWT
RAaToO45Ng5moJ6FXEZI2IjAB4uBclk3nBCJiO3knVfNSHqv3Wfx28QIgqp7NJS2
W7LDHgHMItsQVUuub4JaHMeenKLg31Am+iHav2XoEYK9YDdmywx0OTKEn8dgdTZ4
cvC/wwOv1NQXnA5WEHeVVWkxd2HEFUTc70d5JCr9yd+ot4MZpi1Bm5DUF2R4iCJW
gunULhq9/RIrQLcpI7Y0ftgyvNF7kzwSDJ+c1kM3T9ai8ak/hKU8ls/HoXL7sVJn
hAhuluP+HjFmDhPHLD6gbc3v6BF8b0hfy60kY4rwwNgwFD/NR2nFNKBSWC0qeBSx
HjXr2BKptqYnUGA+5OkmsIwI71EArLFAZvpcGQvIikTwF1Z5MoXZPbpZ3ERlyf9F
gyF7YKAysCeZYt80R2WWhzXScmEu4aAixx0shsns2oZVw3RL5q259OYMydweG1D1
jP/wpkuDmQq2OkAoudmvItQXAoT07vUbKLmUxUYcJApeESHrJU7PZRyITbBEEdt9
rGyplF8Qv6DCqzKbH9Ij1SWBQXLYzOkD1NgG4gI14gjOZTpmWOScOvQnQsxv6abl
ZrN/1nBV96PYPfEbpKnt5CU/zqJHVsQaClQyaKwTmEit8iRb7apFlmeaeVoejxxw
ra/M/G3XbebswJtJVMKawRIOSukL1PHa0wpldNb+tlDwyZWsCV/RXmRzL9fHgymD
bmH74syEOSCYMZfGVweKhwzw2n3ERGYhKnOJnJqNTc0FgBHu10hw07VSAnqmEmGd
RDir658MBNXVpPJm4nYIbEwJgqxK9dEv1AhaWN1vgvzhOY6HAQIS8rokhOJpEtSD
a0xZyLuaZvmlz6w0ZWQulw39rpDTznzBmGZzhazxTckbjRTXXXxpNIEyJUUMh7yt
/yeekIrO6EI2tWt4E7AnNazuwI/mC2Dz6HjHE8AWyFyiuOiDeLS0xMGV5j9/v/Jy
opfdJr5Z6RcU7k/ArUOD713dSu4KBBvmTBLuZMXdgQsLd1uyLshDXamzsCJc4u7V
2/NSMU50Yn294hxJFSKFYc68VOdLHy263f6b/tapLu0UhZ59jL1+roik8sRKPfnP
mHLlOfQTC/J929u9hJM1Q1XLM8IZdngRnb0apxlaKCkEN+52+rG6yKFlfm7R48fz
2t9l/ghGhJ2vPdhuttrUa/Jh/+pc4HC8Qp/XdSweWaHBRQFwC+7ntxnogp8M3A7/
QKcaF3uBPrLbbJQ1vgvYK2QhBKBRDDkkRFeiHPBrkqluEo5m3OJxAJr2Ao5+6F14
nhvrA5ugn4kIcflOIe6G4h6Asmx9LOmfjd+DeS2jLWMXq3dXhWRe4Wu8BltCh9RO
Rr0GlQh/fGPeOASemxK2DJeUGHOcSYiWIw+I+N5OSHjThxwHWSPaZ3gcfqPQgAYC
jMncZaY4BVUFhcoOFvdLKlO6c+hZTObkz3c0zxf5hhum/j/42XQ4EuK3YAQUxp+o
BucW7QJN560ihKl2aJiEte7ApeSzuvj2qtLq9wprOq1tLneuXUiYGjNReBISas7V
7a/sQffYeUsoakKvm1ScUY154s53co4c6fzabyHgGbmDiAW1rV0ag94rn/8vxCcm
VKsZm6OEqsDzyiazFMbqweOTxMybtPEyFHF3HKGUZ/6KT9rkZqvXPhVAjNPlTM2u
+wBweEmvfr0aF8ZTOuqml5zNAibrFOhYA0YOt0RW3AMP8ma4If2d8o1yoJlq0Xjg
iqWtkyLBb892xoqGV00/sakJTLAzb4OrSCNxt5f77B96FtF7EcvwF0HLqQpwRNVE
MMR7GINgNgCeZ7EJA4pjIhlzvgZipDq6lsHVtDmsUV5PRoE8a5lChc6HabqOZCb+
USVRFb7Enn+8MJt1HBeBtoRjsuysFPEI0j/R4td3SuDt07Tr6iN0UxkacLyHN8jC
B5mx9W8zPQr0qC6fMo1VjbFm0UlSYjKC9AWXYjeX3EYnAsnhYid4OoKUBjWJ3GdW
vXEUNlyckmkkyW2SBKhgXWUeXUx4s0spxkISXIdDIWLPol0Dyn9Y3a3pABq8A7SG
SJtMhd8fhridou1nj2HZxx/XpKtY5N5lzXbEZ06J+lfxnAPbH/+wWpRyUofZ+Hz3
OtMFHh/14gSjy7C9ZUAXmrKAjR1qte+khCByZ8bDEX/9lKzhRy6TlCtWiGOsr6ev
HnC4sGubKEnZ5XZL99pTBviRRt/+P/caiJoR0FATrkECl1GVOp48vnlMFZlZMOUW
uk/iY78gP4cFF1hLP072kthFXTtSVhoo/1KqSLUBvNY+F+CnjwvaZsWTA7FCLz8u
JZJGfJiRSWpBan7RWtXd3ZNdzSYzEqVeLkWoyVMKI4eyo7etKMLTa5X5Y+lg6HYu
45Xs2hUqmAM/6YbdI5hXx+pGlqpMfJBnfm89ha5B5i1L5zL9KMr5o4bxJ/1nw3Aw
4BBIDnKA8xxL9h9qe054i9Pm/Pt/fwcI8P9rt0ucKSRjaSU/xmfqvlsc2F6Stbs1
MJjidhh4+LcGh46crHIUItbFzyDnild26NVYc+GslqweV48A2vSi/RbkSGzmwrak
/93xK4Yz5bStgGXKQqcif0sSKXzV+lgeaziH3mL4ExGos3s9FVVV9ENwb7zHyfES
rBScnefrNDksPmufHgqd4VEzT3fxnTB4vXMooBOR0UwdDGzmyLZuwRmllZ/KDIYV
0NfF1ykOdCv42UQyf4CUlz0fdzUp5sZREyPE+tk7S8LQWRsCH8veil2iVrZcMaUa
98+LHnsq4Jt0JBXfLycv80OTyPTwSImwb1VELUueD4+I+JYqcOtG3C8kO4hxSX+V
IeI+iHlK9c0rqZiPJXbusdpYKLvp0KKNHXhyY9rCidJjIQNSIsaEq3Epb4lhXjTp
L9DGu2IC+FIFFzVp4XYwpgyp6beihp5vtsyrHoruR1DKOiev3oMIJhz/oBVSTgle
CZSDBOgm08IOGi9eco2tGuwgB+tkM4SVTZa3y9w1o9af9QoATD5TL9LQEetngQPu
hZeeZLsAHuc+mW5pRWzB88jzrlRqTBT6klwL1zkgWH1THtXoxH+/sPykR0Bm+YKH
arb6pGguwiJr6S96Ser867g5Prx9LH+Iuw9CwStV7r8pr4mVQGfrhvBg7e7mgJcZ
aEFnsv7PDWVPsiaYBQLDZxIGtMuBEC+BwRoWz2rkLCZYH71ToLHKIoPsQeF34fYt
7G/YnlQ1w3o9nXHE7GV6nXnc0Qp70Cu/ww8cSxB7vs7/BJQx+5b4KRlgUDbTvEwk
NB6w+HXmSstGrDy9H+7wu3XzfTnybTMiOnu7ctwLRrX6+Mrm34ySxf9vGO4VW4iW
ArCib4qX8QTDhcK0uEK1FtiGQfqRoeLZlDC8TqEBnouSVE8cedxH57aKMDeUgchu
V0MNB6KIAj8gUPYKKQ3E5n1m1VM0KUirLD+1jqiLvaL58hNJiRWk3yHXsp3LUOzP
pBbm1V39DCSUFl/gE5hZbsvfAxLovwAdXmPLz99abXaUrVFI/rai928ExIFiO0Fb
q+SDzGLaGGjmYkkg9aeIup/l7tkYqGKB2pgbriOpZkTrXCyRe7KO18WnuCn7wRi7
yc8iPad7OrsCHaOXFYVRNZjFSk87NlEYAmZBcFZmURayCMirkS2ElrKniHAa7jvG
yXEoFcpXbErm8ZoZpRjy3mHyiFLnRppaZpdwuvvshEgsbS9z8k5unonNhOpWA9+Y
kQ4i2a/gbRifdQ42t3Owi9zVEh2CgLqpihwgLWEiUbg82HhXWeSa/2M/PkG0EbaN
K4nvfzwxxjSJKXPXYn+xfITMQIhtzYeIQVdr9XOv8U3sGG4UJNd2nyE8cnfgpKyG
cBn6YsWHEe0Lovc3sDhWNVzwY87xK7sc2GtRRlMPaSpfryOpwob15oMkz0Nw55Xn
rrEG+IV0Uwfe+hG/bxl7hKf5N/VmolQrreiQfNrYXpk+3q+hNOJ+DBD7VwHqVZNY
zVJf5TrXDCy6Qv81EGv2btag9Gku/nTD9Bs9zioJoElAJapOpAB4+MGhyx+w6K4J
NGa4W6GXw9UsbXGItmPS+a+iyllL3dR9dRFkzErpO7aG6zbcHP7f3DWWZWKpAIIT
jfgsCOan292gQa6WR0LnF8WzZ09QjcHyAZZzM7/3lFJ8lWj7AomIWYI7LWGlM0kt
uG+l8J8Q83234koSQ0kuHzcBIaNpq9PZjDPTIvrd+8yQzkPKhEyyPHbl8CdMEcrP
pvNBN7Xw8B+BKI5W6gLwWala1/XiCLTY3XTFsOecJ5EvRtpVmNSfAu+Mvkzwqgra
ehDIY7Q/DtUIrAcCbKjeQZw4tiQeW63mrqgIx9/O/mwUmDc/PttaiJW6CC+TVeWS
tKezcY4ZGeT2jJ47hVl9zzPxUSBmMBq79AEHw2AYDj3v8g3oLmMaaOy7ksON+SIR
WM9PdFCQH5DHbw17dd/TznvWYJ/2yswHKoDgN5CfwsKxcLo4TQYJdbsKZQc9fSCD
n06I/BaZSyAx+6mNgUieQIhlUCIXdAYT0wSRZtT6bQWFRis5OKzj8Yu8d3AdUYBv
3caCDOv9IH+5UoKAWk/uu+xw4uU8iIpl3uNyTvbY72lTZSWUg3Kjw83fCA4RSrIg
nO2vnF+HfOfdPJYJPwDr2J/XIgE1S4y7krNIIOY0oASJPTCm+AAmG+M/6+wICOrm
rVKmt1t2mHLZIrlwNaPdGwKZmrPyK0Bc+P+pTexqeCi+pw7VbC/2NvL1+JhE+Kib
kUx8OYfdhr/ggD386SwhWAdKCGCgmxDAZM05ktqi7U3k70aO1VVy3vpMu8d6l7sf
y28Oe6eXgHgJNBnXxjRoP8LlVCoxUYOx+g2nLVLi7fEPeRl2h7HrIWO8u/maVgsx
J7MOotaDuZi/ySLZyoQN/5oaRkJLGutTXBiYS2nuTvyoXzwi0A2Qu/FeflA4h9W/
Ts6lrUp6mRRaLbdie5GGb2C6uJg0OJymnaALfMz7NLl5AcI9150Xq+TO7FLKxxqY
bno57tms/1zZCKiFbWmZ9esAoyPtlf9SM0HgXeZSTicHz2qQw0274gN6p177SQ32
+BYMNRttzugq4re2pDcSSvrbJO6jnzYn1gfA+FEsmGonwMlp/gbCBLTOHXYq80r8
+J1ViXIqWvwHfGGIDGdPUv8Ox67sw4DJJF7Ke33Kt6kW2uahLy/5iBbDGZDcBonG
Zk/OiNbLxJVPfTMLzWSkeYwxP/yw1OI9DrikLlxYm94YyguahFTx7eQqpwgKZR0g
5EYUG1Cj+C+vCpXn0wEtvwphamEJTx5AIaO2ogLVdvLLoKnDriboKJOVJQi+TYMX
m832UJO86jUXw7UpKgiEtDak7Nx1gVXqkWCu8sHhBAL+y32bC8q1XTJx2SWji4v/
OttQoafDF76tphfy9q4ZrwCFAjOn5tr1/lQCksQcWiJSqvSujpQGmeAF+MMYNKtE
MBqW4wcOY127e83d010QW6qlUA5mKkzAdhswf4cdqfmkTI0pQrUBqb8DH8W+vAAv
n3cgkmXMHpnCQ+8JR7jinqA7PzgNRKh1AWJG45AkGAdADc/lbk6PlKj45jJTMxSV
mBHZ82NblSTnfEoT1hjTcqYWnc11bAWmn5ZHEF1+WPGIeGkg+MTo4+nmIBMofbif
BVjDjAykxa+Jn/bNyuiQMK+wAhAfucQa4joL9PQbAM6B9ibUtg5PcpEAmDmAXo8d
yLMnzNLjSrasy4gQ3BVoDW8B6QE1+On05Zej3Da4aaC0hY7wLmXtz2z5R33VeZZ8
fLOw9LXdjRGi3FF5n0Sm0U0A+64rjQ0sserUrLayS8z24neULztU1r+osoKIT6YN
pQ50qHKVydd/kDea70AMM4Jt0FlqsAAOazPOkqU9MNLJ6xNLjMEiOSU3hB34/owx
rFp4iV7lSvP4MkxP7nv4jLuPgSxJs/a1Y8e/dZXy5Q2pB6Fx3PvD2PwfxrwZYX2M
u2pgMJ6/rq0OxHM+/cZZCS2NijevZb4cP3aMHCtgjT7eNhihllxWPHQvdJcOl+h0
1znCNxJi6XHbrwIcVtJq3DgOxYYhMiadAcgWa10FPjuBd7G8ZPYd1YaNawPRXXkl
jniZlgra7fPnZw9n0wCui2q/iUGlYf89si82KyKFosxH5l1YmJxdtKdyfrPp+eri
bZcxKksyoAQFzdWYeZoHwsWX7lxhRWU/JAgxJqykRiZHrLLN78G/wRdBSg2WZeC1
EDG+u4Gfp2HHDHNDvQDww67BGrOvUtEclnuu2pj0dz562voOnMpyrUJz8WMeEhnm
c8RUxkMC22YHYEB5uLphnZHaKLXSKFlByetuJ5MqfqXDVmcC0m6LyUiA3fbmubrc
xiWnexRafV41X8IA2RJCr176joa/qrrdZ9/Jl/YhoCJr05Do5Yttu85x7NuubF7x
ksDId5pjO+ZuIJRLr0DO4uS7zdLsBHDnHE1EpD5QJEMw0/2gddOEunrH64BHWFpy
GjEGem6aeaj4iTJEozr9GLPxkUKqd6CGYMXtc2YjGJG+dTsTbJQeCoCoB8UeaiII
b8xFNJbiYZyR/RtrdhU0/IKvin0tgs3KufTghx7kKo0X6cKvy0J+ZWwife0DyT4d
g9HZq5uEhEPDC0hUCIAvdUjWhp2qt3f8nqmdee5cOq446pwz0v1aOz1oZ+Uz3Aaq
obit3sw14G5tN4yXouN8IuSnVZP1auP7j7ijtvCiHrRFCSDrsGEVUyfOFQcl8on4
NMyDe/bKhfI20CPk+dQk0BsNwh/tIEgSauiQluM+Xvl6KysnUW/Z+fc+FYSlF57K
jnnKu+QYoDXxWyFUFA48ep8EhCpdkbegMo80wS87DYq+zlxzo1Ga0hRUtk18MMNz
HuMOk9GPYnhiA+ErlCe6zaVeKIyotHs9aWnBuwdptWSE5rDcADYCi5OW49tVflbO
VsCru1S5xjZ24QE/vM7gx+rXfe3UmOsa7h7nnNOkeuf704CkN/E+EuWK97Nb0iIn
uLgSLihV3ehmx11G7B/0KWV6qWvy0AjcVuReCzN/UustS9q+Yz8EWv6OxeDtenbm
e8wCaDbSREVKiytLItcgXnjuOGQ7LmDY9ZCZTOLyvTBIKKVVbgJNxWRyLJ/llLPX
9AZxmVmpmX+ApTc3IgxbKaaN9p7g1p0KCFsyom6zYT6Yc7CtFD34wkxYFd6B1VAW
kXiLHUFC0N3DXGnMtcY2NZhzCbi7YdnqCFemH6W437UHvCgm4u7vDok0iAr6jlfc
KsHn05VdC+i67LEYKzdD7zKuOZUP0gNM9GTUxbocE1BEl3rAUNJohIQKxrTg93al
OvYWARNn17UpBX+WxfQdYFQ/VqwfqtHYdZ3WGb0DgH2SIp1j1FAlQiHmyxF4kl3J
vVD0/btHi5MPtYTppcR2rxRFuKC55EyZOKcDOr5yBDL6r24DFSSss2/V1vvt6Mjh
XypL7hfLYLv9f9X7aOreXe2Z3HLyjdGLrOmC5Haf813RZesP6q6n7O8L6foYo+N5
9GjqxG/ekt8g9R5Q6cFkoP5LND0j1tGJYrzaMdpn704ZxjLKNs7Qp3p1RMEYf3nw
To9gCq9NZKehtkY+iKHW/tdnN1odhtU7TuLalqJJJe1+TEQuXWK4sLfhQ+XMS7ex
u73LEF73JuBwbxfzEbT16YonC+SaXOUXtmZnihM1h0GH8tBS624vYn8xE74LYLE0
Zziso01aJCuhJDQn/R35bMSPMyBYmg0fg0PBeRLvajyZNWyweuwKir4T58zIsrYp
o9auQ60TQv+O5j7VdnbGYDc5yfNGifGLFaB7XHoPDHLr1Es5k2J6JAM00Gc4zKts
8CykWyw/YlBwT6VnGyYsbtYH04NwOHF7OvKrNJ+CoJCQkUN5lp7OldqQfUYHya/e
m2wzcdloDA4VTfloYxd/qECNDjPlXZyk3wiNuCB4hvmyBENfQthKl1fAFhCH5Djg
y5g/Z/x6v/S/RP4GqSkqq79CuW4FDER5zUDHKyRDl9GsQl2BCB+Yo5ZoAN2oITZ6
uY47AxWSkQlA0a6qL/vKEBAqNj6KJnZ88vJxrnAhc5nQSKVDcCH895GnMnquIYTY
s7UDGHb/9b+9BzpxVGyEwPNweoCMaV3qSZWebx85WyI/367v6d3GHeuTtk44uJ9W
/mQY9UsIuN8wjdz048CCt0/ZwFwQZ00TPytVnaEbKweigqNJUaNzde/y1XmZGR+l
LwpqhEkYOPT3TuGK+SVMf8Txd0s1xzTaoNnFKDeZtWNt6BMWLtGLT787lpFM4ztK
8yAuyi5lkb9w6mVPcoDMVVMSbS5SFVsLdu8aJFj7s5PDLZxKTPm6h9Vwp20TG9oe
1kWGpJAHtS3MHLg4EmoL6EglpZGKKuN+xO79kPVbJmHvmPOhRWFCUYFrcCV97RCT
XndquUeUA2ReLQD/0KMcvTGKUJ0r0C7gFyGvuhm7M30El3wr+bDpH8rvHE2Gt6cO
CHIhGL1RAOsP7yjAcb3AZghUxSlhLp/+Dd+fpaToVI2YYCwXMcbXIp06VV2qp17l
LEWOnGsSB01QoA0iECe0XWMxASU/8yNlRBfrAZfKwOorvKpGhXr1QTjg8dA4YztA
VxJ6zrXzlYk4jfaehm4GJ0Rszs0p3svS4IIGJRW7QYBsG4RsAKZLH2cDGf7sX/9p
6PgNTssYa3ihGctjBZDI1/qOWXzb8JfiTq1rnvq4cLKbbRj4aet82GypDZhcPDw6
9fhXc+eNec8xOwMnH3JbOIwrHIPLXmDdAaHTDdv9CR5wUzUSHtwB87/W7Pc67xia
zTYa/KPQ1gCHaqotbN+w9fuNV1xqt8FGu8Gc1sQFzvH8udi07k+HKt6iL+errOJI
SrChMEo2FzuAwzkC44Mzb2dAFPFV2kLPuoiDUmKJSk6dmoiod3TGQtVlo0sYiG8L
mVTYcEiN/EH8bd63xTpHv2pF3RmqHgMfmwy66VNNSFjcEzOE1JZsWRUxSvf/Nkse
wFrzKYuKqPpUntulsw6Zln7N+am57iCoR14KjqMevSB1k3jQhDblgmD5S7B1jLBF
Dq3EIyx5FGPW3KznxnCGPwTM6CYxjSpLLqRXY5wGl4maYs+O96PW9ZqLthO2jXXM
FSVE49BoeXEFSFJwbfAclIJHSEmIzxcNueAKaip7iWKlkwJw1Yu4qj0XXjm3WOz/
jJPXo+7ZcEIgvhmi160AqdEabGrKUOD6dMAZ2U9nv8u1HnsD5IOOXH8cfV7ZlTkt
gTvkF2yQiYKBn7n2WIQ0LV2kDu4e4S7gD+Z/zhOWGXaQqlm0eBKY2S1UNTFH7Wf8
dYeT61uqmjcua/Bw8hOhMqsNC0H3ZOqn7xlpUZ3dyAFYM2KWPl/DWmDnrMG1vYtV
vIdXf2W8GWB6HI0RSuaQ/LlvrTDlh3FxS5AAnyeeH3SqCuXTPoShREUQxuDVR96w
KQsaXb31iiMjW0UckOlT34ssQ57kEqzpXRqqWMe20ZjO9akYv/zHmlElMPTzRxvI
Hs33B4jgQTVXUAy82fjQmDkiXK8OrfF1pkrCkzGrPH71ExKqNN8MtUt9kONiDrCx
FEtL1xpBViq0MNxixV+aEADnGY9A7wyecjjMzoVRArWUH53smPS7r9HRs7Oo179x
UmhNXjqNOETE14sScYktiU1YFHjqfyhKQRqAVJF0CedK92XWW0UaADYCgaQwRh4S
OMNrfV0nUDdZrDMf6T7lccG5sytrcws3D1ojNZHnGDInNhB4KYTIZcG7uFFZc5Rv
Z8NHgok4Nn6mADRErIS6FNZhaqod801IPWvePEy8cnY8MTI/cBRaB5TDzhSluqLm
f7yfriNaTRcyybP695+z+6HDAyCARi3e6T9+dSA0OlRVgUpusgO6VrDTsuQh/ed/
KOj367kObOzG8Y0u1rfHP3YoBPDe1B4IS6cf79kafH6YvigcPrQOFAtqNa6JOK+O
A2EW3uMn0pQPmFRZDT5WVP8Py9H/cpHRyKI9jjQfQrVg00Bqi/ss+m9L6F3CiN2E
+z83b2RvrVnPd6/nkZDX4LhbcYA70DYGqibp8IXeRa7PDg2Zlf511S5QNbW2X228
zwrhtLQuGuxaMRZ76pwTDmm5RcbVpCeYNUUDAQtIMHgMLDH3Cd8aXUM1zPXYK/wm
EZOSt2QiWysflHhQVoNg3p5B4Ktr8rTV/HUoe0LKSLRm5rxZU6GLVAOTB0cKlwJ6
uD+TOux4VVDCsJmIyrKg4WqVA+48nbLFdjSYcFzfpMfrvMZBoT2aI4wTeBBbhkd8
cxNhyPLGTroResCHGNwyYQtoS+e9taB6Z8fHygmLsBbBnMmxK8TrAhbMlelC3LFm
Qsx/9bQ4QmZdUBOSlKDtaNL7rGJzLOamilG54THL0Boqob/yjiCdLLdcc+2H2jS/
/o0LjmLkNp9Cz4LN5W/M9hFB+mfT3ZbdR5FkkXTASdzyqsDhbIpGP+Hnf0XzxpvO
zuSlyNFT2/GBVmsWr/0UeQ5wq2xcQMq2e0fEBqfLwBzcA0ZV7vRS7Goygp0faC05
t2Bw0JlW4XnmSqFncMAzbpP2PtD8HxJZhc9UBtEffcIDsJ1hJZd/Cs0NCTMIS745
ZI5FUFwzlMFhvLgk5Lnw25Uzd8EWFPlAXTHRzNBOW5o6PmU2Z8M2d/lhg6i/Hq0L
LoXX7Fxndprbr3r+dl75Wsy7l45wn2qf/RtOdzD+jQtss6T4QM7Vm3LBfJ5tn7YN
8bEcE1f0ZQJ25O4+MekBnCyF64yX0Jc3N61Tje425tCdqlf6/Vy0YkcFYz6NLdO6
zAjJuvjxcpcbwBDkk+ZtUvrrZR4XKj2+oyQ1N2JbVueBKxxYxtFp3TMzER69AZd6
Pn7GP9tNxtifDOOk1oP0yr4CCZK9l/qx+9JZAFay9OE1Sw39Y4hF0vb8/Z4O6TbN
tqD1mz2U/zjMTnWIT5W68OQXxxbOsVKNSDNjHwJhTVL7QiaS3vF7iG4BqYn4gLjB
DoG26c6fr37AW5wy2Y758mso2IOmsLT1LnFZ4TOA4AOohQnMhriTG6BVVeHqyaMk
UGuWGU2E9XHnoswyQRH2kitrIeFC1dGAW864mwyEzMONR/82Q4kF0KsUd3+wCkkJ
5pGdwxR+8W7/L7RnEc50zMdguS0WfK+PjZZYrQnCxDDb7XTcHqQ7gujhYT7Gg6R/
DEWmsRI3iCGjGCG3Ky7OrpaznDh6i9BO5UfLxaPeVd+oISWlRTCayecvFSfloIUY
YFfa3CQo9GJh5MrTP78Z0CxX3vqDLfv3P6nK/WIvp4zyiR0WXH9ebuAvrsAwp/V6
hJEmwrsyjnRlDX9LgQDiXngpheeH8I6w6g33JDR3W6ujPV+I/XikGueqRMxJDTzB
8JM3IpAGqVY4N8Ee/TiYtcjWeZTVgDsS1KmuzsbGj7/qxp8hKHrnRb3D46erwvc6
q1bjhqCD38jM0O6zjSYoc/xAnKIyQ/dpW3U5mvc34VL/pUgMrOW43FbYxYjGipA2
FPtFgTnFVWtzK0q99zj7d11WS5/2hb+031v8G3cQVGc0BF8AS0DWB52v1T4pATF3
kiQXHOJ2bmtNQ4eW7xPrrdkZOfkTFCgIwp0oj1MuNEfkIRhZQfR8fGrj3Vgy+j8L
4+NM0zEmHppCTB2yhVo8h7tZEfU7PiFhG8Z0ta+9oy0Lbp0MxbGIMeHWDsahGJQ+
CoRWUwdwWszZpcR+ptGIcKtR0BqiF+OgXdooeHQVNJEwNpneFizXVmfr93gSrZQY
t80F+BUPON3qr6Ea0JjSVfxM6RSjubnpYXdsdBNf3RudpKAuINzdtPCZhoRGAC06
7FCumC8hC1fljarP04Ulon8pvlnYox64Obter2gYCqij9E3xNjc6q7rD6hMX/VQ2
5ZZWzpOQk9FHv1nT3LJsiiZ3FYU6s/QgT8BJYYt5NpBJ1zk2ihbG5VnKIg7C8AJ8
fvYiSx6sfB3gqThlp1I10+IdPb9orC9FehWjmBLUBPp475DEhVyrWTqdEE0ZAxil
ejffy5T7lxnTZ656u4LZ/xqhVA+fFU0S+0K5cqba7/knDpzGQODBJU2EQpmkAADV
YqwWpslwfKC648Tzgiv9E6vlRZFGfYSbN/MVZH4RaGE+yIm7ILrO/ywlfwLzjy+t
imGjalAOuZGmm/Jv3L+QTV+kfA2JEaUmGCnWPJ7c3PpD/ywb0plObdxVQzv8DC/F
UfHNIyuFihh9lZ/+6bcQAnSbT1jXoP9rcWouLmEQACnAZGyeyRlP+yNaR2oy6H5Z
hqx+89H1b3iOI2JINjgZACDuskikDo2/qPkggDvoqS4Pra/Jw4cXVoU2ZbdkyBkR
Ct28XPse2oxbrBtWRn16c9mQyzrAlSA3ybE95x/78MOuKQfP6ncb/iH4XSdPPZ85
HwXhFWR0eFcAPNUZGCmcW1B10Q28p3MPfAwhoJUUkeXNIAz5L1I/jXc2yEj1CIs0
Srww+0a7YqCwVHTqxRXNRmymTF3ZkfUBF2e8ROFrDya0YRnxbT+5SJjdeTdnK4tu
LqMaTYmLk5uV4Vt/+duVaW3QSUGzn07OUq7UIJAky/8s+i9XdpZty6bIThuoZd5p
p/0bAvlR6a7sjVFbDLIMjH/uNks8pK0DPArG2ZVH7KNqqdQYmPRS2aEdlc8v+Gri
rPQtEK9DzTo1Rag6cKS29ukeLLSuMeWyAyKctipe4BG7Fyc/2w5RDkU6Eq7xWF68
WTTVuQgqJlDulk/jniDYkhnr4EQiXQmhcS7oAtxg8tGXxpTwEOZCFB7/oEltsPhd
AjBs/awnTdlDo5mYzbghRmVs3OzOLPUA/qzaTB+M8mgvobZ8eKu2Apso4c8T705k
LuShJNJzhR8ePguZ3gZswfXcUSICBwVylx016umQ3BsDtoyd/9Xr43CENL7se56l
kM96YSo7Qp/2X4Ttn7iHsHj2+aoa0h6YiwUd+9YavsiapjJY1qdExDXLshcR1FmN
kd8uaOuUZgL9cRMrwAMGoDIhZz7A96vabm6Azz96X3ilmjg3E82fUCICWtsbmWrB
vVSuwE+NcY1bV6qJuMlYBT1cqmq/zcBToe+Wl29N4M00+L6U4W8ukWvB/Bi1SpzB
pFrQ+vziOmEojYrP2hdkhKoTaBZnVnsvgqe/kl0GnaZCRsgtLZQUuPIHBXR9EzuY
9qVrEakeDLF7IGJfBroeMy+VypWxQk8hFDZQHP6cJRb4K0pssvp6tPd9GzNdKwKC
TQlRymD2imCP5QvHHd6r+snEc1jmdjmf5ksT4nIJ5uTvjVJmwjn8A2aTflkc4wPA
tt/suCiVbzEHRW+BcqGZdqmBa5Oqr0guJAiCyO0Ppv8LBgfx4TZXw4s53kuKXP/l
qFpbtoW15wIMt2Zk4kMrGM5LoVd/G8km9WJZRiQ3Zv8oxavugDF4LbSBF1Wmm3nF
aMdV8WUlSASN/LL3eIN2KmmEScxU0HE5mRG8j71/yC+dA8t9ssQdMZDTSkNyn6W/
SoMhykgm3bdwJh/YKLenHXQRUttk3VyNcqL1TgIl2iPBBZ4808rEnckyXlDOf8hm
6aYdWcbEWLlKWDu45VDynbPtG0c5EyKrVMQ//xEFcg4aW6fHwVKfHH0fIASli/RZ
FZCLrWbUBo45ACu2ECzWzjV9mlthEWbP2i1stbFNeNBq50l0lwbumT0wSdcn5XZH
0ylxZ9gXatg8m+q/HNZqM4GTvRDcltGwnDDmAV7Ww1oBnoeJmpeB1eXYhM7SZJ61
Ju7k1C9Z7anBaFpIucanMLPTdCStL6iJ0fSQIk+882gnnfKyABPAJQCb3qf4XbTY
HpsMxANm5R2cUWFIFD8CJAazCZtu9hun5AgI9069/tkLssrenkcEsoUhtsgWjRsQ
WI3cvSoyR0jA6yOGtXQGAZc31Cvpd1X6rGtzEoTp5MTDhSinjxmzd1zc9HjNMy+S
acaZ4RWcX+jX7zSw1QxKQHmpIS6JGOWIAHqKtt7eIeszQtnQp9W0ePpRls/zfUqc
f8V5RsatiF5WM1NiJ09D2WleoYBViTyjvyN1bL9KGOIsZxl3vzWolxJEGVJV7Jnx
R2PgRZEghTNEmxQlfRKLip8OLgPlU7rTNW557vCMI9hVy9nU3+EWmPc4L278+q05
1s8ua0hL8pIpkogxfLsDS2jevx/luNOSCtVlX9jWsZNSamqsnh8d6jG5d2UMOcTo
uZ1wjJatgRYzVl2r18N+/mS6p3sCRXwgHAA7qiCWehpZfTASvt7n7uxHm2nQ74sm
XTbMznzgsAkstV3HrrpEWu5FCMv8X7jLJSbezbYeQSdpNbZqZkYnK0aVGxz7gPvD
ygvxQNqADKCxPJm5He4CoCxVx6HGgvzha6QRdBHyP3koGpoyUt0y36+JD6+LePBJ
0zJ7K36DxLnlg3nWcRTFAlieoZY987eyODH21hlcdc/L3Ih8opFrbuESXCs33wSS
wa9lhSLki/zFtJiRP6b9s02aLHFWXSSvXIkPezNpJxLqWiUemb2xXKE6Oafa4Lw2
24XHu1wzZTfGWqrAUhOuCc5n0huJT9hdAA48pDO+/q9YyoRMgCzA8ijBbFt7JTVj
PGe1wD+QkPn5tITrVQfqpNsbHMXfOMsCt6PaMOtnS6iMHX7stlIDSg9nK95wF8X6
hGbRGpB1pSToFVdX8pR4vBKKSwFZkUdpb2AIp98vcfKfPxO8X4c1yckbabUsCGxy
mCXSRK7mA5kkLJSXMn9CeJIc/Jk39Jzzp9r35UYensFp2Br1F7EH0eFKbFuk0hrS
ToiARJhpS9ZM6Jwcg10B3AcAy8CmfuTsq0UF9txXwmBFscYJOqgkaeOo/0uYprVK
DCz65F/pfMzwvrva2Yvr7+tTZDCSTo4sCu7NJ95YdtGKu4MmNjkzYQ96w0e0Sw47
1tmCScHKHpxJbVFzsIC6irP4O28WY0MlQYmmhAmikduvXwa3cXE1CYCNmp71i6pz
wzaZcGALHunNpWEOjizLKodnpbuh0CrftmLzSaRGfXt8RPEn219VT2TyCRcSjOXq
C7ebte3qRlBNe1DMO3bDjF4aStVkH/XBey2/NJQqkNqaR69IwiIJpG7BWxjAVhbS
NW4Xvooh3rKJh1vdNAyfti/RtIt4GQw6u06Py5adKs7oGJ9Gv6CvwSp7jFR//yWf
beRrjopF/WnoIQ5s/Djo+HqI4QiI+zUucR+vMHMVTykav7BvJoOQCIUBQY43qKki
NE7avGmLzpGS6vSprYi4oVPX34p1DcgEytVPJMwUNM5J0jVXjGeb94rNQawloQFh
gPAJpDa6xCJKi0Q7GZZp7UwaPWxwj0nQHo8MVdEbOIZ4mYCUpjgHKKtM50kHIUkd
MY7F0qa8xZLQXHpW8vn+pPOkM0aCjPOOMhJTROK531QT8UPgKGMcNu3nmBSbfeUg
4SelqdCQvPPmpeHZDNS9fY/6kG9XN5ag616Yne1WVsd5dcO5cZqJehtnfBXKOVlw
IiIm8pP6f+UbmD6KhYuKgL25714hniTUGY4o5GBkiy58mS4TVpkwlW9c+pswnGA0
dXE6YQNYJh1GGsvIaLs7ww6H4NqPVATkQrwgm5IpByAWvj2J3zHW2kkNKiXOJL20
FWxs9S+vqrzzqRBFj4EV5XxNIrMKO0XJ8r8BX7BSWMuFRL14JA3WNr9Y3M3RcWb6
Slv1havlWsVgZMfdl2IJF/gWH0I8mRY5nNLekscnjcqEmmnq/93JFYv3yVrNmP1q
pgy7W55bL8Aq5cGu870yEKONc4eDNLjY6LICpVahcnpKTsfGmTLNAzafq5Atc74g
22oe5uiyM8MORRBi7CMUwq6O1mPSPNvA8/QJfTK/wG1LKkDs/DUdNVQorXGZy1Na
GCo9zR9eWdQ85ZCbB7INMwX3Ueswxq1G/OepRRD3OZyOJ1oyRDuHsHRKSh8Kd+Lw
JjOJeig06fBRNHtPcgwS8eTBIqEf82qf1wMb6InSgWj8zke91vu/UOBIGK5Enm0V
nF+p629EbGl1rLcULdLBltaALUBcug2BbwxuDa88tJmTy/vURgrKw0POKrSBTuLb
zXSrOjONYp0AJOL399vo6LWck2LI21qjnpw1wBrbrvyUd6U/u6457XX2f1b9MMrv
OmD19r0eg8qOtwYn5Gm9SBwR4txfmnbml3a/jcIfzn18POzVVDdWdPp/P/Xwa6+V
X2tN2e3RUAg1CkCOcucqpytRq2uKgUD/WanoToIkUoLExjBncK4oY1BV5/kIV77Y
gXdqVDGhX+jAz2VpbP622d0UMtkS/dh8s7BM01EOOgq1e4XrgY9QF2YkV7InMWN8
hhj+nYrD+MFuZ/NZ97h4iQCAQ+5WFrNI4JjvIGQXgFGxENS6dI2CkB+dBIP2BoUD
mn3zCs1gl11P8q09ThNokltJqcY/rrw4FBMC4stoIjlQT/Bm2/In90w/BHbf345Y
06+whHOHbmt77wpRgeCEcCZAl5JuzEP+LQmZNu4D9ai8LfhRKugMcoGjc/ZRPlCc
upFSM7H7/WaUlf39rFzrWjxT8zyurjBjZfCOx4kFuAiaRXx84gM+0XzTmEhMvNHS
CiCHoAFHXmuvA/pz2gV/vxLhUqdKDSUrsIeeEPCslBDgz2empjfvkaGSbmybm2Vs
RnPDHY81X6XzqZpC4YLDInbqt6sWI5B07+IZ/4OTBAy466XZ/YSa13YDXYSEkuPW
L+MlDTsmRC902NjLZno9E6BSMLVVS00miskZTMUD/ilcYanclGgy+6kWCS4FKPWt
EW6Pp3d8rEaQXXg1QwJCLtfjriYOgdmLPugRcfDVJHLTSbm3r/iBXXejKRvvpNAg
cvQIUx/tqGZwGrvV5Xc43cAvbIkkSbP3bz+y8/vULOpKd1zlvBTg4LTj2KIIUDdU
Z1HsGTS3yTYJTPWAjXPcil+T9ySm/yOpTPYIgIpuM7+In9xqu8RlO0Z+vIWkwjAF
FvtcC/B90W64cRs0i7X3AlDB6bIOr9xdUufRq9osuB35ejhMB79dWC2tG0DDyTbc
gd8qS+8DEC2+cqDr28EyCffa/8PD8IYYoSV3HAN3mH4WOj+A/Fj4EeZHrh6+FPvz
awV7ugEifdtZzk/GHxWZzqLPKjHLB0oAzD1WVc00mrVzf9Wc6O2Mm/llc9XFG3/d
Wv+lpXwtrS+6ncTKeIB5PatBpZGGaqYeuTZHdbu5dsO/p4EgOGU9rYzpzVaJGOMl
5CO/BY/Z23G/Jr++BcKq8FARedZQlhkiPtBC9tHD+KytFaYKkvPafNS7N7QoLMfe
kNsrGWEpUKE4h/ltR6e2WZMtBl5gipgQFj17Kd68021XMM0/F8paHAcKbFicywhF
vk4twzOH9cmeXqyPv6ZRhdzq6g4/VBl9HzXQW27PJ1sWyE0vRkjxszuJKvvMh7Jd
/HJgOJgT0ouBMgHyHkbn9CpG/ZTR+qe3uuxHbWYvJTUHCZehIFM2rZ59IhAG1BFD
LB9DeYlPvxmk0s5WeZaHdLSoqYLQYOWXZqQjejKBQ9ErsaIfuKXAjHY9842xAEAr
Z+rK1MyTWVTltJkIZaPyAQizGmTIM9b17PiNHRqk1A891AOj87I7LlZkFuZW6HfQ
m8KnDMpjmNHXIevnin7rinGjtbQem+aVOYZ+SrxVSDa/L+ylAcOoYjUKEVN9P+pj
NswhQia7t1loBBn1IpN2CXMfGfFTQ1VTn+JmQA6coENr/Shja/5ekMW2pSDtw441
djvgjONY32MrvC0Bi5xKTg1D/TWj2qpvON549LaBD2cBkUBBpThr81s0H6gWVhG6
S/xa9C7zi8yXCQvqs/led762Pjl4gzxN9sfSr3uoj+MCds7E54ZSjca03E2wrPXS
buHs1hZzXNhlBOfzEAemdWAMTTtVG4WHPJXtxFsd0lqh6/32KBqOYEcMW6Ie21bG
+I0G2M7rG7Y9MBMzW3l5ZMUNen8JeWInZMB5Gp1WwgTXo9dGJf2kvL6qKa2YsATh
zv0iPSDvjT923LMMloLPlgfKvF6YXaIs2mx6MTNJspbeOMLluQxtW+uRMZ7PSrC0
UUm3cwbPYAe/AWGbGS+x8ieY2gFfPR8GHejzT+wu7FBzAoEn2JQHEIVRdKkr65gE
8g6vbNLq69PqWHO+wkYhgJppw4DFnXk7hPBqnZJY8OT8DOLCVzBTn0R0x7cVzRBR
FPtuJI6G+e8Acq0vPotUeyQr1BcgzHQnGw31speIuFfOWTkiQ8zqulXkXaVfTufe
XMF/8Cx/ugN+el9p0OUCsgGQ/Io9LebstRyxCZQUUN+kipjG4ARlR5WsbRqhiOfu
p++3EeMQiBjNkjeehxi9B3Z1d/IQfjmK40W7GE6V8nywztnbVEfh3QWzYNl9HZl1
DFVuEXzZAfR0fNCho+yhkPQmWbCCALltEbr78OxyRCVY+vjXStet8bIA/kQXSjp4
eXiSrqUMkEMcqeUg+xQ8MORdQwJcK1PH4P49GtgZEmq/u1xyERPGBUjVgfTawBfP
oAJ9Pz8QaueTmnsMDbJ7lQ7OmoQCEz6KdPGkkikjdmAVn2pF+QeHft1WM+jv2PwW
uOBo7RKTUKwfZqZ1/AnCtvmHhQVK0hJb/E3KyBCiDlkefkfkIFinArnBJwrEBSLo
fvrMPMkzPrTFrNm0BGwWNM02neu34RaL5WN9JB12F2s/eWh2kzGXd2inwq41Z9Ym
x3vktk50v3hdP5YGWA+aubEAWzxi11NDL+lozvG1PV+y/HQdqJUhPcs2MCXpIfEr
Wy+BDpZLcHuJA/m2gQ4TyRkFHO1KLeKOb/Cdb6vyt0LWLzmhqWPbpvftJcWIL9aF
39vXiM6rXlVpF3wD2cRpRAXVtm6IyWAn4b/h23+g0G1TzqISaBezlZiWS6BU0YaY
zapg6jQK+mCAPD6EoZTlN6Jmxecuf/zEQlZVNMybRvz9XAaEgWOVClbhqoU5BQbL
4Ldln21q4g0+ohaJ2m/2KDsah27t2YQm9+9Q01jUY23vymLcKrIJv2Vc44OaQbMa
3SCV1X3F5DAXv6RAD8jl/B/fUU9g4Dzztfn0QcCMQ36e3ZibYp+dQZdeD+IT6JHp
aoQuP8emcgJguU5Djz1ANVZpMfCtsVQacOB0F1yqqxi9f250e0YUqphU1FrX+utN
l1zjWb7c5uwQ8AlzQ20h21nCPsA1YofFkawuubFP/6f/MQ/O6TXgnswLe1DCORal
+efYXy+2lEWr0dLnKW+3H4jfyvntCFPiX1v48XV3N19gcOPgWtZU3bd8bdvLqMPy
X7EQn3PGVMYdxg4X6SYIxheUNCnr0TeRoy4bqbv2li1jG6Dvk6InnHJnCzrA67w7
3AyRF69KHJDwuB1y8vf4fAuTb7kz3qBSHY0G+rF7bsCpDik7upOHfXHuNHGGvDLD
Zq7ch+gIsUEAuyC9YA+mnCbDI0EkrVkyAVZzI1YMpCw37UQTUuK9fRxJcQ3/IOJI
Oy3Y+gB0COjOKEDoJCvk5Wn+WOPsBpRcAcnHeeD6op5WtUXQ66RWRsKe/u/7ZgkF
Dj2oTb+1mrqcKpkWFOGfHhu951M5VLrVMp4M88qkaOMnI9acVWWH3w7ZRm7keGLt
ZP43XvHY5yN8zlN6rp/8QfVHaEytjvwzwsqMEGxSDagUV/mxyEL6aqcS6jK7LcUE
7D9/zh/EBTn2nPwk0qzWO+rDu1/3USrQgypnep09CdJlUGXvhY5OT3bg54gLGe2m
QPlAT8AxfBnMpE7bnvBRkR+zFjuqjq321zezX3QAipvVcWiNhWfIVjX9ePPIOxZ2
uaPJU4Su98ySJ5BDL9VHrsT4VEz6seATKMXqIu2/rHhs8K1Dxx1rMRn1gI985obM
GLhtlcdUGqh9AvC7YzcQnefFITFTwOYnmJzghCu1K0kVn+A1M5H2eP2rWJimMKsv
k/T+vBQts7ViRG11TcjYgiD1+AbUOoeSk2O1QoONHS/zPL/QskYfmRcLFezHit9S
IlHAIbMK2Ns78S/GVf5pHOZ7HyZka39wpwW9jcmEPknkOSSe0hMnZ4uzBIbJPqze
1PgLAxZPD3KFKInH6dTt6cwAt8AkkeNlm0/veJjpoV0VvgTjVyslNa+x7Mnu75jv
bUp0dfeXjbmAiLEqZLJ3FbS/nkofUknyQ04+S6aWn8PutvqSnVuiSKZIsTyFPgvd
zwMlJRu9d4sN3ymbp2QFFMcMfwaEwu6VeUIGPz8KYDQjcmT/fdym0fObP+K2jC8d
wa/pSFwXxHps9X/f1lz/v4yRdTrd8J6R//sOAZ0qyS2unFLKqgqeJeN4fs/w4bhQ
XX+f64WdEupQtfMz5A6Hs3p8rqX8BriLQxRrJrXDcKBq2IDiHip2FJNDk14nZg1x
V57zTTzHSiBRItCQ8Lijd4o3Bph4Lr8LZ3iDqsHYkbkWNIcYf3nZu0DAX9mwJq8q
fT/tLXCimE9YG0zZnmVkD6BBl5jCFp1+Xsv2T4sw+1rI4Eh/j8L5J2bKAJsH8cZM
ZfuL9czaHL1m9OnkBpk8mn4w5CSXaepzHxXhhZhiNHgDFLFFCdPG4pIGu3gT7ayy
zWqXxwA7+hy454hqz9Q/m6bXPaW6O1yFtHxKeXNdV4xtXwMkvtVymVSOC7VU3dBG
IXzIOZ74KaTVvl+rxfO2D2YmrI5YVfASy5sT+oQlE3/K2It0OENrMecEDCZXBttf
wQHTSQRMKMidmF2mGZKtzzm6yCCS6AWN7pr/+0wexaADRlcq10s3TB03Jatj6tbk
w3scCLY60AOeFQ43MqtOJaeHxNcDze2Vxvj9dM5BwP4RRIMD58Nb7vOXwK8Pr3IO
EOaz9gJk0FrrJ3p+fMWxiwrBYMDbqOyXYkDtOfUUXp1XaGb5zSZZz31sfzTrgIHS
TE9n50GGzE8dB7WiTvird6tsM81skZ3hObdkAPEgzmKixPzkpteTEyPvrntP+Xd0
Uo59WE2GlLsDkVMAYrNVa5oFk4SCsNQKuQsrX1kaRuedeRGhY8+ABl8uY5u741gA
4JfDo82gc1aFHHOytGz6KcofcvfMRykWzZlJ7oS8NtwIwUTDwMbMrTLPKvR61qcL
mOyAcDIctysWxQgw5mxBKRNO0n1wjSCcYmrs7ZLUThc1zqZGyfJAjlUq3EDR/ZiP
1ITZ/S1Hk5tQCNxOfC6Z5Pyqziujwbp7eDOZWAzJJFkmQo8FYyPqElewdRm3g0NI
QbDdTzAkfvLxRfWi3JMz5uR/c5RfkCS290rxh0YRO9g5QybKv/Rf4SkyGbqknqRZ
L3nn9CHKDRnxHaToquUIf5Y5TZqIyTj7eKw4iu8SYL0U53pG8RhkZgjtOxsiYtyC
45DACFlilZfvMoQLIY8kqvWsWfXPhlYvyD4YFrvv/P7/wLOCR7JkgcraBphzuQKZ
p65oAwBIgdZf8EbUahMAXzEjrBRzOroHtqOvfvDcrGYipMAL1GfrETLVhgepyphL
p4NCjycfXm5Ry4mPsho4H7FQv3vDV/9N3f1cFVNwoygOhAzVsIsgSir2EMdYnrdV
Cty+uvcNSR7N5sBJYEgwwDjeG8Xp3n6gR+kMIYas7u0qKfNRW++dHrgxGjyIh6io
/LYCOufvHv98i44hR5+ILqauBitWAuWh7voyOBm7oigU6qDpo2si8nx31pAPeqtS
Xs9N5as+1MGdCgzdyjihIFZMgB8wObPply8MXe0/DqLwqnDkUqhSH2Tg3CgQgVNe
pShP8WSyOIhWBqiXPPXUS1CW0u2nMEuYkR7SyOGtC5P/2KZJtRH5HzvChNkXX8g8
QI/Odx273bPB59JJrviT9SWdvJKZXlRqYw103DyECLMFFvjPL1gsWnW01L21r/j2
z0Fi1GSwK2LpZVYWN8LevN58l7R7A/WEfd2FFXIvRZj3vAAmSfWgeuKkcBM4oPP9
JaAZZ7CbNzchT9AkYLwb6V+Rx9vl1kbWnWB2iZT0STILUhlyvrzQOiot/5o0hW7/
9Hqu0OcP+koiSZXhKyj3ppZwuHb9KbQSvZTXykw5xdkdzCpcWEFuDsU7kGYOV+kd
pcpTBu7xlbaHX8FAJ/bdDTA6PraqEuTstUKbj7U1gsu98YAOdG3FvtfR0rRjAV78
NX7ei7q/AdOtiTopgKifr6W08QvLVZlYuqgWomSuT6DhfrNVZ59XCJKd7uERUw6M
aSunHWnsNoRpwLgLblqCVRz8/WZF31QAmAvsEeAt35yh2f+YPGcw66tbuIhAsVHa
GsFUM775ml4ht2CasFKATv4yEZCqwvCS7LRQLcyMGxD2XP9Tc4oE5m3qQ2h++he7
gw32vlxc84EqoaggNyXx1Yhmgn3oCAj3kPcss34MvxobbJHOJOk6LzNzTDCH4l47
rCjEgN7KGqfsQ5GHNZf5UNGRb8syZfcrphQGAR0KSjh80+tgNJNAfXoubF+XkUic
eqjpQKNtGyN/k0IF3qqzv6gEmTXUBdMDyQ0/RW4OeaQEAgxHrGqblW0DCK6J6Vpc
Wp27p/mh/jfaY78OY5RfR45iLgNeVBa0kbfW2m/P5kVU7Bf0SOciB6mKWoNdwWPR
2fnxM4JyFtTLZoejDcRAtarWfyCNtYcVaVoFofe24Mdcubb6wSCq7y2CEKa4n9Cb
6q4mMjorKXoUgQMXfGlrHqOHOsxNt1DDKRv5yCcPKQ/FEsoa8gfBirOssAYmRlh6
DJbMxiX0fzk9l29h+UVW4GoH6URvccqmNNIykE81R81YsWeUQq5mEqrey7kFUcqV
ODpbVg0fwvv5hzczGUPcCkHFqoM5hHcYZbX+DftsPzM8rjuLuLABrC80imHZfagX
OViZD3gX5+4DSMXE7Ld7mpLisGYrkDPnBJT6mzLOo8vF4gTQvnaiGhvNR+qL6S0v
2mqUna2L7nZRMCsL8jb1GBXALf6ta2oSwXbQdLSNOjPOk8nThg7QvaerMavMnONW
IS6PLZqrVOXWFZ14ZxVpTgp/51qcHROcNSvBNWo2xN+go6qah8kpQnCsk1jTPSYg
97qjIp5eimdFYGbYbykVZyZ/OLakSqRDQLN1BAyrA/zVBRHU04LkK363Q2WvMBIG
0xR6Zm+83uKN4NZ9WdQ8ybW29fnC/E/ZzfQ3pfUHONs8ZHc+U0JhNYKqjWNUjKgW
41v5d4nz6SV70tmjGoLYh+GoSqKtJh2P4gQIhLmtn7ZwTNqJ4zy+0ri0yRkQrjSC
JvY3xxX9OH+h/X42TjfGYxD2aCUZgQlcN3tDuRpdo3Y9JEfFlRrFQmkA2p09BTnk
xUtPLZT/K6BusapyIpUTLarYZ8/X/vhDBWe9mXoobNFSeI6Mr50cXsJN3L6guIW4
X/iozMZD/6zaZpU/lPS8RF5gyNMT2TXcodSFb7N6wwqeb8FXDhcSaueGt+dmqGAb
YI12bXTRd6DDa5LpcubLmolS2R/t65ZD7hYqHQWrsLS8oGa+2BaT3i6OzzGq0WFB
0QB3n9NQ3QbjDbFWCBBkZHulmHJhXdFNuBY4ZGGbtXs1JTusYWogrAtpQSpcQyQH
Q+IAmosT08In2bOPuNlsX/l31V2fHxxGrYq6DYBdCiYc9+kTOjzvJ53PaV5PU96L
nCE2vRbdWwdCqIUENaaPaTh0fc1i5qyraq+76LWisI4M9yzd9eeXg+LmtRYRKLtq
xknb4+SXI2PNNSsiucXDTv3jUZNiI6YElqfGLpcl/MQMs6p3+nVYo1BYZZoU+m/D
oDBR2nM/+He4a0D9XEER/fEcE5vjLxhiCLE1dH1crrmdn/P+FGRlHiWJox6gymtE
qp31kYLGpjuGwt2QwhDvLr2mfRUu8ohyM+aezj21NC2mFmTKi2aZPq5Ly8PfIN32
/25uAISVUQcQt0QKJLFL5uZEysOjj/DyqCknra6hOQFFAf0N+HdeJGqjvj5OgZsA
aaQq1hQTzb9C7lJno7+f3MIsg6xYr59CVqQILSUpi/R0Iqbu/MU0WuiJKeZKZRZO
bW/BdCKn1OVfMkQk6BiiIKx669CLeubgItnXuB9B0KCFzWfUEMv/OWiF1czWN7kD
f9kP6shft0fN3SBF2EzJQPoje69OVBnFmAbH23cNaz1gPiFer/rQDal94/8C9MDy
JRYSJnhcbGjgJYo7+Bo76Gg5/Bh90VwwoElt2sijPGoSmIe5gk1TI60Ci8ClrGwR
adMseqDruUH0R2GCLYuWUjRIDl8ecStlxFtBo4+g7o39X72wWHneTeXjt5wOtkUu
IrygWMWZyOdkNL0vqYg7s4nDvvda6crZWrmFFEwXu/y7l1ITSLf69l+ANuJZmjSE
LdNRwNlKbRKWwIARu+Mfdhufgz2YkC897pfdno896apM90vrIn7y2mLzZM02VRq+
hsqvMUtoVxbiEhynBGEtOca6XNRqBpTjGfGnBORhkYic4AX6PSye1hDsC4Ntw6wj
rJa385Inmx7lIZeClOUsc62VkZ2lpAjdMWA+EL70/145ui2DSgnGXtWpo/3aMy2I
DLQYcBAsgObql1ZWB0pMxIUbSBxajj/0mGFYJe9EWnFlxdojAdl76PkAMWYLqO7h
qlzci8h99nrmaAg84S9wI0HG7f6wzdd4ttnUAamzAqN43aTBEBcB6wF3Wfk7Iq/S
ffPmZwIIxvWdAN4ymqoBzUInMMD2z1C1I/zHVUZLUnRo8eJ54UU6AmRCZL6MMOU3
ckSlIjJvst68w3ztOEflv4nCnWGdY1GxuvjaTk9DQZEeVS09SVvo1bTp+J3AFE7j
uFcRmW0HOkPRBhx2xgLUC+jzEYB77ftjcmOM+KJNpdqIlx9m2W2lY2Rt4ZOwVHdu
MeC0K/9rbKvTJIc0zLCre7Kp57qEhlv12drG8joKsmMPk5tRn0W9rgGq14gRj0j9
uQ06pLGXnJE2tAXFIzKzNvG2TxWZh0Gt96KksVmqGCInmfA1FUMnhT8YVHpeGv/a
EYO3baNLzID5ZscUHKz06p/oXRwKMJt9lw+GQPH0TvpcDBz9rBRYIWGfmI+0uupC
o4WYIZO67YZ/MsDcNU5AhftFeNNukKoOBndW/47qYkKL412xtV3cf8m1GfoolbDo
Uzs097ZfZLIdfvKNiOVJ3yI7p1WviLk2nHFqVNLmCiLVgSWxQNh1EswQ8ku4EkJc
zIbOV7VoVYUp4z1W4miBeOd5/4HADQEeWex6joMBNpVTjfALTw3AODec6bydOGqP
0oSnYMV5WPl6Cj5JhoofyOeoauxxpU7F6PywKta8G0BbEy7bixZbs1FbiY1svEaY
JvdR2g8dB3Zcvag1vOYCYkLjl+w6lFuibXSUJEA1t96rjl59cnLkm58GSsFJzP20
JwzOQFcMIe+gpnK5DFLMZ/w5VeNv5Dxb/m2wKg3CQx/fn1lRHXMZoxtawxDs7QTY
EeYqJShBVGr4CDLyJ1/2sWlZa+GOvotta8dnz5vR6k6rNA9D2odj5zK+TJuZk7Vi
rEoyOAYhDvMUqeTDidYY2AGdBvlv3APAKGWmWqtbQ8SC/RovJ+D0pUQglb0w9zaj
PctOK5iPZNSHhsgDzNQTGyJPKFt3Lcw9ljq+UHUsIll1Be4FKiVkWWYiJrqfs14+
0FHnVA/KawRv1uFdnzwxe9MRwTcR1QOluvOVP00s45G+jQFya4qPc2o8LJYK9/xm
gK1b+NXF8OejZ1vBqPltHP5YuiqVXfSblsIx9kG9pmKdxCuuMGJzbobd0QNev8+c
vozEADf/+ScsPLQMCmJpx14fK7Nzw0w4QO6PH+1/5MH/OpVVNK2ym95hYyvmTH/M
1wZ5Abja/b+kY5l0huTT+wKFK+UEpbrU19csXf9qaiGfw5uBDGMFzXbZ2A77oYJl
RX+HnRQWV/jqhIDbmJhZuHqHd79LLuZWJlhww4zNTbtsPi5Zg04p+fb571Oa+jrU
wlcvjGt2qtRy+Bh6TY2NcGLy1Fr5lCka2D/CVbE4R9dIfDP30YvURKVOuIFgI2Xo
aibXw92jcEVHV0rm6Prf0SbsGCyC1FniP0rsw45x/c8fIs7dqFldPKSEZ/primtK
hHMLPSLUpCrmPsFpVnF6BF2LDBAtvnHCQbBO2+ipslY+kd3jujRTYHU2OiOOZwMq
BSe0BKDOkFZOS9WV6ZtcqSWWyD5RPn6/UANU9tgRqJOe10UPAsr6td2BoUQI8JNC
D66Mii3ibesHdxlk+xzQt7xa5ICj4b2hLSPOCgQr9ks8dy2UeZmQAGKJP6/dMIpI
AZDn464jekQjbsEzQ58bDzyXprrpCh8AdhhayuPWEvtCrO46A+z/51Yq0da90LYX
JVExqZOf0zlWEHu2Q70SVlyLrO5hZrP/KAcn9DBFIDRITWdduRqFUsuYb3VPVSPJ
1y6NV+th6zcblRENEIf7fCh/wHJUw4t8GChZGy9eQnrYNjkT5Oe9KGfMy8hpf021
GXLaD94gOlF0+xVHw8M9tujkjvBpRKCPmn5yb4AQ9mBf/94Dw/QqmWNJQuWgnZ16
+B/+Naww3jmLm8+4i35ZyVGlkCnzjNJcS0O2ZvxT09M4xrJ1poh5WfsNosEpoRjj
uzpjz67Z0SAd8FvWhIs2LlN9M9ijb1+MTQcA63J7RIhoAg1o+qVNRj8ruIUOivTz
Zqi9WqEFaC0Ne+Qrmzm2p2ZwEYAwRqPf9oJgxoDZTXqK9gO4ZY5C6cmC39AhZmnd
zlvTuWTLyD7OusmZGwmIe7Op2ufMiTyqlt+et11xKbld3+bZiCobdeWw1VNebvbP
lGVB95G6GozoSotkT6JmJQS6Pgo3GMuQJ+/mnNxQQNw81XH/CwoSGcYVMNCK8QqG
onWLPRQjW623latYTJUD9EW8gBLwx4+oIyR1hr+xs6FhRXlqPlKofoPNGEHlxPBY
CkPS31tovH6GnIv5WGN4rnsvUvLxR8clamc3f83PEvQKAY0XwQbEsgZAk/GM4Gtu
tkBBsICjzqYWnWrNyxqipu/Mby42wZXnJwj/KI3pEsRZ3qnUbyRkGct5HQL5ecDw
mkCus6i+HHn1RhGa9XMHNZVC27KIGIO7Q+EiRpH/E5HgyLaCMV/nkY41L4YB3ysv
1EDkvQmAsCpT5VXj2oQkJywq2Ylik/vZc7jAS6gTiD3UvNMnqe6cUKEZjbpSud9h
96l5t+KPIsP1tyLh3pSjYDc+LAiOt/ZwUWIyApSMn2lqWqML+2aFfN+KBHhfLDUZ
EE9LWBF8+ZcBqSDZ0mILF0zu7YT3clOVNm6S3fXmEy8cq+Cwnp7oo52JLgaGg8g4
BJrqlLZ+N3kKUsZ78sZI7M/fEet65LbzU9CA7nydWQp4uhZfjNNw4SEmGafAHd4r
t76RUbTbI98lxnrmieZtGP2E1yVLbXtC8ZE/55nylO47o0vWWZwW8BXK7juJLEqE
zaf5QdbWN8znsD+/d5PRPK+VQNmcThQIrjk5fF4s7SGnx+6vvrhTuFqtfaxAS5r/
spJ3l+/gGajh13TR3iDhOmE3IsqhTs0n0PtyG/D2EHCE4r7kD8lpKiehGSVUVre1
M4P3zM89nRA9lobOxf0OfCmJPMePnTMXup92MubbyAVJ81re8BQJq9NV2751aef6
LLV6o5xAh9uFa2CfZhRW4lcraQTTkx60g9y4uiQLaPk3AjYvTQe5PXzrRYmfioeR
Z0/tqC9fdw76lCvx71XtUQePlmTYQeNPl1YpmkEt8eIaSoCeIGmDTmPD/Bnd9i9g
Ip1ulfQBkp9HxMNpG/dW5V4GcYT625Qg86PWTu18Tq+yimPnWlyy9WiPftZKaS8M
TutClgbCnywThz4a7BjwMninoUG0flywAQRvTEvVqCQ11e2QhnI1C9kNPpF9MmbP
Zw4UUsaomZaLY4jf4GXuGrkKgPgWkV5iA+/pdmh2cWl1iJoexkUhcc4TtRUnw5av
IwNiG3C8kHruzFd8ZLp7GADKkYIyEfjLT4c4e/JEOlXlqZBIVdZAdXWLK2DMDr/L
FfLBvb7d0mSnQdifCIrpmAU5J7iBnxvocRoluoERYxJVT+5DUMsAbKSYFkxdww3w
Cgz/XeOh+aK3BrBS5CQtIZ69osCxgiM53rEqsOawWViekT+neV740UGtgIEfO9gD
eSh+jkhzEPS11veCMERs3b3rZ2G4LtdMEB6nLhDgniiT5Z5+40lF6+yhAe3XnQqR
fiMq8dtzLw4mVmgXvoimhfJamc84FWhY7sBfwuiK1HJT56E7SfklOBYcYAd0SNTT
aN30OYYw72h5f9AoSiNk1qmPvEmi1QrRttz6e229VKNJnh+QUSI7YLB17y/zbrCV
2Oh/joc81f7/324JI/KRDN/gwwVFGMEIGGM4adrC4+bgHv9KWOUFUFmMVyxw84jn
b3LksT42eLUIDWGhHjj7whr+DrpE2H8g7YH64ck40HTYyaCThsKYQA1DD4KDSGa9
nl0lDMX8yYbBGT/D1cXK41Ac7+F4X3BJlSXpEHXlEkj33ghbxNoHOiIpua6q2ZYn
56zxAqLkFDCBNUK6hUafOem3QOF27q/9X7hujDb5SJs8wv0HmvQcSSF5iAIdeO17
0/b30/77nGVPcWUBvE/gqNuoTwm4WRLTkS8le4MKCtTPXdUuDELjHDXJiagSoOao
TD3dgSSw+ZR+Wd2G30F0/ywLSgCELyS2mOr/k+RO8Wgs30RVWdBrCvCTYHCev9zq
dqQoTC9nFFay5QokAwBvHOYQDKDIs00aHwV2e/+faBiTR6+LNYTLVJyE/xHpy77p
RUU3hmuJmHjMRaULG6g1Zvw5Y5JRWqiscudV9bAeCWaWf1ZUcTsep2pCQwVZkSAH
l51DVeuLf/d5mFd2xn69S4Bez8DOask4QyrVk6mmdrVrgJmT+8T7CNawG8hi1Nj2
VjEflyguNay6mdKMab9WuGwo52T5+xx7hHv/7wXYleCxmzeZdqOLIWTB4pSkitD0
MEC3trJJKPbToPyr6VRRUKAvlJOZIFjm7it4pUxIsiwxn2HZ5ygWKvhJZmAjLt4I
j/OPf5Pv1/NuOEsIEXGOcIlSsbEvuV4A7ERrjbc5ha7X73MOVRZQy5Qtdku5HK7t
dnV1mSC1YtAR6eDV0sAmR2OyxRdy5k7kifI7dGMgXItRbUw625z/R+gJTAjGx39W
R/G13vBuIu1+tha+/qBCJo5CY6zjZoaWAPheyWeZ1zRb1c3AfGDsurQfnYLDG5Jq
m5XFbNBPK9ojo2RP4sCN+x4mcnUM5gwL2EPC61Ny3Y6COqr8EDFnaHggcTBV6ELG
ScfJRdlK0eoEghFL4REjAizFdUCXOZuV1soxJB8R4PR0o85OmCMS/ajo9QI5Nv2g
IWbwyHes99Rz6ieLJK7X2mqzr/RgpdW18x0HAmEQlEz+ewwNL98/5braKL09wzG2
rhJBLi6i8Y1bZhu2fSP/OPnRCRVrd7ehcScdSEsZO8aExdj++GQrqEFmqpX4xCPo
0h9NwKNtKiHOo7+LXpmtLswpJIz9J6zbpLie9Z5fIbzeRkxF+kGKQztGCe1yIbpE
baNUla0tohy2sfJApdKXQ3u1Mqu0IutlrXIOWEFNefeWnJQPNqgbMk0N9xvhSTbO
O6qVQXjnwsJYy2z5qQAJYSS0WPyveFYDGxAFcwCML53hEUBP4Dp4hLzGGNFAv5S4
J0xsKaFgu8qu1nLbslXIJqtbC4XUeDDwowv6KS7Obi3HsL2m+aml3kjUqZEPbbvh
PZ+Ym3QKGHI5JlBHbU+H0Ht7qyN87vJZx/L+4gQ5B+n8t0ZmWEVN3jly4Viy+7ZC
OoWpVO0h8+op4ynjHcU675CVjwshAqgQZJaYXssJ/vWzrVUb3800BoIHWnGGlJsF
tfJGvmuJji3ZO59ZL3/DtJ0YybsZCZIF9DkxIikP23DXVsGHOWG6Juf7etkJwGjo
KZzjNz3MEGsqkUq2rnv4SKNdtFGlaSABY7Bf5QXULFXhhn1wRt7Gg4QLoJOnrxxY
ojQQz3heHX2Rxotg91UN8Q21ph0t8hE0A5b07oKYi6o1cXje/6WI5z1IaM90WFo4
BQJGf0hiy8jSJ9Q7gSUTxgaTWQbLNLiZKkSXf8vPPUcS1MZ/OXd3RbjQFklqlxo9
+7ni3lCa5mPsatsiwxojb+35YV262LjOaIxCqcLLZz7fJQekoV0PmQs03pO7v162
Oeuvr9nQVqju0qt4ZBl3e+vJbwb1BWfQkCpe5MuIvxW7C49zjuho8D5RGkRVGYpe
2zNFlJWsOuwiEhFrDwj+g6Jj7TsllEVLbGUaDdL7yUmCQ4W8LTOu6T5SZrhm48d1
zBblLk34SSl/ZSMmTUgKsNLghOICe1sjtpuKW5zEPdwfjEuDpRO4jkUmMMOpmcqq
kGSY0Y4ufTFqNdmFqAXsJXtWxIvYj1zLMOvtGFm0FbupbIC/ghb8M/3ggZnxNrpP
PrFXDw14Mw/Sw86IAW6WbfHFnRQ7hxaKyBgG3qfNvTTNgS/HCxtPTO3YpTkuT15K
TAz7h/bHN9rxtbT7svQ33cm4bbGQ5sREPMH94fzDsOJSBxtpBTDV+oPTJ07AYQOU
q8mkkr8uZ5H3Gof+PDSdrRncOx1WCIeq8l3ET0/KOsigka9wUpzr8PrSXdVVLeZ9
3Tr/mxQ1dZbUCvq1FWNMxkrb1VG8a8NpjJWahy8ZQlCQ+ZtzsC2E0Xa3M6Yk5S9y
A0LVfuLP9/nfEmfIOPODOIaIvAaTVWX8bShBU4BjD6TslP2bP27wP1OuEYH+vHWS
EtBA+tylk/FbXU0ykaWPBGWF7ljtGc5ALPTPqvpCEh5R0j5Vpnf33PtaOpc5cR3w
U1/4MKMyV3S+rPR3jW02CYma7geVj4vxc8GASFOv3cxnbeE3+gTuHOWrqoGuwAl5
Vw0KB7weE7d91iwqlrA6naLoUgkLAOhQYYZVY/peATyiFv2OvRbs14sgEp1i77Vr
KYjz/wRUbsaVZBt4po17hbmfPMxxRAkU6to7br76VKl1WFKuR93tHgjT1Ux9mNIs
paSZU4GxzrAme0bmRywXauF7Khs243AHO/LBb8xdDKOButkdFHBKxzcYQcf+llU+
eveZXB/Klm3Bkg8S5ns6ttr5PnRRzV1I01SCVVoV/wfZ17dYKgvRtN1fdTeoglRj
J33LFStgLSRPkg2vqVlg2pUvj7/vrVxAhpWoLiYGqHy5SaascC5HPJngQ5zFZkLM
AWYat2ZfIVb6s2mZQj9TCe8MeyUJrhX3qSPk5hwvPbS9mdcRFnKCkY5nobDoM+x8
Chxut/ad3Q33kOAl4CjL6BhlyJ7Ik7q80fJd6mCZWmkkRr4MizAXZjGB7R8lBsWZ
mJq6hyabAjktC5tG78RV62hG5AGr2trZ+UuNt0JoyMJvDlGmMkcODAcg+3WG2vTo
e78AZs9OgtRPxQ+OeErOYHLQYlt4G+1Wlv89mHFnwK3p1xwI4KvkGZ7v56ed84YX
YPkzS166XixrrPfEjJcNPx8Izp42f6dPaoRTxGcKzQZNG7XWRE8FI4k3vcae6iMp
+dMH53XcK8bEOSzyGeMGs8ryqGNhA4S5kd7CkQBtkPLAAe+iURJWTBqlWQXKs1xp
CthLdtllqXFlM+Y4tiK0kfOfPsJrBMbqmiPBBzvN493NxVWLxd52EvpyNQzyrHx4
krKBUU4KOGDhZmj8zCtFXp5o9ixdaIKyqghWzMAHBHq49J1zDiR158fgo4pMMmXL
Qt32ih1Gv6FM5n4LhjW+ypenHkPTG9KZsdgDpOQ56+d4c//xhKJLhMmyzGCpUevW
sOBoY6oceLvZOoaO5n11THsFByF1UAeUebiyl3ubJ9tuG9t+AOjREeeFXn56y6ao
tb2LVJtm7KpGaUdPVJbgQSYAurQkFCUZeOXj5Qo4hyPO2yXyvcuW2NRCy6wBgdCb
NGD3pwiIup3QCesAbfVimfVhDFqL+wPn1fzYtxJelrMzTxiZzlT+cMHQyuXWYk46
GoAzSf5uUKEEBRsth2tNBFwheXBDdWHpMwSj9ikLVuOblZ3csDgWmSOEpn2rf+gd
itO/yGaQwA1NzogVnt0q1Lxg2ATUfY7w+6A9aXduXFi4SaUxdbkrtJnaIxQsB7ce
GYRwPx0ihzwxLnaQuFaPzrx+J6OqZmrrfaPI4tBuOxyj59ARHTh+eKrrPJV38POR
UsIIpzL8oVN1Vp6AHqosZ6P+wbBodg3xlH1LpcpG7qcbKmkoJdqGGjJ0DS3pvVC9
xGznt76zzRCrXNOkfl8QB2NnHXtwknh9gVEWYMHUcGOd7Ltj6aXkn6r2XtMXWcWk
sisd8OkmvTZQtrR3Hxc2fuexgP1kXyYBR9tSDO0JKy/wDF58+eEjh+ncyzU8A+66
nsUhnsuOutCS0YIvIfR6rqU9bNTDip401lMhGosgJzQnVjStN6FwTbSDd/ZW+U+k
75aOosJEDP7HuY9/z7Wt6oKJATvbyZ9kZbCBu7qDM8h7MsLgRGWYVnXBtw2jgJvF
34zZNl3cSuh+oMFugjE+MO6N+ZIDYxGMMSuZxAo7/88SvIFdx6kNgoTS3T3ogznE
8xdowGUdjIzuxFXSSt5YuVSu2KX1ilIxR8pRCnGoOSGxwmEJ8RooKVUYL+hw009c
KddZMV+QSHn4doJw3W67KuWeI7ap0S+gePyqa4inNNh13gNBeLHf6g7unmLoBX8o
y8wFDAdMV0cE16kMaRDFZMX1XC0HLsav2FpGp9f6WgJXhCAfRMNHp4hrtp3mGLk1
Rjoup7HGLEebqeE+Uv8wbpLtYPLMDBBaDCOShq166DlA2qtrju3ldMD7HuURU7Sb
JDzxZ5UQgOJJTQ/h4j8FYiRfSv7Q5LQToul1qztRzlqHBkNZ+k6PNXZEZoR3Ob1Z
Z2wKnksHxuyWBTdmMmWETkZ5lV76YsyfFc5XqkrDIU/jn3rVtUTProPozTfefae/
7McFU2g1ip0Or5s20VBK+dwnOWFUV3OVGoCSUYwnQxuuCEtqmXXWDzGvMfJB0dnc
1WfHvg2zzZHXLZNao3kff4NPM61NpKaPFos82229WBV7aI0RcOOpjLXiVTZ3h/7T
hwN9tWGRYQbNnOEPWc9KZKs29rasoneutnUB1xm0FZKBTMYlllMaucqGBaj/wxvI
Kl1WZ9uD45PFwitxdyCD4mx3lPsnfpl3kTRR/vzrkekLvWzqvHgOmNGIUxAkCy1O
52jkRjryB0UxjcmYe0Yeawm9O3X0hdAXY1tc80OLrXFR2CbnTLb6rg7Eh8nk4R8X
C/6xEEWZx3kj6lrDQqxDdySUmdH3zBviJYmglWPCLK5iol0b/TRpHx2aOSwZjS0X
QxDAWUYxmSnkIUagv1zN8lf2MekRZOWxsNUesQSZxsLG4y20W62rI7sw+M9XIq22
U/oo530eRqtYTY4dKSfBSVK+VldmPaafkvfSYsFuOt9O4UREW3k2fxpieAqR843s
P1PPwa3uxtf5UvJQsMtWl5NqUU5g+rE2BLVydiEl/ngl2kkNkN0989iWlJrpwlkz
qTDk0VRGyvccW7EIOd1PpDsrl4Vot4SRWoAPNGts+pO4n9rMbUROuq9d/EacRwTE
lxcSn3nry+KkBU8n1ihAnbgS3X1d7m/sPGpXK+h5W7yO2QuHt2Pdaelodl4UKLTB
wb5mtKBYfuZYEJJvCzoEeH9Z5r/mTuJQmk89hy1CK332FbSoEMgH3bafjFey1QV9
p0dwMtCIdb0QnVbGlFA++4Im6K8e1Xr/CMfKMFy2OLkZEchPeaTzOl/hWJ4y1YjP
llWmwTUfrRqa1Vq7Jd7LHv0ogJOl9n9M5H22avbQ2vR66WTl6ylWfDkGlpMlzTEd
oemCgQrfB1PjQeVPZ4t6aM+ixkxCkiXbwZaVNhY8UF0CP+FpYIx5cXPTijQrMm0Q
/sCrd/23CAZfXjMu4BYcL2gPxuSumwdUl+mxncuStQ6GUrQkG4xVPVysNZCEMOPI
Ag/x3LEm8yK+gJdzCuNe5p/wNNJ9fT45HQUEYqqqbFtiRB2U1FQsxWS1S2OTf/Pd
xSjQkT8qtcf8/hfMFVgaZC7w39rXaTKv9hUgtGPWM+mtEVmYC3fnaJipEfZlZJGt
D42oW5udgnK9fU/Ps5BHLLSiw9B0dpoZkcw66rdSKAtlIb6Z95ohMQSOKul28FIt
dX3+YEipcMxfoZ3i8nN7RcaTkvagSoWCe/XNm8ak4RrWO6yu5f15gPjEa3pJijIK
oKENgm5abSzYLOeUEzez39qtYwlkoY+V9iJ9Wigery8SNEpPsQUa/yLr6Ad7c1Y7
pAtXuPSdxhwip4f9AR1QdGUDIM/MT9vdiyIEg8NGgdC9AUTj1cOmtPpQhnvS96ew
rhFEx+PBvkcMKiriE2mTm4YPGNioJGFtlaOC814HQ25XVKZs+2l2dtYkGtwMWpcL
4lSBYzyKcZk2FnIHIXQ691mw5tSZxoW+94KRUQTr356NAOE7OY60kWOgXbJd+bt1
RKXtpjdq0VnSeb6BF/U/xcknso0ft5bkErOi8QFF/Hz6ZmWNwsO6mkpLC7+U0iV/
onirZ0Zh95gRzgl8sqtradYKsF9Ige6pDPbp41EcGtRfG7USkZ3tyeaTjS9lb7qN
OpOS2a0UkjcGfN17lTWHaXCXClK08j4xgZTgmw+BUKnV1QoLqGj2DbRf65QDkQeK
3UEi57j95CouG6YVgF7U2mAOwWqiMGmTaIf0GITsWjzNcPPZjn4ma+oNuCaXdMA+
fngQ74C0977Gvrv6WrkeGV7REcv69daUzmDcNpLh/DkPr6MaUUUqBo/P0kHT5J2k
8h4U4ackRsdYp7CowN9DbYTvv4rQmJ7OSMG+ZggrnTMqp8wKvMCpsD7D4gZ0t+02
swLuIGoSDnB8Zk2cyDjcpkEVhj1Z2CmNTX5G+dA5q417Gt4ibuYqSg1DXL6LPbol
btMm8qcaQJKri0RHG3S8Cd/PbP85ycSvdvWx1RDTAEGZmAL9dp6qRITpM75Bqc89
tG48BzSpY8qTOTkBlsBVLQl5kOv9I+8OyOLpGUZIM/ncwS49Pj7OQChm9/YwX1M2
puXCSVkRULStE73wNptHPruG/lh1Pe7XjHneQ48mKNJ1cWZuOibmpKbwUVQvnBmh
xQtxBKyzExXrdmu9mmALp2imI1MKddIbaCxgaTPDxo+BEQRM/MMqKtAoYG2ZROs1
2nlhJ45eYBsRflOiQgquF1+Ahv1bK2BHG23HmEZsILllHbhn2RQkk6VJ0v5avr3O
WnyglCuLRNMkEcXod8YphUJeCsufi/e/LZ3eCjyocrYjBd28LpQa8LqncnJsg0xm
0qIvniwqQmkRIgmQG4OIietjkxrtVVys7D3h1F+0YSPkTyrqRYYvC7XFAEsuPJUj
swup8ZTNPOmbnr8a/bPQIjt9FXHk/ZEjnQizjKS+D4bOtiQWKcxmWQLUjz32eE9a
ZNj1Lv0vIC0TByJizSdom4y4I81+STuUWbVCaimByx7BMkiNq1D63e6a4Hw9Jtfz
O5p2AK+MWRhS+l4EYwe/yD3BV3gP9wjjYAq8XeUXObUYu2ayO0aKkReZK/CvYMmf
2IlfAjQCeCZDGvRyLT5jVKNYL5NzUp2ffIJUbFAt2vriW7iiTrPBS2JZJ+bZMvWu
hE3KFrgjUrv4YTIyNw9CzJu2DfdR1X6poRvFhqPgeWRgskl+iWkwgv8LEAZg/Ibg
eScCZJTX3np91EDYmSljYm6GBtm/WsAGGUYq4kB6lzAq8ys4j091exQ8qwXFFfmB
v6TgrnyN6ECB0i2c47zLDP1FAwRJ+QZqX4UpOOTaecgclIVbNqSgAPdEkSXB9otR
WebXS9jQtS7mJKQ03yLnsGx+jBmYnajp3dypnjPQiKx6QZ/ByvmhWZsvMReP6soU
iFN9Z6UI0vq3md2IQvvH+3VbuDMY7r3Wanrhm9jIHYHC7zGZQyGgLY0ohuVtX1bm
hw1uNasrHryBWpNnjlw3RvaP+dc2ga+rsv6KC5fv66949QVQUyMetpkGE5EOrnsW
3KfsmbSo6fj2GPX4+HXx8EWREGTTw1R1YpEZXPRO3SRRsmT7dc72R9xAE8Narlni
fc6nuf/iptvd0yHUIiPrYbphn/iQRnsY2qb/d/hGwMdRZ3tjP0Ggm5T9mGvXdkEX
NayNCAoG5WDkn56BzF3bM7MOMY6dVHFivccFScLlJ6a++rFbmxlMrHxes3+uYp3U
L/svCkz7Lh2gMPg5woHpicVFhaJiIklovprs7tW5lfqRsTZr6qFSWWTiUrRUZi0B
6rmTNo+T8w4jv9jZTldfGUpdSKCMAtDwAAx8Wzdz493sH1ZJF2+OlFRkDuqh5bIo
H8/MMCAUH8XgJ2Ks3whwmRI+IymeMdTtOj2n3x2I3JwFV3hHs/Ht7kFm6aBTEawr
2LjEdkf8/SFQMlAjs4/b1ozMv2Rcegx8bCvWlzj69sAIch1sgfU0NnwCWC5fvF5h
U8aCXYYo+dX3/UJPc6dGUYsvE7A6zSxdZc+89x66Z/O131ntB42LItNcOHl3NFDS
xNPw1CF9I5AtsiP/tjGttqNb1JZNIa4Gvb65fP1hLwVi96s9CcIP4sJVGPIPnew4
y+fUSjJUaoOQwQauCs6G+yWHZtUK8pbCT3P9UUnlBAJpa2YxCXoTtPK5HxhtIXqk
ekSBgC3mkxWJmKbyTLkzeOdR8q7b/UdivV8tUo+kqB5z+EbFabS5Df7wBS/DHgIq
Xmi4MV3EMRUOMKL2vEuK2OqF5ojmTY+mLmEAazxB4fILwFW5B8W1mVLdxE8xZdyb
23p6NLaoheDzWS+Ij6qZx5fqgz68/tRpJSAjldUYXqxomLTHiNHEjNUMOzJw/Y2u
wyb4p+iqM+IG8ooBYCBtMILKAzchdqfzyqwTpbZzHpjhS8T+5ZU0sJ/2oLRXK9Rp
NUMtzcAdJzmxeQOpoz4vcFhYPvy3lmegorTJJB6wFHze0am2IDito3U02AHStSFg
QA+ucNsyFKrVdgOhRP3Xhe2k80wIYQMH/P4rZARWWQIhKUmxKy6szREuXnbfmOuC
M1HXoSVGivLHYOvjnadutOvtoII29Rk4pVnZNicvSnYCSi2slK5bxlG+QbOgSO7G
30DHMrQwXv1WiFHPjfUuu+eu3yuoMYTb33iNrfOKouXW1krrDLa/2ysUI9yk1+Wy
r4zTRtYPfKyPAc1BGUGlU9Bl/nlTPLWlvagFbrCG/6B7kKudNCp2oSBDK+3CxMvV
EwuWlSi01qOi2Ul7HRCfh9V9Tnwo3OR0wIdhFKQmTbP2JducFvwNoEFuY2qa9eTZ
ujGOWHROoF3dtubfYFz9Q7NdmafzNgyrs2hbowwq5u6UNKrafqXLIRYdMHhgDW9n
aGo+GyX9E9B5Un7jQbJD68s0ZlY/U96q5zG+d0SQEF844lv+6IwgVv4x7GBYLIQQ
yHAdO0gYig0OCnVe+tDVkc/+aWNoyXxyJNemXiBwQYDNfXzcKCVY7G4/z1yQKmVX
MHVmuOxv7m7YuanE1hW1Qs6f+9hIxJdhIw1U6GMvPKny8OcAaFEsOCQJTgTnuhot
ttx0R7Yyq00OUmz02H+GwjX4SgoicRIqyd6396edHw36GTH1bidgkTZaxt+X/3a1
ucM0AJ0u6eFc4wAodNkFfuUQomMgb/twb+CwWxA11t2FCA8bXGAkgl5zIW+duA7c
fuwwSy5SPtt1/YhO7lnSmIclO23/0RYax7qYi1Tq62WdAqorq7BYGkQRSDO8LBfP
vATHH4xOn1UDSxg9N/rsj5lUNnVL1jmJ0pYG2Rfl+gCEfbAelqKw8sBPYiCgoXOF
MZe4I6GJ/zhTlg+XGKRP4kc0lFUEzhMKN9dBkYiIghPs5HWS9VE+W2/7Vd4egff3
XUT8V6i/QMge1ralXBCJiAXolSJsh4l3lCTEbb9qcPF3PLJnu8sq+fbD+GW3vQVG
IMvN8u7SOA4Sj6ugIFtM6ZnAmVBX6Ql9aaEfJTeW+zvpgJYjcTG4AZSyUGbwhgMt
UStqs2Htv5OEil1964fqO/iD/1PLJxYmFOjlLbTLDMVI/IB9CqxQZLpeWq1xgW0X
GOAFjZjsVdCexVGE5kcJe0CrNxPjWOf7kNrt9QoinRST9Ib3DZ7DnRJSeCA/6HGJ
vj3Dp+MHX6rnWHwyBsSDl/ZWZhSDJBxIdVJTtzWXXXuYMLYdRme72kK0Vuf2hLYI
EbSw1DuJkWUvqNWzQECUGfycEskh7bHzHoLyrDQ3rg0PJJhwL6O4d+8Ew08J8wdf
o3Zl5vNsp182TEKFp0bxv/zGGdA4O/ija9tdpxPYDCvpP11aSNdP85uYIOSPC4C1
BETz7XrZptBH1WOwP2hQfMFsr2O6ANISaDJHuyHiE5SorUIA+hP7QVnCe1nq3AB0
MOd/JjA99mlN50ct3OjkbSDTEloZkRojpGLbJC+/GIrFS9lZjQ4tpunjQ0JL0bv6
ZFuHfVrMi+aoN7i2gpJyYoLceices3+CWMsmZ6Qd9rn3L1AYhpoes9kpw97tfFq7
c+q9r2/iGzVB6kmdfx3TGDtc2HIpo2jKX/Mp4BKw/+2yAY4dHivo/LNPSwLOq0QV
nr5F59Ltw6r1WXKqtGJxnGimeVBx9ty2cnfOQRiLa9BkcEWU8vUkxQVk8yWvndz9
LGel7QCMaqcaF2l90WjnOyK6mFc/dyTqL07kJLI46kW14Plkvo3HYOkDc/r3lOM/
j/svPF5Ot2DXrurgoznXCRmwKG/LZaQSZnarwsrjRi+CXyTcOjgp0vsuNyj9ieUY
SFMbrk/hSjGrI3EAStmiOp4NGyaknQUoaSzyQY1Ml2bTV56xIMDv2DB2HAUD2jIP
DDGWTk5/cnxUoE2IVTvKsApdPC8OcFGBYBzNzL0N7VRpoZ1KGpgXIfanRIGOMsk3
R2JEy5nMTccTm/XKn9+vwphw4g7/fBLGXVED/5sDFGjHyyPyf1X4w8Pq8KA5DxbU
Ie4wJWKmDtF9pw6S/5FEkncKChGPMtqUfS7mkSSrAHasGA+zjOdc47zqUfWZ5hiR
SZaZUrKnxc1eBCNTUwfW0/3twdL8ysN6VRDvbyMXtqPkVrilpFkZhe5TKvI15lxD
dNzOGBXXckRwelam9ZcEqw2xqRZwW8HzldzM9Sff8OzKeXv2BM1+ZIO5gbOqV64G
+NnTP8zFx3fWhkfP/FZZGHxwn5DIn+AcREZpV1KJju0Mv7ROgO05J/mLSZyrq6l2
P4fJrVU3ffYalc1lJMwCTBYPd7cLctdaWzMhwj46QHBdHkocXQ8ULheB3zWrqve0
ayhw+CFp29J2AeQWGu2hWxwMcgVNxqTEDXqPByqo83gzgjEME7t3HmUMEVvvpRlT
BLEvN1AzR4lkEJrcs9IkTkKMpCHRrHrhYZ4CJ1TizNcsZqLQPq3SFPEJbomiaFmn
Ylq6iwxBcbTAEYa1YFbz26e799yGZromzT5uwRF74T3YNkG8gZzI0LKqKEaPdtvQ
hzAk1wklsNZZDbmZ0khSQAzXDAjbkUz3gQI8BuqY4q75/56wzJgyjulvvAGNKgr8
aGHgB48BpMU7g0Vvgx3BkezOGK5rs35UpW/VEgslbV5j+LCmTQFa0J1M/BZDOjlz
0tMAU7Tl8hPzXmdpLfrteRVHseMT55TqynhYEtia5+FM5tThYmVLkUfUlI+hZmxf
XkOHHD6lfMz83t/8PRpTdnIzb7pBWPQgE/T84vA0UytmR2PwRaFdRLsvptOrH5J3
aRsGiInJRCnTSk/bBJx7PdmGj85yBygeBAl5Q+Vcr/nxzD781Ggg5I1ndz7SniPX
i7rJGz8yz9Z9KN3CaEZv1UDParVq8K+9sUS3DUI7RGWbK376Jn4abmMExO+X1h+u
+k8w9v0Wo7sbpaznC9Hu7Oh5HgzMjwztvo8YEH02++FrnL4NYslXGTWzbPECuOnS
NlQnsYoBt0X0sw/FbJShghemYsDHIZC+ZDvlCMkJatiwUi3QTdevE4Qq7uTD/KlQ
KHCE21h2ZLngMiv2BBKdspv6KlKkqpDWlxgdKCB107QQErayysopLdURd4uYl786
39NvrqtcKvApw78l4giZaWza+taAZAOP+vt6oL6uEL2FaolTzqJdzNWPjVELHpeX
gNslyRtDNjpB4pa624xZSRBazSs6f43B436rKdsBqcZ1GclXWM+8N0rTnrJC/fh4
YfPhXAs3XO8fenNDafBKOc1y3ndRzFYlxqk8UQlNLio/dPTDcahlu03rKPE8r2H/
VfGhAsH+056qGPCDx2O0WCYOqN8rd9XwCoG962vhkAez6QmdmoYZw3i469ObSmzv
4BGnV/ktmnqyUN7kfsvIjjQqG5CvmWqNnHpJdRPsHnvwmmlkIFdxMXxjto35bk5i
udoJgNNkjQdzvnRIhV+gA++kiOju7h3lj0lO8nldtLOww25fAtlgPsyt7pdzF1tP
ESQE5NhXimA5aUl4PoyvmEJ180bxw9kHqt72+pvorb/fklKGSKN5Bc8REcAWNHAs
WDMuNp8Bn4bBRlzNObsXQMbfoQN4yaexHMxY78pGkR3ACCBiiSZuZT/rZPcMhceb
+4XeMnGn5Rvm7fCD1q6G6jV+ObzNU6pw5USqHrrFe9ku5ba6KSlhjHt6yzERrJCO
XCY9cAfqPrvJVz3sxmbVrUXQB8bpkD4nrnTgaEzhcQCTMsbihLznR6t7G+eEHzA+
M+oahhQyHqorodzXiC93AWyry1352rovHRxCoI2Z2e1k2CSp8XzIhEcpFb9gGMYj
ViEX5uVASP5yElT2TiJTZbm7vG2HijChvh36fFTxFH1C9PWXI2h1iWlAksYroNFN
VGoLSMCAz0PIa/fEHCdZ2eRKws3C0XEnXqpDoG9BzU1SaMUH2J4LIP2sUBDNmB2l
oqv8kfE/ZKpeSE2Oz8Olw6xHdo6gHRleDKlrn4Y0IiA30c1dkXHQXfKst2Owmyg7
xDt12E/hiVEFk5lGxpz/hn1TVm+KGst4BU2t5phNPh8wFBsmwKjeHThtzvuTQj+E
y8M0kenokogVcSFRHcq4QkKjYqq+NvIod6tvSJQPPi9ZlMMAVkanMV71SID5hJUp
Mrm9OYWoyXJzm4UrBpFYYc8KbK4edpuN3JCVMNYxwGCpOwufpUSx5a2JG4nPVz6X
QamM6141zSzzn7K2JI1+QScxl3YAMQilCHwc4Yh7wbJKyCw6Yj5SoNelf0eGU0D2
JuUwIKuwcXUSPj9V0iSZBFO+/p6BK7ocUZcxEnnkXZl3/y70LetYEQUtCrg/hkvg
0naVJuOjTA7VJLPROPL8zncTBeH/VT8I5+HffcWBGOC98ITNb9CYILBpWzOroji4
LHP8UlAp3Cyid8xzRWSQLctfboBezP2noRiKUrMcA1UFtyCcSZFe240UsDyg08ei
7J1WVsZXn+2EnfLkWDDTnUPCfSqT5M2Zoce3sKCY3GJ0dJmyDiyoEGCO0Sr6gxEE
2zHmd91pnFm8tqzdrPNgahVJ4+m4171z8TOsYX36rN215tS5bVlBZThjn/klc8LE
nlTGfCxGV55cGtjHch3DxhhMzE9IIkwl9ggbyA4jj+Zy8NO7VmEH4+XTWTS6fBsm
g4E5mya1+Jx7QFiTj+RCqK4ef6uxZDUNruMbDtFBPh/3lxNpQzGs+jbDiwtypKwJ
5GdqRrzr2ntOpIqnKKS4v+YnLnxbL8o0EFaaLmN+3YRpQcR0WxiETUbzuQcsocG6
qduIK34+LrkBbyBDYEVKqNyDTmfbduTUl10TB5MeQZsXIO31nv3fc9DIPCt/6Rgf
/oK6972MMmlmUqyVPSJdyym8wRVof976FyXUrKlU91xZ9gYKZ9NdcwPAgANyjUNS
d8dZfYKZcP6LukXxKwwmFFphFkuIhhIlh+EMtJoZmtRVfX6Fqa7m8ugIXxxIbTuG
rnEdKdG+BCB5qZ7OAmdjVNCbrJgtEbRpFC3ckkdbesrEn4Dscwu8WDVkLiPkMaWd
JBxcDt8e9osL/56E49mSJylsGW3DJrqPBY2Xf/VDRDiaMar3lXXBKOoE0LNX2P5G
RmxMjmlrxDUH8EeCxVjkErj6D1m6CF4DJWl6lo9KCWPZnPxsFOLw1TyahmVYeIkj
hvaV8sdTfHmd9NuoWwatptuqyUVFa0DMWXaIZta5yUu2ruTvs1XyRtm6J90G/m18
9WlQUzr2BwIsVVg2xgxcbvWJRhgtlwU1+5UXktmpTsc1uV9BJxYCs3VfG3WQ8u8r
A0MV1bO/yMtful/3hKPC4me8FU5dlXhSL8wAOlGl90Vt4Qf7I+jQOoXjy9ZJQ1TI
8TW7O5Mzo+ifETZnf8xW1o5Pmj2yCVk9m28xEA/koVktHo8jeoVAK86KReniR5Ye
BtMdTozpFLtpNQKSwoiHUHR0sC2LHksVIYBV9pYgVTK3dtioTcM8C0PYbCwB7LLF
RUvT4G7zpq9Yfi5eAYAmyJFsC6JKddybWgvNz/eMo4ZFy56c1oBW9mEu8AJKU4tj
xC5S6eBxeTBv2ogIWa8urTkK97iOUHocGBevS7LdXqkE1odXOh9wDPSgRP3yfNrD
mPl5ppjXThuO6VrOyGMDgFBzBlvK4WqMZfk5qsSojtLAMHG7LVIr6MVhYkv1g+ry
cTv2bC/JnBswHJVlAtt5joYFjr3zTjE3fPFpQDBOLPllJBgf2itHzk72deNAAe/n
n5BcuV0H1SK2xI+6iOEnnifeWn0Dmi0HPDPvnPyQfqp89a5aj8RRlRN8SrhqKFMF
tvTe9iJPEtJYIimA96GKP152uCHll+zccWwKjTRvZhWqbESPmnTIcZEk234uMjzy
yUoVwSmHtP026LF1GQhIAz+78mqT8SELuwEv0t8VJVTDrcuZTMcxz2PUR1+iaxDw
i97xU26eM6RTQIPjuXcfIGgHYLkqPIRD/OmsPIzvTv5GhFS44sQ4LTDk4HAYRZ1G
2+s4mPg/T+meyG63ESIRABJE8iOgnVMSRvETj9pUtu90yxzYj4LXkpvdQDDzDCV3
EOPo4zwXAYARWj8BDt3kjnYWs3F68s2m2hpyXIMKVHuoT2DgThet7NbNKA/saPg6
i6rKzC4p0bGh6yZ3MhaRUljNWtL++SQ9nOyJJMdMpRU4VkDE4YuBBHv5sOunDGD9
J/Aco5+hWRTUD1Id3R4jbx8WbaB08A9n7ZfUtBWWW1zj1IcOVlW+OX2QrAiR2Du5
KbU64olE+zSWWn1blzcVzKvmwcL5Ju/5uOWJJHW0zgsWlzERZjkguxRlQoaC/gxn
OeUdRQ4dTtEbcLvrkjAS+02Qk+6CsMcm/+a74drnP1vtt7+CiDOSJXG57aclLLCP
LnQ54brHYUEosFSPCg+rNIA7MxEkADJZPKAY/FJValZjJq+eSc1fXSYywr+vfRJV
z14EYBFbn19jiWDZfXwplLCOfB9DifgOyDLuRUj4AR/URr1fJwCAFvFFaKK2cEu4
FJ2MwMkX6hQZRLxCxnTGM4ave1u29ZGlJI30poSzV6xvxWNhDdt6l5+9hrWVEBkN
atXAK5glx1uwSpPIuN58tezqpCZmDg1b6Ao5YO9T4Fjl4Q5cnRAbFJBVDYbNJeLF
jpKvJCabR5xrRtt3L0KxGs47WWRmgor3EoFikBcjP6aGEtgfuxkwy/ormnchO5Ot
LPs6Ei6JYpNty/xXSVUaEZtGKbpYtmmp0f2tD65jyrz8JvDIIHMuYn1zNu2fv+EE
56ZBG7vmCuOHgcsYr1PMgEaVaHfxMYb3EdJLSaw0OkBjF3XuFhxL8GHvasWKM0je
Rpp8UE+jR1li5PZi1pDQ5Ju2PjoIBv+Stmn0RP1s27kcItCEVV2gJVVuxz4Qtxew
NGGNJ3xbr5yjGiN2r1BBu85Jwaz6FHhB2gRTsqNeEmyVOgtP+pxCFh90VCUpf8/p
M0yawO2fSFffn5eJAziv1WjCU1RfJnVTS/2mlK/Hhk5uJKSwoatExnw2obHwJTmW
gx9ebJHqSlTX1OBAdBNdEf6kSyTRvCBgMCgxLjShAucGfX9SVMChO+P1mB1+gETC
vQC6eshNeRZCEkJjVOgIrlQEipD8cmhY3EmZAgd0rIWuXLoESRWYbW9UKr9liJh9
Ecifgvnjq8ZrTnICT11Dpealo5smDiCdgAXT6h5RStw6SlaRy0m2ti+B11JJAae/
KsBu1sKuZRCM+g7RynFmGB1z6uqYdnLABooh3ceBOwfdYspkyGGWl0Nysju1Ib8e
UriBXwMWSCQRI/bR/Ei9lE0ptmv9rf8G/A7f8Sw5ykabp1XAXS4z6qs+4EEXLyGf
k5MGnbdxRb8Gje+dD4Tw+OjWMpZl9+4F/6Aqq0d2s82O9e5MpGmF1GqQRW5EWFdE
7GHK6eLF7J6m9sR11St6GSeCVjy0211NPIf6mLofO+P9EEquRR7XJdadCOvHZMXc
eltXPJsFB8daSrAKTvzq75vNYFwgiiP3M0tEjRYvj9gXSvPWqigXqZG7XMgEUqKV
N4q2sea6oQjs+BlCzEB9MRI2rqESG5hEiyB74DpX9+5DEnnZKQ72WMNZOxgmQjnK
ymw0gCQ6ILeGQ7dB9egMTXEm0zPJuQkZiIbEK6iDJjtDOIBDmpu3nA3yrnvpQj2R
jWD6rJcsil6VMjU81lR5DGkLULmTvxYaXecGEDpmyx33h9lUyiDEBDu9s3BTff1a
0+PAKVDnSosLu67zEGdGqDUSpcP6Exbldq5tep2LbKonNumOQOmTCRtj0v559CKd
PScpXyJC2eNIo+P0d0Ekb7NxmVj6uikhD95yf50nr3cr9k/SIOFK78ZIPZ/LToCO
GTPAIXsHgmLTIep3Inbrh2kQEoA+IAE02VbSSH37xcodbiVpxDt0ZA83/UwwtcPo
3pu3YcboscfVVCZu001hqaXDGPIMHVfzxdI1Towes1tjaL6uIxRBmBSDpBJn8Wxl
r1hPlvuK8vFxlsXvLteOUrY1ouh1DgxAQliWGFp16v4QPQBOjhlvitZg+rriFdcZ
GA9i9eUeVI0rHvC7eUt+AuY62ezEVMH+bzjcbRXkimLsCOJDQTqqsDDjUQDend/J
APnXyqOmXJnI4l4oXTDx5MGR0V+AhYntzCZIdJOxHPWw18To7rhpr+PXomzhpNP/
d8GVoHEZkva1ZeiCqywK0QTkoIg8gSg1iCNty6jVrZ7y3qIfovv2gAkbcvuXlsJs
YQDZ9VL5z/tZNorILjp5TP3c7tSkJDeh+ZDtd/WfZRRaBVIzSNHUrFDC5FCpsW61
0/iy2esHbjCqZvktfZ9VcHvxH6P00ZnPEmQYUCuJhr24NSLEJuXTlWOmZbmp+mzh
oKMVkZj/XPD/Ar5jlKLYzgrdnhvE4SN7qa3suhfWY+cgNNSiz6HBcC7aX94SuZhT
FtgduJ3r8g0ntezYcO1l/FWYRht1XjtGIJvfQPkF2boZ2gDW+m025VAHfwZ0yqjM
yEHPBJClmrfpiuDcQF+2cMw7wNf+gl8+x43gg4UpShZszkgI5vt8D6xaWXleenfo
5YPd5zW4ROapb3Yh/psh5Kp2RjrzW6EvgMAmIknKNUPgBDvORIs3WRHUNP247mhF
S1yeTYDJMwfXffX2qMJ76CjamXf1GlcF+loBTne68qJfqwqgOQMnXdkM666vWiIx
wdlyfnrAmSTXewZp+/XbTNhLDIM8jYMYfXDof3tI0Uf8g4yqnlgMlqpze0EsbjX7
OQhbfpFqiVJ0WswnlLBvuBSJsMhbdh0XI7COfb8Y/+mflvbiUZjm2hWtGY6SaGYX
WxgtHyRr0P0gzEduIRu6JxRKj5mpj1DkXjZkx3PMDOKkzSpuE68/8U1A/3aFSZC5
qAxnMMGQKn0v/WLHTW7Ve8WbKAqHxg5+6vd6WxWafuoWa5WrP7w3BmiGKTZ/VTpl
PergMauUU2CaT+vAPCdZz510o+jZ4hqY+0EI7d+RJh1QKOuuQ4i+l4eJQE/JsqW7
ccPyjcZv/zP1dsDT0M0eHr18Ncphkl4IbGcHeCeblYIs6liK51lVc5BNplO74Uok
i/Rv9fE6j306faSLIgeMseqjvy8LqOzuPOVtuxCQZ4NO8KZ4l5AseNFpscBsKtCf
c96RGoaTZKSkJD/J8xCZcUVcUHqo4+vg5gl0cca9gTEypyzXYgynXm2L6dXmEmXH
cg1WD1nEcVsUwFg/8DjcKCgY6PMQH/aTBqOJ+UUtK855pZ1XeJj25JZubxv8Mda1
xb/cSV8CuGAVsNlGNPcku3URvHXIvWYou/bYHQwTL6DPAkO7it3EwEbNl+EQS0Nm
jYCnWcoiGZniPNkx9N72EAHubfcTkDU9u/fjS5cGCchy4w72q7td5NyqJdK7/1ln
9Dke606FPsNyD4+bEVTsqQVBi3AeAi2OGf6l3crw7mI46pOcg5vXB0vMvCKPgYV5
38eFaDwDJT4Kq9HtNqlVrlc4NgJ0GzBOP4GfYfwyyIVrwKg8YGxtmkKGin66b7pj
OjJ6D+0G+Jyju80oA0sMzAelCYjwmJYWS5Oq0e0F4Kcm7BMvwE4acCRbRa9NWjv/
GACyJtyqVZ3tmFa/FHPI3i9B81hK0QwOQEM+LnJgIfQzW6lyzYuIGqCCj8MfcFvN
aXRd18HRObwAOgV0Oa0wwim0e34GOWdiAqOAGsVypKIch6MzsDZdUyHvJEX97Dj3
Hjq9/wPXPVqLk7CGMMkESZUuMRUyET62YGbgIedt++DEd3hPtc2s4IIIwXmTg2Iy
uZTj1uXbcUugNZRKf91umD8mi4WXGslgm2PhQYUeZd8EZUQRPc/yXXkTUKMijE5J
H9GnRz/Md4PM1j1Cnzea3d1kclmZYuRLKSgGC4+LzzkJTr0HlC1MMsZS6aSModei
3LzgGl+OLeyeDK9JEMr32VurwsKIqhu+/sodbQX11VUDzmXIAkEeGIWWFQ2nhQWR
bOmXBaS6GAB+z+8HyPsyNDgr1vsELw7E2gBCVfNZTzXTJQpu9/gqwhDRqGf1J3GU
LJivzlOjsdUbj7om+Fwx//wmoFhC3xVNeCvANYbwXYiRNdJY/iqf07c4LiSCeWni
4UV4bC1/T51JXdT4K73LsDCk+1Jpxv8FukiO+gulvSR98Az9KhLClkxp7Y55P1PA
y27B6aI2yav1wD/bJd8E4RMiYbeqawsdasImQriBprE2QQWjJSd5bYFiqQeWrt5z
X+unz8t2nUbYlWGZCfCHFB60YVaYNr6ICefyUv5LDAE+fnkA5TWVa/+WglF7Y9jT
6DaliZb8FfbdIrU96zbEqZ4M+s4s6mbWs4nxLKtYgRiZXddjd3aOeTI0gksuH97Q
5cqk6+gU+mO964A+iD8QnfASUThB8sG60TfPVT9OZbc7n939lb3tASzeN3OgDqpW
MhCfvC8Qr3ZIkF0FGZ0wKEWLKffzdbbspixqRxJPBd3MylgZ86gZ9EKdH67YmnXM
wftnHL3bHyZaul/BnXTXemxoVNMAknQmYXAR0nqJo83Pcwb0xedV6KzPKf47kFRh
9ivusj9yXJVtR8PI6h+aXQkijEEPr0doSRwpPNSwlCl6EMIlgX1guvE6ZL2A/G8I
x8JloBD2TNdBrO6AYhW96okFKw1aUf0Ov0zBba1EWxpZVFA9wPJt6o+DzQu446gZ
JkSBe9OCc5wiMOu6t+Q9ka3XkTIwry1kwNmqP3EhuMECBKQk0m5xg7fgJ86+I2/l
bPsfUcigtloxQ5BV1lET4dYMDfzmIrFFEUVOS0M9P1Fl/PjOMBvbZWxc+Vx52D2Y
6HtZRyv023xFB4/yIQ5KcJ8HdljSs3qYKLdRcbcRuD5jTFS49RdGB4debNmPNFM6
NImushktBf7nqxa7SvIuZuImGTyT3SCLdYxrrv6Io3eEcP/ku2xsgcRpXiu5ji65
iDnTIqcpGkMxu9BauNTPZeV0gFzXSR3ccFh5sHi0EZ6B0kQBHmWGVp9FUxo3TocW
yCVprWcymP0PGtcwoRslOUwRl9+PucBxn9+gXMpjHwg0Y+cFB0eHxwXgnNQYTJZs
NTLaPhTVeWGUUuzvVJHCtuBydXJolVtONuedTc4EDhxoidy2rTOs+9P7pAm2oGZi
17eteMPLagYmjB4noj6kLCFUwMO/zcLJL8rEtApTwAo7VsuOoIGOia6Z4EUtdusv
TfJcgucmkRWu2Z8IJjewsGgaDmmWmvstz0ic4roXCLSgjQ2/k+2KELg5/cnjhQ1V
u9RH5VxBjx4o/9BljyNAP4T0JJ7SMsHqZD+OkA/jZI+6ikoNnkt4fMJ9umyY3YtI
g3JRjgUHWAu5adnUxsCkq8Ynai2aWP4c+7ANdBVrWHHE/8Dqb4R/Ng0FpSMyKHdi
ixoMLIUgtpP6WK/wQBecStpC/9A1vCx0wTSp4hfytHsgJpaEUH4YuWvIGvItD6ZZ
1YXpmPGE6tLoE4HPYsItOsfP0TdckKyWHPxEhASnQz7hXRLnMNr7bCTSVo++FYjb
BQqE1zuZjMJ44NczZcKOIdKXOacbHuBuzfwgrfqLNdHmSonoAOTMIWau2fHh0rVR
E6cG7JdCBL4I7iXeuNR5NL3xGRjstpy3dIz1mPP2fAyQeC3jeRr4PUogVNUmLsx8
dVN6+RKZwglAReFpOqbLygMA/8+c9Lifn378ZbtCua198mbtV+F04xVvoQ0341+M
SlFn8fW+Nj0TmJ1Uba115C2bIcVnQqOFcbkPNDmQy4weSXk2eW8tYNoBstT5iba3
yoHlD0X3PYwGWDYkyLCJKPPW2+ozqlmDS4ABQyRo5igp7HohvlvPBcdmbWK8oPih
5bkX8eu5iqel2T4gchZg5zrvtOAWixSZZSrGDeg1F4AMzMGScGh672Kdif5fuMhF
SUryc++3CNCtlrKzi+goPIxLWgMk+blVipZaGI+ZfaqtbA+DSnpa/kE4oiJnQEur
XJYM3anvnWurGChN31oVeYsO38U0vv9RL4Aso2wG1IML+7N+uKJR9Zjpxonijr35
yUTWlfER1jAhf5jwb7+HcLQHohI8My1TbCISKNNeHEjxRPGuzdMBj6KETNl0t1dy
xvWOxoil+lXhvMhnAnvQ0gaakAoOkZkU3n+LEJ8QrmbMMnvqmUpDZW1wisY5raOM
xfaqLbUSGFVQUOkWQSZ3zcXjxyfsU/8lCi1Xhey2cSl6NAb5zHM3oDB/vMTcv0hz
TbxXdXUz0EPdRdBBKkzHQF5PpcCyh1UfaaulQp3QFdBl/k2om/EbV6X4GUTClAO9
PuP+vuTtad8SSeRYjD0ByLQ0Awf/0+zLwuA1y4u1sIQSL/7gfTe6pBDTghxDwWsb
lsSiTLxImGGCedD6K6Y1nYV6tRjH96Z4nT9yt+u1WhUochBwFimyVVAzfY6B21eA
XKU2RMAZBkZi8OUkvyjMyFRc8JjFnT25MbwfTM5+4ZK4cNz1y97jYuKxfKjXhrfM
obs9FYNxEknhpaw7/B6aE+FaJ4UQY13H1JzOiVi4kNJxnSWedPP96i2TIoNSKZTU
67bc5XCAQBRQOemDpNtr97lFPrmPLBAuzjSd+6iXNAQx8Vy4MeoOBujbLg7ipsc2
U3H3mbYAbU65n4EwQjVqzf3lHWQgFKSDtqnRGfQvE8+prMZVUXOd6V4jFNvTuiM+
A8yGWmzL8ODeoAHfsmAhUiPPQ1+J8GDhqIYepY6xbHb1qaLTEYLq/vknNtP6Xcgm
5+mR3sx8tKXZQeuJ9iRGONhKWw36MH2FNU+AQHtNBWlRjlpwGWqwQbo9cz9BERoL
cAvF3/8C/oOIzegGS1ZBWaAl5lp6MeRbJOgjz+HFBehf8r/JRoUjTraKK2OneDRb
iZjxR4gPYf00/CldQKvkWBZmDCEWuk08E5j0vLgEihEQMCeFCPSOrTY3+JEj2DLR
n7ZCqfvc8cGQgbtYMK38Mb4mhK6YZXwikWLbzrkY/P9tY8MNFESC9n3DWvBtSTaD
EAKui0/++kKPDQ4OSXZFGNJ3YHOPqXLTs7xspOMQbgQKZShqn8ZWLWGExdGJK+FO
iyRDbvwq76yvngXkwyCBgUMf4M7bkD4i2v4tWcumY8RnFEu54V/Wbp/cw47n5Q0H
hY6SYFi0+dIDSSbncjB12nRcaQAJbzyjY0P4OwI79bg1ZpoOV1tmMqhYJkAVXDbf
wMP0+6Zpe+3bstnGaRewPY09fSgdvN1fUVm10f50j2eSpAtW1S0eGQug6ep8yodx
DCTW5w/mYMi+5ibJbnLtjdozCf7PP1cylz9Bdbn9jqgGUkn2SMmH0geoE04V5At2
Zi1ijmdr/a5tvfDhTypvd+3r3Si9C0hcDqywZ8YjxtpiXy2hlzGaqxI6dnjfYgK8
P0vqfIMzVSJ40LhHwgGO3/y/reHQ7MkhpLbSUbTzu2QDaOrI0OhReaKs6CZINprD
R5HKhy7wqp5uBLL41ysRCRUva+w0hreEDSpk0U4GWQqpiU1BZdBXamxL5yjJXLuM
7bZg59KWrSHqlQx3K9yYyILGmLtpvtTFkhbsahxyiByPZyzVlnqX1Js4iuiiAUJG
owa7R6SofRa/fB6Aeos5wWuY6c80HZ2+v2y0wDmM0vkOcrvpGGOfBXNI6l031M+p
FbZrYEeaKGcwogiwmwNMUNSqaqYG+D4iMW6iBQqrDokQBWfpkCpVMFSE5vkzmwgX
mzcraOPBBrWoxB6nz02tUegqz1jEHqeqwoasSK+fL8ev9PkOix5tdK7KcHCXYMPY
jci7k70Jzsdj6nftrq+q4fvnFpu1QUtGPfgNetxcUZq/8gwKQiBpOptONFskPtxS
de+xMQxnm1Y3x0JdZlUUwDbL+xFROrBAOlzBs11GjZ0ky9mpy3oyXko1F3NRXdYN
0PYn2NLN99iaBh2zxLnUF4Yl0BoEPXjJK9CA4FaToJnSuYVjhh96cmdwhUINk1l1
amw4pTKUcMQLEVlBBUgupqKDcovFYole4LVSiwj7GE6UeVt/K+IFRLQpUIPy1tpY
CkBWGvldq/cNbMVRI/2LP3N0lfw+1Surd3hjRa6CNx6DaZLWfpm5FeTgJC4Z1FO4
eeSHs/BlP8BpArk3MtKbzo5iKb67ky0d7V0+5nVHAf2uKhERrZQCJzcCz30mMNt0
9BP8j4ERmtO8l4s55oOLV+B5TrzuINXzpdXKliRMiwxuJ1g1BUS7TEt15Y/XUHsM
FDoxV5nGTHIbVcjqMXfJj+xO6rR/xZLRtvlmPaWquutyPfFIr3ICKEMuygRNeSZx
Bw0M+98mNYpvxGM7JowzglbmTcUQrM91QBx4U4t0EpbwLnpYaDXN/FZVmTuKr3tV
T8l61kN87mhIPE9aRhsklV+LYg/b4vZH8e/+tOyAdMwjPJF3vAZK8l89ai4OUokF
C8dvCYuNWkAgXw8qVYZtKTDf1wsNWtlZHwlU0lMoQYmBmTer7c6Mj51QjQJYPJnR
QSoZMeoNt5YzzBWQY68UkzZBrcxfOVYlaGD7ZCRAOqWkzaof89P0j37jOrQwfXXg
bl7+qJhDawxHKSOagRP/nEgWuVIZ9TOnmhIRmt0MnNVV80In3x0zq5VenA6wxyU6
jCYyjOajebu9SrkC1mS5Fv8b+7CT8u7gfuhxx9XHGlUvrx23hTxjCe18yRKZhu/Y
MJaeL4ulWRZE3HAxtn3drIaANxnMREvTeNY/uhHH90+nQoh5kzWjeoVBQ1Tddb3K
6B1EXU85l1X+i4J5TG5RspbzhlrI3tFwqu7p2uBJMSBt+TPUIwf3aIAleQHjrw2g
Qbh6vR2z6dhKASvXh7mPjfYcvYAlmW41OwZ7QcbJxXLaWfafIq/Ao1cxDGKhJStt
conQmKvAGxey1wRmNKFAYRBUrA8VYgDTDZuYVd6DIJuh2L/XEqGlJv3xs8m5GqwS
zfWeqWD7qe9v/h3OXbaY6+66x9lKqDhFQgp2pRmVMj4WjkJS2o00RjeyZ2UUn0qu
zYXnH3Zgj5TUPiENP4Xc2jGNUa5cAagfJqNEycs5etHwleFIXCgFsJhkibfF29+g
3adUizL6Sqj9dTZlzFIk6qj0mr5he3maHB0NqQSYrZHOj+vtl/YbuJmTBNBHTeM7
QEbJYmoq7oFEZZGajfJ5zNuwMR2JxkRnuD5vOJZ/kM2X4HKPohLDclOBBIzdf+dz
Ba4V7hFbzIBoqM1r3rk2m8Dr714AZpx3B04ZTj8yMqbDpaAdwkcAjpVMg7Z8L54A
9GRyaMPDStVjfazETmvMMMeZl5bYhsSlCJHW6rb6oK/Icrh8b9aDvGE/exNhNDzv
jLHBIauDmIJsMB9fQMufwMRaAOqgq69lPajvd4No6c9kvBl6u4cT93/hq5WXej6b
iYk356DR6/Rzm475QP/mskz8zAMXjx6vCb9ejDC7yDNmcYB56CEbh1gU6bNZGvA1
by01Xv2KYCmbT2gizyblahwXTPsrJtZOcFtzdDSkJvnp90+NzuQ9omXvvZAbHNoJ
lwDu7yjwrmHJTk7yLq46xr6Lms9nTXh/39GhxwzXx6xOeNCz5hITDfLb0M1GBYi/
+4UC0IMld9jb/BTpWKsQj0LdpHWUMrsyg/j4TAwkTGNmXpJ7i4p/oP9Xcp1L1gcW
uaVZkU6YxVNd/YUtxKByc80wRhpXhIgKYtkJARIeERvDMuPz1MZzOLoa4rjM9q+G
kvlmcuCqD9WI04IShaddeIKO+2edQ9Xh4NDTuYLwMgUcGdMktvqoqLVZaVhgIt+r
9Jxr4OeSbFF3PkXF8bbqigbbPIrCk9iOcnKMoBIk1NInZKR7H3Rf0Uq94tP1pq9O
mq4j8PjVrkxgkL1qBtaj0P9IH6x0Q6MRU69PRro3NYMG+jGmwfDtlq461Nf661zP
QI/vkv0psFLNqWw7V03ITI8YCVHHuNYn7HErhe2BZBv2hJZ1bUAYzSsc4f6+TLhe
Mj+N57C+6Myc0E5XLLaEPp9JGyucr44Ne5wcAVKceMJIHUP/Cxfrcb0oyIY6cWq6
jo41XbZ83AAHV1sxuQbITXs5PfnSx11Oo5JBWsSrWeNaZHOzrBJPsNhPS50BzDgR
k45a5XbTyif8f1SBfXJ30aTFvTTHG1bxfzLdSQ6exZzCroowbYXf0XFTrafrB8rZ
ywLuC3RB0rHMV32JkpiXXwT9E/B2mwrp+0YgeskmhcfM6jQxT1IV3BQXPTSqKC1/
rFZ9fSVPqpJqTdxMIvPcGd2+1SKjvQxi+YUiG1RoKyFwOKg27+Om7G3ENeSqfHWx
b8x0keQ0GClMsoSxUAxCPqblCsSVBR7AcYRugeWedyldMxwTh/B2goUO3OBsIXBt
ed4uVOTxXQb1DnaI9YLbtpB3NDHGDzkiZMjh7LiG11+iwBSbtWtf9ltY04T3Tc/V
Enc/sn4RjEbhlullexUQ8ywg+vgVb1+nxixZmeFNfdy+ZfFgeQ9qqS4SZwrDnpkZ
DgHcEwdaduskwKsFxO+2t17ZwZNe61Wbv97sVB4qN4aaMyPyOjhk4TKDqEfjRc4F
KcGytxh87VtAB0fUV/Jq+2Xj1ldLzAgrqy31VdO3YgJuWjaHRuYSifR9eCdUGC0r
r93yWQpdHiLTfHt3yF/DcsEil/OqSw2OW3YRxg7K9Rq79uGJ1Lq/eGI2g2iRkm8p
S74TjxHBt3NJZ6IQ8OL9d3+8U5rf/OBPt6PwEsDs2j0mnBZ+Ot3ifN9YPWj/AUI6
n4MIwwqvYJLtBFze1VcdMlpNrcIhZVqxX74iweVoh+VISAXe/mYSbOfnGwdDCg0c
jDm67aHXViou72mrPrvxatQu0NlbSplbmQhFNsuMbqwHsfa78z0xR8oXnID0jdod
hA/iiVxfSvqR+qeB4hLqD9i4p42WtWhieKqg3oVysCcP6Eab+RWvO3cONhCVVr37
qadD9kmd7uHdIhYuov/NJ2lznH/BM5GjDkbqgy2zzxk+U/xKCDPJNNGKAUiwnFWg
LOrwdKTy5NaqnIxA/6pdunTL4yorN6j+boXWUnuSYB1WM20eCZJeogMREvDfbXJJ
0zPvNI4x1rHge8FM+29MStfaAZFQCEeLXcag6WsUqVqgv5i2dNlt8t+rSxJCijA0
Az2qUV4SEev2ukc4S3ApGFhPDrJkRKoazefUddGSbsNkeLZjMfGInRMhOnvqM28S
x7uQ4n5KUPKL7sZOf5oho9Ddec1euPJEInxCQuf+q3CQbcprlGd6IVm8q5qu6gGC
+GChTCsoypukfG33gOoRqQW2ZL7jdrNnCN+lSDyBD1ULUZx9rhxx3MEeYadoxgjm
/k99yWUo3s5O+6WpRwaFLq1pECt4C1rrWpxp3CCZw16NQ7vafHAJEhnD6RdYkAmk
/snx3D0Eur1czqfFJWIx24JdLks0mCakQ9qekxzIfqXsgF68ZGnFrQiaD54KdQO9
Z048Jyh2K/7X2WDa3b59Jyhp1Px37cRJlmKZgA3M1VUks9sSc/rSqZmqUMen2wBB
NSeBI6XWSo9UiK4bEqQ3kyOy1gPC3C8BuqME3ZP8lhRDf/GtT2ms2v66USLq1jPt
crK0NpikDD93Xm+sdD06GdpUIa4bi6fsHk6YZOz+mltlcFvmQotf5B0M5R0a/vVz
C8kSGelXvgjjjQqX+esEiVoJj2aN+EUQ0U71crGdZjIpztAWZv5QG7QOtoHzWEd8
gqWcMHRj0suQ3Xx5/MouPPBdH/2RkTM8JTGtUiuZUeh7fKK23vdiIUoVcQMpBqMh
71LrC64OSxFm2kLrk4BKEAKBxsMI7ERPhVx+n5aToOPFUvLTuIogPO7CNTVMQsnv
rawMwl48cTM6L65EwzoGhh4z2GRAetdtB7O36Nm6kh+LicEecVDv0BubgDTEDMmD
Z+7wGqoC2e2mRMOs9uSa30S+oXb+2h70G93hIhE/w/AhZEybNszl0hdShvYMVPuh
0RuA1BHfkgx3HwW9z8+8kgfCyjG6wyHWj8dDv5kjO4b/fkkOazQcn6EWgBXI/c9k
DGQSqIa3GB0stC5JZYlwVlJ+35Ts9xGIUrArXAcY+fPPvr3pES9yABvSAAEyE6z2
TgH6OYhO/2TwcSjRoNCzBpLYFr62u2mrY2bc0lTAy7f+CKuOTYxcQbVYw4qo7WlF
J27/oLS00mCYc8edmYaqg/NhMJ8z06WZ0dv1xuZlijM3nNW3XmXKBGg99g3d2B7A
2qu8gviB/KoFN6L4sBKRI0d9s50pzfQ0t4EOzUq1qpjVVGPn+6cLRMsc4YxxRduH
/xvUD5Z4NjXcBxsO6+Zg59weNyRpI1DEcdnSraXZm1X7nqYab3jzktAkWVC3eZu+
ADdeX1NmeuCkSiQKSK4wEvDHEPa4MHfyQc5W7ouFp0VhTEuPwZG5+iZCz7/P8db7
ojPUWH3R+mj6txEbOPjKWAmNZWi1WbS5TGI109IH6LI5SBuIzg6be+S2X06U1lrE
WbMETjfceBEqFHp9/rcfinnb1B03/Vjs6gYQl5M6X5JC+UGEnRz0Fu6r/Eg517Ll
uGBPt9juPdzxdNlFMgO87K0/NiahD8yIIawJJIi17TujkwmcSUn7kZWfH8YyAPRz
PiAFrOpqOcKUbEBJk2/6q0fNKT1DWEBm7yckUmNwfIY36tVeTsNyoNTofKoIN+sn
rH/1ln6B+PnVzD/AN34abQEISUOK6rASZH12uGVRK8qcYjnj6+EXk2vNhKRGPonw
AgmmMHFIS9wGIqHIeG9MQ5QSrCm33LqJd4CuFCl2TukasjdGoXiKcOpwoo71HxSK
HbU3h/weQpn+TNgVZ/HOgUyaVuCJUMXoPSwqT9KHfBfWq//+rUvfmEYj5sH0H8RQ
lSagjoQWoXDWGwTg/K0pnx5WdzukX9LfvpNe98AzDdyb04wyjiTOYAuHiU6Oe6T0
IJIDybJSQk6sQ9lOYbQkQjX3vGuLesv8YpyyanipQKTJgambW5W5juqdHjtGQIkq
OGf38PKRfvXX1L+O36539gmWOQipLT5N92Yt9jLjXSUQ5Yq/sW3fZZIsu2MigIuQ
H1R09hxqEPO5RMqEr7PXL06CYtgi9xlPMgfqKDxFA1oy0a27dxt2uj/iuEoCmYmx
f1DI7FlUL4qkxqS3EKhbWP5c5fAFej7YFRb8r14Te3Oyw0bCXZhBbvMb7sPOm+Sm
RLlVcZFenYXBRYEz1RYTWY2Uzf91+sTNz/+vvuigcLJyXbLsdTsKcEv2aPtCqf84
Oi5PlbhAUXvSHpPknnFLw/c7M93k/qy2P32TnJboD+cNOWBzj02tJusDgAFE4Jtg
DNvamkmv1mGcyzG5hcV8LEsBGyur+IdANh1hlAGcfesMqqmksU4QsPKMEl1SD41n
yLNF8CEFoUYF0S+iwJG8Mf5nTShjwHM7guydrvbQMa0bfsc6gBl3i+C17QmFfXBB
T7y2vzaNTiokhHR3cyMsV0RcyTLBkbx9tAqvCkOFLH+PDQAuf4dg7Hmc3sO8f9TW
/NtPyyJ1fXq7fT/EeoDEpoqvBQQJG3NYJ4C9KMXrHEjXbFRXXhSps/oylijrrH4r
sWrnlpYf6oiuuvE1JAgOMjQRepHZoTcI0nBLy5BFWjKAYc0wsOdFBVr3ACDGZ6B+
dj8yVtuRXHRu3v280dDpeYw8BzdpoODkwpQaXnlrg14L4tUDX8bYYxFh0CzeScCa
AmH+mc5b8RxZ/5JcC4r2xmHDboJAsm7eBPU/NF+d1KXyfPZOzBpfZwYu5QkTFtQM
7DiQr4Zs9tWeISf5uXQee2e1idTCoMK+VAXw37QLQyq5ZcgJc97OW8fvAfawUlWc
i48LtO92j6AigU18hNtw0aietBaLwNMVcenkyApOoZG5pG8AR51km8+oGkzYqlSy
1TW8fgT2v9EwyndYz2NnkKmi548CGUadjnOxC5KSHnt2caBEoP7T3GInmxDx8WEU
lJXxoSeaqqGddG9we5fJ3mUVf0vRgHqABwxnJxEKGl2CwkPaPa/rlUZh0SF3fxgl
ZDY2c1Lz3ED6Ise+hvG3EkoA9TKtvuRgVCl1roST+ai3v3HZBnx2Cnl+ZIW9XHok
CIk9/RuCgGp+1XOaPGiZ5m3kP+EOjlOFjYnvgEp3Tq5fl0JnAqDr6EfXta+qrlSu
eRKXQNs1/IUAn7vXsvq/eBCYtxHqmTFGTTjMQ+wO5SckhzWHqpaYgN9kBodR7N6K
IcfOSQn5WCfIl00eo3kOfDAR6gJYHPKUxDP/HzkZUfwlofdJUcLhUNyp8pu28pQG
d/gs1LadQ5iwf9WJUeGO9LS6q7NCTntOKe0+a/Pvjj5GfDCzNe0/nU0zt6dgTm7J
RQKi94lqzaszCnUgogvBoTlgxkIiJaIgHR++jXy7r+apo81QBVnJylggeFLe/WPS
O/HCMHVu182ZSkTZ4et/Td5b4fpJtg7eBqiPOrEbFBk3jNd1vIkmVgXKf55uujOD
q7f6uYTg56ICHJQ2yCRggXy4U8Mcbm1TGSkUKHknWgQ/C+LcnHcxcUcBKqTrUOO0
AYaIPxHuh6zGs5o/toMxW4+NA5we9MK199vVoCqe40gI0gRtMXiYY53se8dRGCCq
6brSYUiU6jGHqcEc5u5ruqwLSJDXvWpeeYLoVxXJLBHAPk79+1HH2PRmtxxWjFzL
oWKs4OCjTXzQSQ6G2I54rwCNDg8+jWtPTTK43YdPBXv51VSICXZqoCmgc43Wia+O
MKR8VR3WrhB5E33RBj2xlydbNzesAsMN1UNgPXsFrTYD3lUD/y1sEaM1wrKIvGii
ZoHGM++C77Mw/Q0RABPL0PZxsTELFar743+NNRgEZLxqJWTaDhmZwRvwzdLIK5dU
gfnyd9mNC117Tm5NGAuXAFSCr8Rvhc/bDwzSRYuQ1DiUhLMETsCaA1Hxq8/WNMWA
/O82bhW8V2m1G+w3uK7CfMy7+V659KJ4IVD20xquxxgGNQuJtImDXDNQnVeTQ7FY
D6VuWsLGgeZeQraRcSGBOJ8w1K6hF4gpx6Ljsk3TwfP3O26t4u+NRCcPyBgwOy1t
SYEossRhPe5AvYl2ac73frOIG2857DxctZbgMdHOQYtyxnWS0B5wH5sHEBiZgYpI
DtQcQCzi0HiZixgDzm5iWXeuMQ4rjZWBiK/y/EtFAMb6GBkRYnCwsToAb18WLXYg
3IksXC3hLSnshX32DaBu3NTGCyVkGo/voGRiaixFBkR9ju/+8yrYnJbYCWAJJJHf
x0whhNo4cPLjZAFlhgf8UhEUy7apcwaWakDEoGXjONMP+L8LbWTbHqQDru21rDaT
CRWcxBuFhUSy8Q/BS+4nmMjH8/LjyvnPpq7oD4htZiLZ+OEDvIn4XT55fulcWwTv
tt1eFNykb/Wqrz40czI//mO7y5kelm+uWvSW2r54ZZ2XmXhYcFm/nQvOuxOfNUpt
mVHlUogNGgu9BDD2iDQfzIAzRyyY3R+5VRofzDneuUfssDJtgGZ/FdWMbw53QHJK
SvOQdmRktHG3eX12IwAL9sjdCWts+OZ3OzokrNcM3AAyf71OqqoaJLFS1L3U9jKr
qN+RaT26BbNoom++eKXFH9H6hhTy51baCasU1QdISzPasnKZ5vP9DZ4ZRvvMd8Gv
VyNhAhcJiJTUEn1IxASlEQyAfamtxz5EK9g6E6g2YRwmfxVKYRohZI+NO1jHablh
u+I4gojSGXm2pMMDHpSsV3PQAIdLe8ntUTw88J7P/D5rXeKFTUZyo8TObKClgFGO
H5+D7R7ZvhS0Y0vP81lOd6sXtHAVnnf7g/+0wO7/DMl7UIEXa37Jcl+ScJXPcx8q
OUTNQunUY3PYuKUG0fWOgOtpwjgOuBW7qzwy3VQdZOMa/Li279rDwxKqbI6cicOp
g2ZTsIZfRrR7qU2vcm6Kgpb7lD74sPMnt8eZma4Lg5vv9FWhsIe+CGeom3zsWSLn
mlynfi0W0jKxHLbXuIkpyDMrNNDc1MMP8hwITpZdbsvdbQXyJDX5y6/j3KMjpv4A
nPZMZ20XOLJtx0S6kLDMTXNb+jxOVBomD7zaCfx0dcSAiFSWIxLEMAHLm67c/QXm
nuLWewMZpURlJSHjBgUg2ms7FhKzwxtzpgy5pjLE63fMsveaGMOzhRy7wmFfJpeo
eA2kfBM9cp9Gauk39awcZQA5xTBvs+XPmcyg3/Hevlxzr+m+0lIRmwkjXxnjL80h
5G1+wOPSmEoK8SWmXMtZhdnQLk0xGlVxYMSQPH2JHWo5RyHng8zpSLD+HjE8tQBT
uoD6t+wIVxeje/om4f5WRthwc5J/caacPgbOxyhOLrPFv3KwwhOO1bHYMw6vlCpN
8JzqF29s7M01BB8pE7PkvnRCTJuZHB/l0iy3L70IVx+tRpefd0L4puHFTNh+h4p4
Dxpc3HL6pPHXjP0nOkQ1ZgxeFy6m/ADBFKeXc2C7TLGF2XJEF73gXATY1PdxNIm+
tKQcUGh6F4VCRq8+fKlclY62CBDFwi7cPg9SnzXpkQCYFR4XzpP0PLjYCA/6hYYE
UjhaUyM360XwdTh87VtuCTcOf/QUWq9Av8PyuG4+is4ogyPDkq9i7VfmPzVhJiSo
dky9AWhKa6i2N4TJ0IFKsy/QZRJ32iWt41KI4T40k+b4kfWPeBBPbtoHgB2KmlSi
un5Eaxj8SIkDPPAzj9nJi6Y04zbki4gXjcIPzwlv1FVlq5SaBYhel69TKRdP4PMx
CkNCDgQYrBBZxlc7HfEW89o7g8+tk2mcOXj77p1/1Fqtu6jeinj3YqL5ZX1keHsk
9Yr7Dzodd8MMZOmEsO7CSnh5QdLyAv/pRUcILjM7oyH2Ntb82W7i5gm14G84jlfG
oDkfU5Frym1foCXrtW/UJ/XC+oOwi1Dg+fcab1b0ovUoqwT7Sc01VHGA5Ugi1IDc
emuGoctMUTlKCUC4PwKFXWD4G8rEaOg3VZUYlxmY7HXv648/dghKpXKmHbYxnZic
wbD9gZ8qP8zjX/dm/oGYJhWz4j7Rh4QiNMy9X06/OWAMvlU8GQgoWcIP4/VYPYqm
5rtunY0VOW7dwcbH2cZsHyz5/D3eRw9mVNZhfVpGsqDbYOsHOCjvoMZoY/DObY2M
InWcI5t5z+Kd2j2Q1FNpDeMkbWyhlYjtLyNFwe366S+qeZlZpsCZkT8EG4jIgNLl
YBBD9kJFaBh8af1Ld/yD9OY3vQnrKEmt2e81OdicJUUBQWQEyk83BGm2j/bj5jE7
7M7AjKJFLO8eArtIkkrZkRtgS4rYVOiUGsSsoOrJm5PkBgTqFkx/262sYj56Vixb
H3h4MddfLIqv2zHFTj8OCgehyyIDqClEPuK/f6c3H1bWaHWaNzsvSllbkobAGSNr
CFl/GuRoU99kq8jL27QfudFfLOLos/qAk3psn3uW2bhOPV5rpo4o1ZqJrd6CsJCP
Bg4Bc1tifBlYNaYCBX3yUWOlu3OapD23mmcJKW4wzPhkDXXbGGWDPc5QG8/O98JJ
JkHVXfLApz0V29NTJgH4IDL8Pv7iuweFM9xMz276Vo9mMsam4n/wZNPRsBlyp+3J
15FYicKnnOYgzY4DFvttcbYdvVObzXFC9CSPvpQxmoUi9+4GjhfVd1EHYLzjrZ4+
XC532gHsWZIwcOefl+jHQ72NkWWjs/heuvkaxFmTjTfedKikzgoQZVlh4g1U2UKG
jmUigBV96yVyVNF17y5EPgVydMnL+iW6l7ypC5kjj06f2nBKIOOFUmXfw+HJnfxP
jl+6+amHceAGCP5tO88q65NdbFPfuf/Blu0KDNX8qhOiDc+M0BUaErMcQEazQMFt
2PzLvFdAknqaQW8gwliKeGRVpOkA9x77qMYPkZqCRSpUQeQhzoOsd03JNGHvic5W
9XOqy/Qv95ZrDmoTxihzYMWWS1Yvobkfouw6caQpbmZZVR77rVOEmh0GZ8qvHmaR
ZTDuyGvPmsDHGDQ3J6N5Tln7tLRNsu73cERYEBTVrEmcWg0tx2hS7cnFflcXmwZ/
BgRyrE4asZq2qrdcuNj80CZ6HuzAf5VTj9ml7IBG2ByZfAbmlS9Sc1YG6HW5VcyZ
mBvKR8wOMXjnXE23mIunGFddjPgtG5U+wAQMeaGt0eeGjOH0JmxpwUPlz6mu63EZ
WAfkjaoOGOUa1r/7gGXmRETY3YxmHvgGbASQ/mAFJFVvpL1TKjear4SwKVB8zO8X
R82xwgiPp0PWCRAvv4PYiN5t92kZmVrJSK4hM1Tkrwei25tVP7tA1rs/c915Mf7K
jsj0vXBK/ltX4ujwGXSwhhI8pXH66kv1RO940LOhkb+AZp1dqbwT6UeP1QAEsD9D
5NK4ZaZNJFwE12CIiMFQDme8lhldT4TFXS8cxyR9VpX0oQebirI/Qipv+5hBFD0G
WalcyBcWPoD6IO80wR/QEw6yHsDmrTGsjLa7poT7faWQmjbqQlneov+CS+ztlJ1a
IpvEchqBM2HIZoPPkpDWsY0WIFPp0MOKL2nW5EgN4jE7bl9HQVp0qY39DiQFN7mK
3gQnht6AkEt5FMz+Pyx3WSTKvNf9+J5K2qn4pJddq/HihwrRGlU0eMDe+Bc0phXB
9gpyl6GXAIprjR/ZiQiebI7k4yMEIac14JyVcZDZBaQMK3tyWoJ8I1O+/acuxYGG
eyUw0lKy6Q0nP/HIjpuAIWbROMzhdmr+axykmdeo0iXatkNiSyCqQLwSX/fDMM13
m7KUI4FXdExy6YZeJksKFxDY6nvG89eLifttl8ZSw1u+uNLiBcdS66nvgp55Msjp
er5d6NcX1VMCRF8ZFT+0OzPS5C0EFRGXeQWBgYdFI9VcBJj8efJ0lKF9ykmXA1AF
82O9PC6WaxKv2IHolFV6fwL4VtxQklnuMp8f7uaUxaCrNbRAXuEZKbieFCJqsO2Z
YVwA08Fy8W5qQ51BvXdDOreu5fUkazDmza3RpB9fXAh93GlN2JAIZOnSjEgmH5LF
GCGybeBZQ7Y3y6Dvz4hRuO2U54y3TL3QVpQKqdv74gHevFQ7lCna2iRHm31A+yhZ
jllR7F2WtymqIuTUBWKfUSStrBUtPUlYwUeqY+/FnyJojYDk4aiwhCadSi7Z67BW
FFNXGC3hqsAyNp9ey+qzn+rxdiFeh/ENQJkm/n5aoDyRe2lS3fynIeKqCaTwRhgR
uLXwEZdtMRc+5BOTuIL08y0XxEpAOWBk724B+PCdApGRYMKZFEbot9swYuKKBpCX
JugsvgIxLk22FMyG8mTbPvliUBbcwZxk5KWcxb3yhbGOp9yokwJaVFzBw4F+1s9S
Jf2+4HjC19Ptuyt1N4L/MPyU0yRZOgypk9wFhI33S+9hjYzT4BsAVMYOp6FcASf/
m0ZOxsp0NZ8auQvf6GqSEeR1/1NVZDFURS1d1LW20LgYTMhkvC8z/FOEihdZG15j
D/v1ecEBYoVdQgwrWTzDTwbl4rxrfyef63VHBpHz6GWSj1irfOThho/nK6zffV6O
tR7Bd9iUhSqqbDpv/o1GuteQd0T0/YEVDuVsTSkFy4E7l9NZYQQb+z2MxcAsuaKV
mI9AgVarUpXqd7R5uxHtBSqHhXp4iax6xXHSTsc6GX96ZNE+ERD3qcQJmoiJerF8
G+kZghUWtT2SJhx+zJG6dq4gEGuK4gJ0z8KKUM4gXcqovS4/uAXIeQRIFb+OWTJR
vhSgDcC+RHdv2GQA4aexYX+NJcrRgHeoBhJq9eWrLpt3QkyBckPgSHkpyB7NFDAS
U5hBTCgv8nNq0C8DKfR+Oz/ywcA23fsQYvLblJB8OWhbofg+vlDye/0ed98AbA07
aLgpheIP1pcZk7MO6WRChQ3xezSS/xnfcwqdSuYzTP77WF6osTyOPnKEko5S7gFF
Fv0DTA1Es7DCvH7aOgTAh29aX1z2Jqt84IuiTxM7t407FGCtZ+IxMxRA3mKmb/L7
WvmB6PrY6bI56J+1HjE5AtZGu4Fxi22TQilJHKkFedJsZzXaON3bbWnGFQcGA/VC
IYKhOtFVBcWY8ohgBZ7tJr9Dl2LKQCLZNJ+k+OfdAt0c6dB7iJQOzzRbji+kBiZJ
F+KMhN+l2VhzqUZRxxe9nIJT0NxeBz12qROGDOB5gfT6x1IrAxeVNIbhMzYpXTzP
xEx2wstNmaKpeDCQmjsWYg+Gc2o0cPyUELFqMFQrqSs9mW3azA+dYj5M1vR1vq5+
YTTsrkpN5Y92L299e/8uIbJ3Nb/7VhzQw1Ad4QmHqnTEgcmWA8c7q0hX01yedwfX
PcaTJvWmzoMQPv19wL3z76cRrFgRhKOWHleLEdbio/VyhTa6N5WXuZTBFaei1ivk
bron0NNVB3x5yZhL1tkGNVZ2GeJDHf+QizxbAYELtItv9t5Wl9UGLoJ4exgc+Y0U
iyYdHZCF2NZrLxVlkjK/2H5epMtTADxSo9Fetvic1HQTDulJqD+zDnPY4duWMa6A
yF4GXD5CZ7ZEoLryoiDLRLZMknTb40M+L+X5nQvbaeigXUNRDESR8Z513e+71bSg
ty6tq44HeyUyRvV3j1ZsCpM4EgU6pzsdEKLy8zP97NrmwADUWK5w5TD/0giD7KrV
awip+QcazTDIkAWFS3nah1JNtA7mT+UZ5C3k1DzE0/53kGCHLpPT9MR3gQxrMBW8
/R+8K0FsNiF/B8detsvNFGdroVK10kFHi3OKV2sPmBriKwZ3MXleJFkJYhamF81E
X8Vk+XTjqjaNaN2ZSkVbx3lmPFq0dD/RDFB/NjYP/MMU7y0jhEm37flpDlBSvRQQ
tcmx6XQvaXJNwA8IUyhAmV6gebUmf2tzaqKo5iDH7WSfD1EZncbJWrFJSUIYqixs
68DYqh2oV3ki4kEpYvop5MWx4cNVp92MUL4WClaWWLVXWCrhdeB50Kh6wGrj66Q7
IZywrGM/QD1RN6F31XZfbU+q/Wo6rbM+3KJOZTgm0iiMxzbhUeSGYagII1j0CWSI
nXb19yLcFDZLJaG+H3kUitiEkOXXmFgb44IYaOtB+YiBhL0JoQb3BavSVsmcOLUn
FqpsMCO1HgXWLKNndlYCkyiLAZPiQSekdLiG4iobGGtlroKi/jAX+sDq/qXu8oaX
ZARzNuppb/P7/WYjDxCOH2McG3qBouSM0K9gqaB1AFNZpeElt2A9FaoKr9r6t0g7
TBdgrNYcUWVUEE+aJceci2sn2+RanWcXgtlFnMrZy4ad8B3r61sBmjspdEXZo/Kk
NtZm17N1DYzVxC+snZJtY5m4k0/pj/bnlTQXWaLSbezfPZPlVzHoXf43B831eWPr
64e7FKqJsamKrs7oBO2HMU89s56+2EqwmAHNh5lULklpqVMP+oWjAOkeCd3d6aBG
WgIttYVfdhS/IMJb6tabIZEyer6Jpy0b9TjFSgTraVSBxLf5VTqXJJIiKQdjhOMM
cwkfWAX6xAfczLhufsKTN8jDNdbCxd8e5bFMpExUteGrZVHJWDUO0uiDT9KUp5aY
rOgLAv47uQtkMBBqZQ5IvZXWGra9ZuEgPQgLUuePYD27Zqf839f2xNhIEYe3gMU5
fqW/LeUFIEtCRtmkWrHq+MJaCfmHWHbBC8K3J8KTNPzSJ/5F9bT3jCqipX9my3Kd
GiAjyGmWh01osIZQW+2UZoHSvsOwoc7ZHwepZXh8eDEAXJVdg7QsK0w2rl4Ymtt9
9tH4mwK0Gt8mIoYjZHVt83kdeKpxgJJDKm4rMt7X9HLafzaxwYPxYW44ut+a6cel
suuhK2Wau5IJvKRwDQmVDGA0gKOa3CXnOkViwMtmRtwSDFsljqb8GhKdco6t3+XD
+R6VUy6qF1LXPb4RBAlIrCdOmouwR1tmOv++3AwhWrQr3Ckyk5ilpB7HPnur19rH
4kODIO6LYC1uar9Bwzc74bX3+KYkBt+IRvM9KC3Z9Ixksc0cYkxW370n1WwrRgJi
dvwqFQRlc61QhqG/Z64ZDV3+YbxkKNMnPe47dGh7/66mO7yC/PwSoiFuWcVG6u4P
Ijjj/feuAHvfL5JqLlhnoMkYMLGk9jx7iy3fDgVUpDtgjBvVbsm7TZiOLFEpXSGS
HKGrpK2L24/GNZ1J4dS8xpebuqvmVaL3ZJ1BBbQPXOJH6N3rFTO4CcpYLNpxmmXD
d0jfBFxZ+ELvo8EmYRwuvEattqdjscgd1ZMupRSTNJmWwKY/Yc/lfwzFDgkATOf9
kqOFtHeUa3IuZePgWN5IPCAXa+VFnJvxmmvVUdtJgW22i10Q9z0kx221Z0pCKutc
K8K2s/iwV4YevTmQLbBTchvKMbniB68q/lkJfWxLVESaKQ0/Xjq1wfw6ta2PFGv4
nXZjpFDupPvJlq9yv2olBcmvtiJn5eQ2pPu4LFPqtJuJnpMkoCFVYesrPY3fPOOM
35vkZrcrlk+CaH4YcNFCDkZYFgSFnc6tGQvW8LlbEOccJcDw00BuXmFPIj8C7Uan
gMxjQb7yGjzGFf3B8hVVfS0UvvbEuCK89dFu7tcE7pfZVX3Yo7dsD46eJXwb+Uar
aIBis0UGlWx+T7TOgBt3qUIHPFEPXDJ+jba2WTaN2dAO5Kd4N6nbY66KsS3p26Tw
40hesf02JeWAIUfz09BHLTLjnEfWb5uHSB0aIvTb7XyxKcwD6mq3pLkV/8Wowhbv
jFc6GlshszHFN2VJ3yARra+ZttvklNYVTC33HgfZU0/AqeBZUDYADbbTGWoNsOJF
3nB/pH3ar3uqKWd7PAuYETaFW+tQIuoYOQBqR03eJIhF6BtikWx0jhGCTm1lQySM
7BFIMOOyjn6ymPPwpWRctvXOFlZUeofnLq7/xZ1aHYipSROJo/DX/cmY+UxoPBSj
Q7c3GLUyJ+vH1z6LYyg6KBWtFbGXNLjCs/WOoh+1b14T8ijtWQsN3S4eg0zXYj6K
wlcu4IAQz74ciliq4ZXtT/oRneL9akJ+T2FiLaX6Q9UsdQbOqYO74RFGKOhj70fi
4ukncrRTyCb2kz8jUlts/PkS4mrZUF3N3UyRJ4Klmlja+IGjpAFc+jYrGomLAj63
2r30yk9TcP6DcgzCFtCf6rL920dp5X/4cNBYEOqzYfioDkpg7ym3mfFp/pazTNAb
LYAcKU5AMg89hSvufofp0kJyVZqsqLF4ozi/9pHHoipCmei7AAkQTgMvfmQMCww4
GJIpwWEvryqRxU4pyxdtj+uKT1UjbenX+AdT9+coJzd6ftsT7tYUqL9scGgzsztH
B4HR4weGinf7okmWe/g6Ie4/6Yh3st2s/A692Fz+2MDH3/tEIwsX/tbRsapFSrMg
+6ZYFhuNFLbQRyOnihoRtPbXNXTZrlep9/w3NTKbzCu5HEzpYY4NFoXqTFj33jtB
y+ck+svX8v11Spr8u5V+y3gTgEaPhQPXWCIq0WmpAWimaL8XvME/RZPGbZHoyFQh
I2IrhZ22tJKsyl6kgMx0fsG11ImNlcHjK43+ASZdyhDCChWs40o8VAfjZOo8Pcyu
1i1M9Gu8ZFVYTS3vJjmUUcaRneX9g7PmAWxTbFqRydgd9kk4pf+nPXp9DWDZrYpU
i663vQb04N/p2Xo3MWwkOCKsN+2QhZw1fB7b2OjogHNu+dOeqSkiRobGpwwqhlLZ
2w8vDRqFWNVX6v94PtH26bhPgVZX/yscyHsfZBxX43T8QOYeuljdqtXtnmjNxJJx
8KzEg9hBvJyyDxKnxRXGW358UjDvtWM0XoBQio/eW7IA+Uhv1V5mlEgthTgdzBDy
2pVC52Ni1be8Lg0YQWEyonSUGuLVnLZTuI5Ukn826G3jWoFz2HOspzmiEN7EvqQX
/KjNaXv+10NY/3hcFcto+XZjhSR9lbtIEV+718YaBuLAZsk9f9SzZ0sm/B+mmngq
aFCplPua4F4zFQK1xB1TsJC8/cxwkywpKyTc+PcdtE70wOwGKhIGeztJRIPlqZSo
WRvoCmjULkQBoUuA671QYxaaEFxtKmGXQEMGu6Rki2xz72Xb1pGwySY0NEUQMiQX
nrNcwrx5HkRY9dSozAgMFN0v25QHSiP3ldJUGaCBPuE5BK6S1J+aKaoBLrsHGiDc
19ITtjLtnNammSffHjAROEG4iyFzdWqDosBJWckysxHJK5h+upBOUf4hb2fHPsES
uBgXitDovJUxzJia0jl4aqYyf7tCIeAjLN4gCPR3UaMcyQb3GmfM39m/D2eVa1xA
Hyl+m+szr4oAbPVvmCXlX3L7H3A53IuDA8CpUiNW9MY3a3TYSldXy4HSaViIm0Fn
tlTGjGlP4+aaLViBSiWZUtS9LajwxHxCowIIT9LHtMMxxYEIi8P3o8ovEc3QhXEk
yWH7Kf7wgPqrkJ0QLDTBvdAUqGrhtyUVndp5gE9cmn1OE3iC7R8jlpo9Gb4nB9X9
FC8vNqxzwR2nxvBvOvHDFJEAnyGVV3KxjQMCiaEUsvAwOxukDcAVBNF8ItlCOFJ/
wnRO3a4+Kie7wtMctPpOZALdCv8p0gvfqcckxtLsKbCoVmEFaj70AIgINayk2jhz
oTkwiPvMm+/vf53bwFuWobnsd7VGg20tUZpw5wLzYYcA3XrPQFPlGPLgAMm482uN
EGV8l/H7Sv0G6A8D64HU6WfRio7abcG6Ou9YHciomEH4nmKQN/tASKbYzXtbFkrL
6Msq7AHyo7JtChGZwI5A0nYr6ZisWkATzT4phP/Wp4bHmKTcF7WhIhTRD1LV9wjh
Bt2Tl9+G0AHXanGs87lCP5kF9laMf/Ej275pETSGw472um/8n5b9LmgDzPoEJ0aV
5T//w0pkqn6q38wZo4Lt+/noXXyzTkW5NA3EJZKLSE985+1vNR0QdfAurhgRyhYC
7bdNTdNqVMgeNQ4wRAuH4orqiTEM0oY/x7gQXg+sHyYrzfSKruexH0dMWvDuWKYF
B0pfDdIfN8iiX9Nj4/NK5uYXtOiZjo4FgFE6WctMT3QIaG9kHchmFHneQEGm6aBG
WhwpccC3H3wL7qochEh6m3THpgIvIAj/99hOhl60P0KBdrVdvp7+pjvN9gwTPu4p
K9JwZmbevxMIIXQ7pDCqsW/9LkIqmM5Cp1l2cDLiieEtXR+rIgZ+76RxjdjJTm/a
/DVfBG7ozuyIQU4sqMma9LfPHIFiBbboJgJKq7WtpVLH+cGd7WfY+67u4kFh6j4r
P6qh2w508F530J/oz25mmUHq0KTN1NldOWXAYbyGg7YPfzKt9+Ia9RF2BN1KzIJI
VDkqeZUcDtQSQl0BLfKMxOMxz3B8RPBDxSSH1mBKe4zHWRO+ui1aagMkCCED4S8D
ZWICXNXsIP+bgQiPan1/9lN5sk6z9mtz7PwwgPl4NzBIifJUX94r82dpijDxvNXW
JaeEIMuEWU6+va6qAaI4XglAfV2jFVySI1pTGF3yBtG40AlhWguzXB3AkLfsg/k0
d+I4KMGIX0yhJj9HYrpQuRBPwb2iMSiOazlI/qwz0uJZsKhWR4sIgSTrVECD8mwf
xNBDXdfjs3RqdJKAjp1Pr7kH/TpAPbQ2UGn46thHpGlhqvOk6jnXXxiNn1wLWT1X
dKdH1zp6SIkhEPKxUsw11PPdLD7AHCuGJ/oMoBFHeydRBD5dsmOgk1s/ebN6Tkv6
1NtLzPlEeZfR1mb32vFvsZwGTTVJUiMCxHfg4V/VJaI2xPZTJbGj4LxW1BdYBnYF
Hp5Vd7OVV0pulenWjahRhS+HQdb3sJHMOL/BT8pCWH+v0Al9Xbt27FwL6mYwbNpI
lD7J5HgXce2AIkBc1OEWcw5GKLpQU/yWsbWVcaAo3ipSa11gLOD9cWnTTbGnsRYN
05eBx2ZlGJu7wJvM5x6ElbBBAB98dk1bQ8tSOSpGg/zd9nxSz1ajDtLUuffryNOm
ae+f8Lp/EsZEJBbct+Q3NEjvDsKhAdyXF3cbj2npaUPDFzhSvlLILyLiTDSX3Iab
n9BjZJ9hZJnzagJVxHu09rzTuF/tzx1NBOLZbH4Xs8OkyyO6WUJWgBuHPzMlZtUY
I+BWpmE86kWie8ba6YkyukbbsoFz46V3vYf+prPKrcJbUa0iVjfm7KCmMkIAANgA
tmX4TaTUeVdeiXMru3f0KHVO8GbgSCE+7DgrGMhOuzKp+mXGt4wHLeXDJ79HBiBy
nCZxdYWu7164WcVxqGKA1dUGHfNqlwVYdW940IhjGKPmoTDJPHnnOtjltalGs7u0
Mr7AyLGDXoM+EbM6GCrkM0fq6NYnTF6GNWPDrfUrtKVF8mWSWjJEPdJDXbxkiedD
eGHq3eLnOn1Uv4r2NKfvrBZdcHRc9DUyLQPJJ80d5OlpMkGb1XGPn62IEuUjlEKr
sj9oh2rWUvQrPG24nLLuVbuwc9bBW7deqnDsiDTx7DFnuU5X5xTT1ZRkw8bbTux5
rFS3ZCIepApLEQLoD7yws3WoEnrhZx7+oggFJc89Xm5KOF9TVp8lxyLj5Z3n0ZtB
XqEzHduJyogRtO3442rA/g0KPCW+mkaYmGzV6g7SSGSBiK2jJDjcf4qIBlCR59mw
y/Vk0B2dkUruicAVDhsCEFCux1VhdFchdm4KjTwZMc3PiC2T/iBKwu+Mv5A62wYW
6AXsdKKBpqx3ltpTkvjloUWXltkLtvZozxS0iekhKRnbkPs8Tjh2JK3W70cchpNo
WzeOBs31pzG1Dyaojll/g/LFgb8dLXfSbuw6aB2epxxMg7/ulU9ukdJhi4hJx7/L
tyXPKJ8R37RaBNrlT5hQ2t3XcppCgZak9ZrTakdMXOIVXaxPTFsZWDBI4scO1lJg
Ffe1gmJLCpG9eskzmUWh83VziTIywlSAvgXEIUK/1SdUOPWp8k2lF5f8dgGAifn7
3lALjI4OSVgvffudoeCHtLD9Egjrw5evefMZCCL5tTzU5hOyXOI2tKmYrvfh+j1n
kKjkyindFVrIBDSNIQ+BWj8Ay0O/aZ4BG76I9CxSAhp1Z4rMaU8dsEkdIBFICp6d
M+R7emXc5yRwBBxMr8bPRp2qbw77jV/GlKmNTIi1GKDNG4BMBq/WmmUOcKmCaHYV
/57srl30OEB714tqLcugWcPr8xUbnlSxnlWQ8YF47HQm4xlGQ44rgoyURrvJA9ID
9xBhY+V8+nhGFh0Fr9v72AfUHU3hQqSz1Vzk2HPa56i0uRdueT/SURweQebPyxhD
D4BT/IHij1fIbatAcu7ctYM9+X9tBeODh1mJALyM8xjsDJOlHmWi9NOvlZzc/+8p
dXepVL44APgs3/gwdFx0zy5Isw5z9rsO64jg+UJPmBnNZvUjlzn2rgiFf2APg6hx
1NLEzHVhhk8Ju/u7KQ1nXncDu//fHJIjtGN4WNWm5WEMpv4A5cXG1wzv0KSNh3ou
fvawmRiTeHfivpLOzvBZLb2WztcFnwsEbmtWolbEqrggRtPMYmlqu0EtLW8T/4c5
qX65ApTi/fQoQy6SXc+JlzUP8dL6r9ILg+kk1kB435eONZ5ApT/wCQjTF+LieqHR
ypJS7o60WEyR0QiE3adFX8MSoAKXEIbekhvM3GbNWyVbeqYUNJPd0YHoDIWau3z5
+/F5QguddMYfIaVaU3LnTi9Hdf+WcwHI+ZwtB1ToWCmFwka9WFrYTADkoCMP1EGN
VA4B9FiZdNhLsDfHSkndO/Fk4Wy4506teoRvMSNbdg4HJS1yzF3DbPdqVrah/QZM
jSlQUq5OTz2LMMBgLq7vwKES4KFTc+YoHcncj9CXz3WxLJhdf839EmbAncZlZoTK
cUBZLVcVmxmdEKCb6BEX0Xv3MvZ4oLdUFFLmkBUWZ7XrPlVbLsd2zDQo4duDhL5T
Y2gxhtsTLvUyE5azRZBicSJbqIYQNWVP43l7XITLc/+VSB1KuaAZj1bM2zKZ54Rx
kKbxVMea8RNgQsEqVap5GiTSCAl2VYFi1jRV2LCC5lbCFjVEcsVVlEN8ieSDboTT
6m7lUBOsr+jo7dwQU78CYkPb91brN3EZlS8L52k+WoS/mCuhrVVT0b604xE5Ol4U
4xRpBfAGg8Wst1Qr8tlMP067YFJYhN55fZnvG3XcXPHwF9wJxcsSG0fgczLY2u4A
zygD7z4r4vy3t/JIDhsXPrwWXb3PQqdiK3R6DW+EZAiiC5o8d1UQR7BCQKNT7Xh2
TWLsXHUvC7JGBpmBO6ddE7zFgC78TGSi4rSN+jENm+M7U+Eq6Lqb++KY3/ZyXbI1
RbBhYtJ8prRGUEydfr42525615LvK6kBbQ3/C3Rts18bm1u1qNuPV6zuPkj3xxuw
LbFBF2RE9Kz6gXeFUv5sEj2KK2lTinQsTnXFjy6dVfOyWfNp8saKpIw8bZggeYev
8hX5BzW0RTV6zc2NNT2QNRn8ofLXHmclxYb8km86Jm0Db1AVe80Kl/JeXU4yawEx
koT2T3rS1sEyTHWZNYvFyWLcE537vZ8CDayB6LMd+pWACpnUrS0BQgK4N2H7JOMH
F+LoFlFb5gPbDY30QA/VjdJz6eXdso7y2QGjkTtKG2ZJpjym4/39uAxXqoBlsh6R
NvMPgNQD6lYkprQFZTO8HaefooMFCSilOMEClN4tzIJpL6PQW9zji0PVmAWChASB
SsnAX0aiytseZM0s59mq0bIUNxoK3cPz6OJpvgGuCZ/kGfK1GwEOv+qdlI4W4eqL
X3XPMYK/Bqr8+xXIqiPhcCnkbllkYH2eHkIyT+1j6Hlt1pI01wfZbr7iwg6vgSdV
xOVfbE5JJ6xyiMc2cWjn71ml8kNMJYR81KwOzVwINN4yDBgqFi2RVyEU2b7JP3Kx
AQ4wwnjh82Cv8097VnEdalYnL9MXBBNQntRZWBmM1D0IaqyHgNZBbdMbPj+9aFvf
XDIpU7405bag5WSElrPraBXkxP5Gb83t0QzhOItLC+OK6I8XYTMEF7fqLf2EF8FS
Xq91rx9JopKhZKGyLryb/2c5tG8J7SYtxJNZzJ3U9RBCNCZNrg42qhzY7cVAzow/
pH6MqWtlZuqex+Pzitpw7MQAXUozd2/t5aCA9FYcLhPTbMYwT7LsXVrAM9g5GKOY
OoGB3cNkSNOeYBDZoKRcfTy+cUjIbC/y6VSBvLy3rB/lPelvxENAaIluHfmKp2/m
qxNwyON9pL7udwEKNiRNcYuOW0b6zo52/La+q/V9V6I78+W4VFndvBkmBy+pHigd
+Yrc3EzhRXr+HVJuzausbK5hX/IQqMaECSQKTmqtEaFh1H/pFkXAzdRNXV6wswn2
FT85bfyT+KpgOW9zowODf3aG5kFc+GZbA80Tnyf4LI4b6bd1HSDQUIzO4T7RVrZj
GOw4TQvVDjuNydU2dYcDrOv6JoTP8xAdOx+Fpx+YoJpyb++Fulbv5Y2B3EZnZ2F8
dKuYyc/GRWsRyxz/IBz5EqNViYwRzCnyMQNliRLhQGhpF4zvpA6kyIyyBTHQOAu0
qL13jPoP785weWS8MXibjUiQM/5nsxWW71CK6Wu0koXPqnL/wopBZ95zywZ0Jgaa
dCb0dIROcj/Wzt1uUQHtPr3Ce1/gkXuKVCvG6wPVUvG9bXOxl68NcRkvyfOTiZA8
CDtNbHId/qIKe2on5Q9IjcxPrgtEM9Lth4HzeB2lHSvL4xls/iZb+e0XwR0ln81r
YivjjlZ8eFEkFbieM3bUCDS2hzWOxO//LxfUQj14l14Vb2c3/M7jXKELV7uWVCe+
kWgI7swBv1UUVVRROGryWbULkJz9/2e+WG8kEV1MpFXfjqXLfGB0rvLwraEUL4AX
yMWxCHae0Vefds8NejSsMiX7cmcEyANpPdDYOXFkbl4joEQvruynQBNe7zPHkb/L
JKhYctXPGiRCnyGlTkOdw0WQzUrsa/InOgzsS+788sCMsboSFT5uoivQu73EOck2
e/11xDrXqm45pmezYV0TonjTeMUGhhTSvrmO1CO3LmnevoN/bSj4UxBnRObJSE7W
H5Tt+lbYiZsu+5py28Cfsd8QoqoPTENFrX7K/2rzTuTEXHru8Y5g1nbVAb9F/Bhz
LTMDIdyaOaJly6amBxmLMg8mWi7/4mj6R2pL3helWFD7nMTgZuF4TfK8lZMjiHk9
j48iTazyUMshk9z48rcM8eROFlfZfROUnr8MJNuHjSdid03dQvEmz0ynKawmsrdr
rrHRP3NPGCK6xuqmC5/9zPrRxms+eZ7lXmdu7qETcuXo37VF1QsCi5vqErdLWyUE
Qs/WQ8gg6NWRqg1VlGvaLgROHRCt6dGJy5M+JZyUYnqEF+BTD1Ua5iH91PdH2HKb
70e9zaHRXq5k+bVeZs9mYXbHdNY2BASFd7CymI7HEDD3xGMrPZSvqkAaTGJteC2F
Kmwxrva9MiYenabNnIlTcGoj/KVJsyAtmVxq/bqzkYxjUFJvuOeyOZXKd+0E5Csz
wKftKlVTvXD9adFmTjaz9QYg3mL1KBzqJketOefDDeDETQa3z0pjTfMOUUexTDF3
i3QA0lg1J1wF570qfAnz4y2FjVoZUw2GyYHlzS8/o+TXgdwXQseHwxkWAPMX70l3
gW/tr9I+wJLOpP9IETCi5iNBQZ3kIpi3vYhjvu6Aa8xOPmh8d2QPdRNg3po2eE0c
/+NWT93r2uVZUHAKHMNwRyiSkWJWrAp//z75hCli3iU/qOvdDVy400mLzySyYO28
laObZAZH0zGzMB4Fhb0J/97QPn1hi0kS83g9IUX2zGi6f94FSdOC+1uBP9YVwD2O
0VxZQ/AS2Ck59MMiiQbaJPtMnzZcIjh2S+qpps3BzRaZrtNsAaoye8fFYn3cGXML
vG34WIIlEqinbMDzn0V+/6D7lsC/thXM4PhHPU40kVGYa6mxmNTizQB6Ue5L8TY+
bJrNuOralVkQstbXgyVQHPKojGobqxOaB7j4J7B7cbpm9YaeHJ3bOxjZuhAVoEku
T2lxb4oyXzSch4AWKM9gw1bAOAuM3fjdw0JPvzuzQ9rzbQ1BjwK9bEUQ1pfP/I9d
YoIJ7vzjfJK9w0HdVEy2ORwylyvr5VIQP0kAIDZC2yRZRgy7PlD0gULfe8/Dy26B
eJg7efRiNc+kp6R+Wm5v8Pi+MMhROmk0/TM4At70M+2ZP12an+n01s5TfbyK3Pjb
8SrRibQVURnTD3AM5DmbFU3YC0H5HXHy7o7mFFsRmCIEzQy43oSSkkqLJ3gxgrT3
Vk6ZeH46jYoUGtB4oORXRr/Ay7qfVEV9M92daBhb5cJ+WrdE5ZfCFG4rHiiWpDDC
nSLEU8UfCRGM3UD0Cuva6V/rhgq/0zTF0M2hFt/wc0lf7k3GKXb6x8V7MtPGQ4oo
ccRu3TzYq2XdckqAPgfyJ0BongnlpmkUaDqFIXS1PdlwtYnkZzzoKpepONs4fARL
I5+akcjEjS9qmSiXcSe2lgHkwYda92+SKOR4uEeMyNWjBzbDkQidqX5Oypiq74OZ
6WggfzNW851H8gjnGGUqNE/YIoU3AYo84twsBI8tEH6xf2mmLNYdT4epJrkj2L1g
YzkORHEQ29QaLnlEOBh4MV4CrrPAa2wmdhJpFeS+vKnG5IMoKllJyrlY73E1EL6A
pO07U8rJwYWn7BzBobva7sVVufFSFDiuvSXZ698GxxxuRR0whqgknLvg6O/+Yxd6
XylkCKhqEt5ZrWgfEqxzQRTMS2AwZnvgi4Arf5vCFs2bxY9z/6WL7DVqP+/FAH77
iGFRpV5jeOk5Ncc3OzEUkTFi14vPb4r6rh1Bc4sO6mNvGTrrBlcbKbgQryaU8upH
5XYlsgmDkLjt9PvnaYnMzDOF366jsQ2mP3nS9FoNLRIsxf4knQWOkZwzaZuLFvpx
4qwf94dEa9VElb29EhYAjnPMXnu0J+IvWAHqF1Smqr1/WJy5y8dNae1GEqqH2/gg
ZJqQCgPJdQtBVXjS5vqtfzNHLPcNAH0nu58tK18pOw0VALbxbmdNUcRI4KOEwR4K
YIZ+QFW8j7AFBeZTcZPutUEec8Nv60zan6Xva3xDK56z02eMMN0SNO1btdamyJ7j
Mm27QBK/YIfgG77PZUu2ssTXLOcFsmyluxdDzHxN4Do5xffHEW7eubqBazSlZPoG
V3rDhl4BK10PtCcEXylw87Qq63udBrn4HCI8bUJNxryA4nHU7lZg69k0zPnQokt1
JttM0/TJ16IJw1NfzjB4gEyNkXuRmjPItiJY1Ybgxv2WpWqXbyBvOdiGdAr/Kdw9
Pg5OJ1zdh1+OLqYHV/kZ8tkTXWXI63Q2Ks2ZcJC227SWT6cJVWh3PhssyljZyNMP
37FBuAlEyrek3TNhtABcwenrdK9weTQWzsknF0W2p2J115UB74tKDR2oAyzXJ0SN
boYToeWKIkYN7OG6UFIAv1wobsEhHK4lLkHL/VTg6c4gBVwNo0GOnd6NNGTsgv2T
ihxiGtWkfm3ImSUw94A7TVubI0KMv12rcCxszv52eUo6ZM2v39h1i6S2hmUD3EXI
j/XawbEbHvSBDKJg7w5Bd0iA2wXpCXSKwMmXe6N0Xt0TLHuKbQOYefKzSnS5fuiv
GB2jdzC+Eej+iroxiDFMCu8H92BS8oKuzCUNj9gO0XOhWF/7B+ecajy6HGjvoTUq
Qibv04Uz7409MFs39E+hUCfu0AXlCDmdIqpFMv1YvdWCLyLzh3+tMLgqx8Pk0Mha
GvAa+JgbgzZk/abXgBRiAgR5bCVO8DI6AoWEyqPQMJudFhLvs3+np53qkeGJxKPA
BxDX3+hFT4Vm1n7vWRl7b/VydBerwz3Z9mnMdjiffuKM9ZX2nrmq2ZmUQAs9GdMo
C69ZV6GHOAOmCk2pCaJeQTquPALtjEadgvOOttUcwCEHjcHiQQlUd2x4pKosuzeq
/lf7bx6tbvbAn8wLfo/rqTYdUkEolgZ8ucOJiXcZWNvB9PAFR6rRxKuIQ/41DsVw
hOrByZaq4fIs2dbyqCx5a0BgBCFeW6HdgzS++63iv1U4KZRtNUulUqroYoxtzGdw
tTiDYanWClAD8YSPZw3/Oj1rKJszYoum9btvenpp21cD4S/r+vQT/ZWDk8Ac84Jb
gX1lJ/6pZdi5ReGbRoiY+9FrSKNuCAMMv/uNWfbTKS8WwKTYx9pFdfIbgmDGO826
rvUD1rjColLxOhn0je5pplRQiYURRHo7wd1C1wwVnvsSKUe7oQEI3b3YoRtZCU8A
IUXpMrs78F7g5pxXnr1YSuZax5lF6iT/uw5kb8AjUqg88KQANhdIqSXLNLgRA0ls
P2liZ8zpGZ/kKEM1p7gSYiH88WZhb7yIwJQKH/NCrgaHoG4cs5RHZ19U9HlK1cp0
W0tDINLI5DWldYQ7EYtXnyz8zxJTWRtPlI1LHMO03bVQEEEWNeFUpUUpMJHLcooq
ypHuXoA8ZpQkzpPU3ON7RQ8CwTPezYJNiVY7YIOycKhFsu1NbFY22036tRYIybfH
l6dtj0UA3iiIIJKpcrLbDzhmWehhjLmRW+cAgoR5FoWZaHH8GOiulkCTYlq1NmcK
83j8fZGAe/LlgHH5WfXYSuPN4w0DtYOzCq/J+m8+bWL4Riq4Jq4MZAfcTtz2iZ97
Zocm78x5Vot+0unfGbq25WoRgBv1wcpubrUXTH/G1TYzUjRSp4clVsv4dJ8jcZvq
C5i//vNl0JJLZRizXiztfMO4xk9mxwysY6qXbSqPikg3c8xX6G9xBfqTQQ6TjEnw
3MS93EhBWKEcXbq4c0nVAg9X2xnBakXwbmCayZNeyKzNxcgWaoql5OwiyYN9isPc
tskisk14P9qezuquKPopRkTb/HBZA2Ek7nZaYbP1Imk8K0GyO2KIy0gmU1FUmHUE
wE2Pc6ts5k8Su6FU4733zWb/cSiD1oN4FVbjgeyP21gkH/9axHHKuob1qXax7lIN
Mi6+aNY01L07Qu009AZPb7oz50m0wgxXqlUS4pkBv9FkgKmUTp2sSWWZIACJ32Ek
BAJJh/Ygg5FllMwZRhaU4mM17GSTaT1A9TNV4bK3DkSg0IZr1phNUv0xNmn6Y4j0
GPK7/BfE3z+7q2GfiWknPAGb6VQD8/j4VslxKvgWC1DlqWci7BqTPjovEfu37HTH
87jqEoDArmLD9CYIl8CSYA2zi7hNdREzRis7ZfES+R0g8F02z8Z9aloAY2aij3k8
FwNm/ttja48RU+9NYyQ2fb3iOaaFJfl8W5eaE65vmIPLpb3HRxWdfs3IahxhGWNP
EaE1v3yLqse7MAZ3UNc8PNwxQZ+cGWO95i6uT40i7AZiRWk76Lhi3NRA0y5xUoj2
jQdp+md3cDimLwQIW5QOcri3txW3W09uX/4LNSPFUaRfKYi1kZcx8nr/bXGvFMj0
/0zE6ZknaN1ZNUZX74U0KL0PTFvYrAzK+Y65wfZV/bfOYGJD+ow+fLzrtJfeE0md
zbzE0ZmBkrCpDDZkDeEjO8vGnQ8T9JR6Thhm9UzNGw3m1ex1eILZikaqucgylIL2
HlROEYBr0npqymm/o4qz1Y/ox6zKpegeT4vHV55Kw6Acm0jQT9UsNSFj0ldYHa3I
hmlHz2K6qS+3nXnahUvBoybY16uH0k1mKX64quKQ/MEG8vPK+nqoJGtTMQCAj4re
kq9e8KJl2HZX5ydecT9/XiJ38NgLI7sEFlSzjgMTu620iDDsSKP1MQ+CG9JKgKSO
q4GUrlrLVUh0OlpROHK19B1pIlI5E5pd1bjWkm/wLXrMz0skD4Shc0tIxOOnFcKp
ao2wnz3luOZ2IRi47NIrjt7tUAhbQI8mprKsprYV4gB7Db86raqwUjmJzMxbkYXl
Au2ZBVLXA949cLafIlWZ+equ9tYyS2HMJyz5VB2eo844A0CaweL0Y0ovDUoQad0K
teJitvnjp/eVrPmUs6aGjr9i7R1A8a6/gisDwJCmBfZB5Q+irnkaqcm9GmtixIki
Eq0KhgRvXFzmMK/SGakE3L6MsiH/AAoq9MH8H1BlVq6odsgf2Xn2E6b96tasLh9r
pqe2cyr6b8RV34P5cgQwUyl5rzNosDuxzHNfdFA7u5UAn4yh0g3ySQ2bYlr8B6rj
JuiFDbMd5+w9KNfF56xbnXx0NmqA0wwsrUR57McKhe2q8AnOTKHg8UqvrhZOezwt
VldwFqiqHqJhfBTWPwdWSgLCCdsUlr4zSkTx5bUVpaFg7CQaJZKuYYrfB3xuj5VN
JEwASi/nUD1cj6KGhl8PzvjFHiGe5FaWz/Ze1UjtlG6Ooaw71DCOiIidpVTZeXNY
q4Ghcy7S8RuK+XzPvOsWgwab+HKy2pF8QZ2k5WO/jIj6/gpuPBhWDAjTSc3H0kNP
yOJDLM81ZGyf9UkiI5PXkq1Vv/0ySzcS04P8lWzGGnPOBZMaOOuw929Efg3D8GxA
Tr0pLu3tJuGvG/ZLqLkRwGRxFu6W9HjzpLrMWLpdQ8hGA19vHARyhZiv6uh/issL
Vz3BPFhWVIdh08I6sYsBnarBeb5tnp/ZUdzLyWvj1EUx3BQR01rtHIZcScPRp8//
c1KFudOKeA4qhlImU5z9Y34A02cf+kJAz2/rAgw33vbKBKNLhAJjRvLITIleyYYg
fLk0zMXs3Bmpj6CeS0H8wKP0PijaXJKptUDzxLMrZC/5BEjJIPYFXOUfEUlMq3K8
7wohTsGEVoiAj06sB9SFqfPuDLXhp3Y8XUbwOjSjufWjZIxwQEmc70UMuzk1uucL
hirO4NBXtCoPdQtMKdfTWA6ytsJMR0Tisu20+fY78zpVEs7pUQxMArjwTr/Eix5S
w5CY8YGhCbAUennX1UJKZkHXNdMcEdmrLLKs+84eNP9HM+uePe3jjGLgyI6QGPPz
QfqR/Q31MY1E3gHxHoos9ayzuis8gTL0mW42WT4A0u32uxbibdj5TGAi8Iv/GP96
hytupiCporAibbXDWFGmXXWfzBntXvWpFl4uOHwbJ7kilpyZNw84HcAkEePaa4BV
V73oxZaKepLk/g7rcJqgYMMn7vtoCQ9DUOiT3fwOVweXayNm50UQWbCQJIQo1lHj
7TY4ilxfw+DLlBxKTX6DSMNQgaE4EVuK7SXFwXNS6SFjzNQozqogDY/jtCae73k9
LKLtNTnwjN5NiqSEYeatD+wgpiJljT7MDjjSPSPDV+r285Y1YblMlG5z8NQRm6L8
a3uJ0xrvvTvXEZxLRiG7hrwyosT3peyp1ZQTbpGzJgrnR6anYzXF5XrcUodchSqY
3bWqhP58KmUmHB0itIdrMRwkQemB/uyR/svr5lEQKtBXuL4lwCDO20nk/QKEwGRg
uMdcI/+7giKuR39mKl34yojIVWeElyDgGhJU+v60fdnrsOP5+oL88fBQrKb7wMhO
M2ODzNoEi2QLxSUzGor+/zEUQOU59cSZRLJH0C11jH86MN/cEYNhjFh7y29aPIxq
vf4XSGMvi6avA0FXeXbEvHdiq3b4qOY46M4Xy3jIaUns1VqIK/dPfPnu3gf325BB
0JFvbWxN5wbi0itzweLlvSDklSQ40od2x5b4BwltLTKaNsJaT/0YEV8hoZYInSDW
AxBuZA6wEp9YsaeQVSo4sPbyLo01FNrULTquIqQB+iaoD8l2kyiIRtIwCCrNNIhd
Wqe/kvQ3fMVA8RtCKr46LNRIndm+vL8TQoDcTjJw/XBoOrrOZT1PucuQpkzRArc6
fHqKGPgij/0OHwH1LlqUtxdUF1aIbHwOIALW9QgBphUV/9TTK+sNmVI5lEoJVbfS
z4p6WJM+sVQmW2vXkx9nQHWoTnCE4z6xMws6TbATPPGkHkNXF6Y3s8ylR7GWYQUW
EXoQagR+iydzFDXu7Gv6D9ZQIeIcJ9aBnUFVXvyip0R4/yLAZ4pPevtDUFkhykMK
LDah/OmNRotf9YE//iHzibL2U3+SnUcwNSRqrrgLuBtpRDLHayQKss06Bh4tQhRW
Qjzv6gra/w8dqmaejUWugBRXduSoEZpUuPh5CkNoS/RTf1VWBn9OjcwMmdmdZ54y
fRdfpf11WRF19otGyl7UAqLWbqYdXVPVkdAGp74+z7ayh37S6WDzEW5z3g2I203N
+IPECbWOoBZwVavgNtqdCY3SHo/ynFQx5xfy34DOzss67VL8kvf0yo1GscxvUeR/
cAYeVqYYNx/lkN6JJ999Z4Qu8/lRLX2iY+w7aycVaLbeY8mRxT/t+SklYJezewUM
MQabbTWBQC+MIR4qEqa0sl/oSchsoClrK18ARDF3nSCv79K32PsF+QzJccJYSBaj
ahEwRkCEFU3qIS0hw6A85L6AyjFdlZR952/dkPcunbufhkWywcYLDdrct65FU3mw
eG9rSPT4jIqsCejj7uGjK00uo0f6om+aqe5+iYOCkgn0kERW8rmd05RhNaB6Cjuo
E0mEouISFIl+pa8DoRA286hUR+aYOcuse1HlaqsoZCbcsPDqVG5HROrv8xy2DRBk
kK9QSCdIdwJzRbyd9JKRhYAE8TXLvgvTxv4nmDsdyWt/5ni9RHtGq6HiNRhCjKSO
4hQzdm/ASctL97+yBbTm+xJDk4MXWb6r0YnrAOHg7m1Oe4mQkiLF4Ylldc4l+lbt
hHLKlBBBbiII0srgulYVaSCgGKo1NCIShZtu5eheh7eyKkhw5ma0lAV2gzW+c4jX
BJKM6Q6CncrEaNtNMwFHq3Kzr/5rYa+GaJB91hVt/okQ7WwxipTKTjAJ/uGXJYrY
YBJtBxxbIycVe94EBCwf3xBAmA//HSsPa2AqJVvEVfAnKMJK08sbNhU69JuePpGo
8WGpst9svmZk54WpT6Lq7H0M903N18kv63JoFA6lZjrdlOFfdkGAv+oRiamqqc5i
FWWIeOPrTAMF/oNIMIYpXPIcChDUHQjpCn9JXWc4W2zv09Af17EeZYvWkpmEaawS
NgBkbI+nmsqMHmLbB6X+QWikYnfsatID4r8o1PJ0o1Trscp0uDk3EsgNL32YTfwf
DeMUHLVkErx9iMNm/8r7xQFDLH/vHYbTeqTgZhM1S/fMusxwjMnCh8nkxmNDBfTi
FX7wrgR0Smx0o+0ZvMHsStBDz4wZrqwJvZwcba4VxK0VyNCwF7cm+9nBtFxbo/vB
axTqjYDHCANlO1cYhYOtidzBrOudN15e+gdpOv79ydXUYeQHpSr2SHcFtt0eamDo
2iVa8tT95c2x9Z7ZecYuJ5oZKaZ1zULY0aVg6KwC/K59orzCN3FkZQRvLFfDUbEK
Zz8l54xSfAa/Kbw4rDJiOPCgMng+DepbLXQBRXC/GSxlsMvbAj6LWPS/cJrXk3a3
3wsQj9TbTb3mSqw6FhdIUH5KPIbVDvhxTnWRhfuf2/BLUTASXFAH7mIRhQLsVoi/
gOAI/qfXRqAxIp1ry6Gexi3QC/ND3a7cJEY6XFSxPeStqk+uiE4iQAHNDDQaKDHH
uM176gp3p7eAt72EpxSApUTkq4x9lmw2OM46nd/Et3V0rwacdxq0ROfj7t+gMH2j
JFF8B7yofjOLkp7DXkeCeqfrO1M84xFdlEKKi//dRupm0XXU0pxtO6OHNWm/d0d1
nKxFfH1bIS5vtQmNllOmGBwqcuqwdK/HM3rZkBrjEBgIte2jEeTdvipok3XFnCUL
vTUsB7kH9hVvMNSj75JbVt4zeFe4KTJsLhYxxlqoeARpPlc2uyJbNxa05HErKwV/
AvdXoQ95Rp91k5sFnoc7bK425MgPvDx7UIk9G0lTNOjhhpnWQmmzmV0dzu78YUkD
bCM8ZnO2wD7c3J3uZmciMvd2vIBKduhYk+lJvYJ+kND0U6Lrmd768xBlm9jm5nqb
eQdp0hLM5WFCOY40csGThZ009cxE6IBu2YPTC8cz245Tu1ITXGsx1ymbmrMeScUL
Wup2hn/kzOnVRGF2EIQnAK+dPWzDQzc3HDKmMGD86Bq+Op1NiD3VT/BjnsM1aV1l
BPLQ4+JR8Nn8pobEYnzWWVxeFr5Q4A0tminXGkbF4hfsLIsrKb07y69arQaDQ4+e
fHT7/XqTdqVKGJYOjkbhVwz1S+7kjKaoPHd9Etq5tvriX4mtOat/g0tqQC6mOx58
8ZXj8cRq3N9mSwJGimomC9dwzCTFgiKtrYUT562MCqDDQrkxjBU/uOAjzYr5VPNT
kXTwhUtqZZ4vCPjgfYt0F+Oc1AzEP+5gSSyoQMMyj9Qs85nVELlY0SCPAwIGf4gc
TVkaZwWiDahdkX04Zis8CrfIOVaGv4TWt0gzOZ+3nX+Ujh0u/dvENCZJ0kO979p/
gErx6emwkJWAjekO1fbttjnv9Fjr26DnJTtrkOOZoN94uW8LFt/MSc7ve2pS2Qlv
VDYHriXr2RbGz+70KmjpSZS+DT2HDOn+18K5xEd8TEh9B7l1oHkdZXbp92dgLCPA
H5ZYCcfp+BlYPDrYZF0Nkf2ucTqdL86BeN8MZ4UUNZPPj5obMOG+JVuWCEBXVDLn
eOVGx+EBDffOwhALzeQVPbi5TzEAnQXtYY/XD3Jo3pgkZ5Jua4DSd4nLiymp19EG
FUaQvmcRpujqKP1eJOG5BTrQz2iPiJx63u92FnC30FIzmYN7H61OL/xnToyZb7F+
VWSYTVxL2/wqMl3wwyYGX2LdNmRj3JobupHmLXyPl+cmuuSkIlUc0MfveDDGg/d+
AzmUWw1nfmZNNI2cDnf5qoib6T4CaQubeModTB74s5fvJKrCQaJm1Z5EABpDRT2U
0/4x8W5kE7rXgOKluAKRToA2ZawVOraXtxNq9lvfaWl3XAhEMZkhZtYQSaYeqxSI
dJamkwWsRxMWNOiXHHMLaDrV6dfbEJPVMa3zgN7/Ih/n8UbWJTaH0AWALnHQb9eh
6o9Dgh8J4KPeWEoHeodw1YfnkEuRwvFo8gYDiSHOfbhU3mdzEOoEwor5v1vDc7y/
2abFQ0a9qSw1geTbR34TwSLDFi3wwqeYaTNhCXn0IpS0nMowgoMIkWtGqPqqoN+O
Y9zwjNzXeeeGtxE//Tl4E71fJcde/FyqnAgtC8ORyaDtNRC53koZJ0tAR1Nczzd0
X3zP6P54cQN40EtLJsZ9qKrDr1sQR+DnLmX0zfBVUhZ88LajVREuHzbmdu+IB3Wc
qdt9nvb3NvlROpvI9RTnVZbq8PDqbGnZpTHAdEVM6xQ5/PqA6UmBqFO/3m+rBBWV
4BYY+bM57asJ3/JnnHHY51qtAXgWxRY3nCNIwlR9sXt0vLoKnza8nkpoha1v9OjO
xU0nNZMDq8NLgRN36qq4nn61tNh/880AeUfKiX5upUC2eD5PGmp5vLr7sr8sKQ+U
6oM6qaM0jtAf0zctUFy67t1XYf5kIPq4o3l+O/31R5+0w34Am/6qCB3qp/hP7P9D
YIJ/yW/3yHwDBvSTyg6LS8hoFhxpClILWMNEdm/feCan3J3oNqDgeN51vvYJwUzC
ZylilSN4/RtIRuc/Y986g1CLugQkh9T669Cl+1BCtKgVlpC3/2ynWIuyEsfqDhrU
7geXRq5YmnrxFUMf9TDOpOmZPf/Z8hw2Gh7BLwR6V1uCHDkAz8badhTMmizYIrYn
bYLXZvdD6eBlhDT0jkvfjc8c2m39XaKzi6LviZHvCVcmBEMT9hVlDV2ZDbRNec/k
L4K0VvTVQs982dHPtzIt4mi1BS18QdDIYaYur13Am7WzU7R7so+Ph/0dsmFfL01b
1BWQe3pjtLg3WrAbV6ab2Qbxnx65dKRyhZwc+SWii3eB2qgDJqrWamPPuxJ8IpfS
9KbQQO4KANwmKurjS133GTmTlQczFMZ7Vm426BBGFZyrrKfbkOVzeJRCeaiI7zoE
pfc6OVFYoH77Qpfu80w/tJE7zIXmp8sHEu/i5EsxUePbRue3SgatrMKhQe9VjgPu
oIlxSdILRYxgweSaU6JQOo/S60msnISQ7+XeXH7dgWx7bmIS/UdmSspPjG2QN+4J
Zwbdp6/1Hy77UyMYXgFJxwBe7CDF/w3qZOKPZmjFAJFb6JdAtWBE2mO310nbApDR
UJ5fddU8a53npYXLlzEjb/YaC8wUejb3okP1Ye6gN00fuUBsq1L3OGpAOQ+7Fokd
3uTlFV1l9fUFRebc3kJcjw/Qe2MK0wTpvQhwpaxdhHK4/4mexfSAs+7xSzC5xASJ
moLXfEV4kg5bI83HV0gQrXS16wsHvQ7Imv6i75PlYHZMfr7I8dajc7hVnN9mCmDB
bHRf585hDgENufdUDWF3UrhjzqMwd5sHQ17iAddHYI4XJdhXlOyrVHEC3b8cF1aM
UX/fH1VqZef1xPBtL6O7036oUvuxI199IkSE6YHhWud2GH//YppKR7mzYFFLgbxW
X/urWmfnulHNBCL9O6z8aztmOFHRWASP//Dl7pcIUy5TStTgGKCvpImLx1szX7jT
ZdTH6dV3S8c/UkxPYHY//8b32lp5DPgbnVugMooDxXG88gCpkwb5709nPIEffmIP
HkubY6z9CRS4PsZdytiZ5iWqPe5CVGhuVfKPt/IQSCHjlI70Bnp7aagGkrX2uJAl
O2VbO6Hn0PZhFR7EmQUQK5gfpxW2sZ9exHBK+gqA8x/NaCZxqVQTozdu2wcBLxQG
MeoxnZQlzwMwJ5aRbvEqu8CJdE3IbVITUsBnpi8Og6MjZ+Bu/Bith61dtpK8e4oN
XXU1bcU9ZY4xLpEqBwVzzlKgem3mPrUP/+jkxGvpCgQA4z+r7W8b+IlWre7khcd3
pwqjzZ5e5pLuGprM4T/HVLXbdWcSSkruDtqfBGyjII2QuYqTR1lonGtnNyu9+atB
P15az/TtX05Yl86b5WryJjm3EsS5HAegOdlYR3zWmj2IdwsSdeTqEk5MOuwMVF0t
EB117Jf0AAQ2B8ogKgH2p9ZhxK/zGdIvoxP/27Y8ewDT7WS4QFWHtRn9lc+sjukB
6BEK28S5lXI0M2RdYfIPdKDotEEsAlc6/adK8W2k2LjjwHFs3EppTMQCmJ5WA7D/
NY/L8+JWbcPDeFEWkUhSRUaO26kPodebJGoltCdJiKGS40/O+oQ7ETEaafMxADWr
DbC+UicukPCnAOVIZLdynzkk81Rk0T5LXpDBCgJbDRBg/gl1N3qDi8U4U1tsO+KF
6jvQ2Y2T5P6XTNO8mXERh7Idv25Y8GgEzN87kcllZmVnaIu+FebSctVXwXNPuHzq
SUCEYpnY8OHFuCyeNufeF28KrJ28kRcrOD8Nh1fb7b183OcSn8cTIqC2WcA93bB6
fv55iZcx6tCzQB16H9PqKM5/wiSdTAk0QXwpNarme/SXnffvvs6uoGJw5pfh91s/
cOOFjrgmM9ru8N81usNkbiEkNtpZhYp10RTzJ6P1e6LnucrgD+StaWW8WjzWgqcr
jOQwrYksYU8ZLYMBEul9UvV9FGodaaUX4uQ0Y/FoVBVzytJ4WAClkEBM4ESb3mXO
bRU+Vrrbxb578eu4l7tyFWPoQP6airg8ontbWENVCPV+Jw6OeeJWUBZ8xW/Xx7S/
QYWS5pjz1Sfq9/XJCLxYQsa9cyOdGRsAs3DjPEaftKx6u3gPKLoHBZNNtma8+s1O
CKbk/Iq7iMziDJCWqLGqWysxeCqwmSdWQlhQ5J//8q4r+aYQVq+8wR98oUdEQVwZ
WfbS2edZHg4qSTSyh3HUoCaJD02ZEfL9Zmu1gtHqdt7h4FB4nx+MB4AWCHZZ8sg7
RgQF0IlbjtO6YdyHpZZBvcJ9+WTL61jfy8DBFtMWXuEf54gVtDv9yNmBbDO11dCc
FRstZvvQiYP8knHr2CuudJ9GIrgNmuUnK2gHOdigstgv3Sa0zMXMqub27ST3h8zy
P3jQWlsBwytnRu5JOoKKOmdTWvKIJnZ6SKjon46HU1DwWipryH8Ojwfkpv8czH2S
0s6FUp+1wZE+9BxvVNgDR9nNV91k4J1+IUc1fxaqn5uitDpIgDvPfQcgvkeZF7Ad
fU+C5OgXrrTTzRMEr3RUAhRLwsV4dOKqDs8URREetZiIrf2CirnaPI2XvMd/KPc9
02LnXRSHAf7k6kDLzXdTeuiq3uK7Ryc7p1z1Tehn/l4PYkdoHs+JPXgFO5KInyr+
f7TDov6SwHAz8K4YjFcJNM+3+qgDZ/zNZyG1RtRzvz/1YTjuCCIbphFhp0GcjDaH
GlCm+dZNRqo7OjOfTB9mavBR0C0MrMlzrxa6Zr/LlUtoiBku1ZFovEYxgBNV587Y
Kn7Kn1YLQLICajiBogl1Fw+h4A8QyG2CYjLNrU7cCJhwZC7DdQeCTULQ+nBGpXxo
B1pAjanuHv/Jqs+t9zOdtg3g7RJchrK1qtgnSgIG+rIoxjrhEPHX49mHMI3/LDls
f/I5/2YQE4APz4368qtUwlzCXIMUNPas+6Tv5FxW8BfM5kfHGXjWoPtEoh7qGvNq
LdM5cXj/MV4/OQpV9XeoJV3k6ozyT2AhmtR1WBmCya9MgHjnd3FEf1e2cOozSOjI
kjMLW+P4WtDKTlwfzAj1qZgAUfnZyFsyF/D6juREJlu5dLFyrn0IhL0H5FX1en8q
aKs4NlGvZrDJer3AbbMXAEFFJIF3FKpt/Hp+8rnMHmSUW2MQBcKY0ZHadQ2AM0xN
DcdowpnNZUAb5uy2GHaB6wuCtpK9LZwhVIoFPW/aYmDqAX0F3kvC3jH9yazS6FoF
K9G9S9BWbgwHcGjm4Rf8TTLkhE+zKLz7jq2MtPpie/VX9JHv8iTVUQMI1iQY7vOM
nZDf2LAs2ml0s3j6fTLLD/SjA/EzYXRRfqkZl6fpZysIUcHnaomamRxlvnmn+kMo
7vDlKRFIWYTbRw1d+NAyDdHHT1NWbwgSPKQDMYAmeEvUNOtN40bjBNZ+AVfRdz2S
Qbs/8Gt0ZoYAznkljYmITkDlhPdTkQYwTs0obFs5fwpG6S8z8xPzdk0/ndRxcH9D
H37jRNvr6tWePoFn2sA1M3fIyvuUMbrmQvjNg/PY9m0eRe4DN8Sv7/TC8gPuHU5w
yMf4yrkGhl2ZNWFC06Ja2F3n98unne8SM/cDoNPel74C+05Oa3dswEFTDLFUXc10
IlG0A/wRZz4Tp3h72Q/+UczduY7rHnoO5VWyM2gGy9bTtk/rhSG4yh6VfIdXW/6O
vRJwFB1ku3CDtqHLQoIvZp/1uyjfQaHj9nWd5F7kI3TmoX782UX7thyNitWTK1tj
X7Fv1UCOcPRqAEvvp3nmqec6irMSRKcxz3wp2iL8+y+nVBtmybjqnM5MmQX7yS5a
z77aXQMao8UMxilqdZbL8xy5BcSArqii8NSi0n2L8ONh55PsOYyzo8vTH2NNZVYj
oqNp5/Wwii9YmTA0UOzk+9jYgpfvEv9ZF3TDpS+LOPsI3fNLEJv69maVd3Cpf7o3
AuQhD2ksIqu2SM4VaKk1WJGtmBvRrsMf63SgsLBM558XFw9BeCk8UqBI/qSbTSF+
aoNqgjrGFjLmhJCX3TH1OrvfpDiVdceeGN5FB/FDDnOE54X69+AapoHmdGPODQNH
d2UKpYZ1oajV+Z6EI3U7wmglHWUo0/6Tw2lBhBrzkHadkQN0JRUsDIyu7v2aJj61
ad1Kc6RT/xE0ZOhfg8IDq3RG9H6ecmFNhmfIrXv6lU7T3HKkUVdi7l5YIpFjIEcP
laUc9p9RR86KuC9SIFpjtJ4z+PGwY2OhZvYw9rU5ydnQ0eSl5ONMzN9nm0omI6F2
XJq7uqeFxc6mum1zoYJes3k2RCUGvB/OtuNQkdVAnfoTJZAr994lR6qzTJjzIycI
OuGMVL3PMl15d3H1DDmunUpdhUse+97ExPx4Zwy7JxRog6uF6JnA/K0TdtChhDcX
hxI/wMNklTtpwSg1w187yA9hlbfNJWkFmhcsNSEOFmCVP7nbrA+VKGnT5EEdwKqq
Dafm3AZAZgFmytj0Ag1Obz10E4m7vKQXJEfsBL4+51CuuaBr4TULBG4ZJy14N9A9
yMtIqVxVnfwipm5o1GZv9ddTzcIIu+VYj9OCEJDIf6/W/+kfdKSUR/Pea2izAReR
7DWJ73BIzYJlued/rkQmeBzQkUnbgKittRWMA48v/tMG+D3ISlnDVvVmL5jHc+qi
pL5bnnsH6sieRIqtIWOT5hlJmOqwQ00n8T/aHmOB/5BKnyiu/TG5vlI5amd3kPMV
mGB30esEM7aQ6VN1/ENBMRyR1DVxOybt98imMTsQ0xbDopRWJW/ZRIYcHc2PZ823
4Sn7cL2lwbuWXJBLRETkMsabhvQgvYqAbRsNwFpx48XqFiolQ7VxSJmKq8TLbGI9
Vu0McM9vv1MqMxKqUeOgIZecMuGNwKKNRKZvUqvpW7eyQ+5g+q53T1AUJiVv88j5
0Axjp2v6rDoyZb5MCCGkQGzTpdoFI6aSUCg0MDNcwq/MZoMHvTZHxvghceiOg7Wy
4kmrS0axrvWBD+yksciHiERjbyrIsOjyTMUgmNwD8fJIZjBlfE8Q3zMm/m1vp+uY
eJRFyF1eFmcbtOvi17PDSSkfMQC7QYTyhfrHeMjpAvbs/Amt2hNsok8ACVZs9K97
xRxiB/4fCb7ZxMaCzeO/8rEbD8C4OWoBHZOgvqUcXhvffCEc0czW0vgtiXyIPF77
eI5S7WYAQU+rgP5Cy070wq0da8+oXyqSF2FclexrMa0gT5qWlPVsGnXgDjAg1xKg
CJL0+i6M0riHDGKW+ThOtyGTQJEuKnZSOMDS4oz8wiiLHbVzP05pw9BKyKhVDNZl
FgOjKKNgrBLGEojl29hZPw/e608T42zbP0v5gcE6Nba1fC5r/HCC5AGrTzddbaGp
o9I3hCCaR8UvjdZJzKGFJp7H43dExH0Ap1rtK/1Tej6a0metjCD6wyQGxkVwE2Pq
p5F/42LNSV91QUMCemNb/Lz/UwfCFIVULICXD0xvG8uLGaF/RDHWzuv3m3XnlBjQ
Rwl1xE9AUh8aJIhIyBhahs4FnsV5bFy2eqcVMJ2BMfOvqWrxkNoxZ8WLXtYMnXD5
Fx2scXmgkH6KuhGsUfkCIKmXWJEScnVc3LCw/STua/1cnv6ZAB6ORV0nhMNJUniU
OuTfcwlT+o0Ymve17+Uhj4bd9GBH45nYPRw1ZdCGoSpm+G0sdJORvI6nBN+i7lAK
CEwULqRfo3ivnaZP6dVTT0G29mAtCA8JbDZ3o6D4rLpm/fpuoZ3ZsgitJyILnSfC
iAc6HdmfQZB9SdMqhat1LiflAc+4ReBh+4m66G1V/Yg1W1/06QT9jtDs3sKeAhPj
ErEj2pHwoYS7sRzUpkxToioBLWqTlPElqAQP+3pYuAtwWWfFf9dJOtnrr1iSAA5a
Zt4mvV1m/xaqdA4u7imtFNyJbX2cy4Ed2KVHDytSt0WA1IOJyOVF3b2EDjaiMzdw
jIWzKM16lQf2hKYWeKuQ7eJdKm1qeEDSUnY3pHTq7V+GqAuaV3RAlWORIwvFR+u+
DyJu+OYFrGssGlF4kFsnRg5LogjOeF+NlX95SNRkSZ2Be8YqOnV/SHrCPr2fazYm
rNw8fXUcLE9rxwqc5Pw/LNK6UlpVLWiQ3bK2GKzarD+XeUGhetd4ntkj8Ye81IZN
CytadPFJOT7dnM5prXAW5ofMFTwDisflZEzTHYpTWFluogWV89UtsSBfmUlhqTdh
C13M56Su7EsPtl60qHQmYccLzn/6BjW7t0EBZ90AyMEYpbHvBnnz6QwH7ehT2G2Y
KFxHJFshEJf9RV6NqLPczaNBbDFqJKbzZ4cpf5zByGHdMIN9AXUuKpJt2DonQCKH
153yyRBcVc3kJM4hLrirhNT0EAYzMoc6yDWGfCX7hyv2CYQFZDaW4qWlGThAFjiJ
1FoBz//NUpRHkaL/AdM21ZJ2boRaTj9NtNKEBCZOhKvSkX0jiAslaS16g+NDpco4
SMCNWjv0jdYfVzTjzuYcHhi47rpSanyrX9oJFgOIp8Jz6xQJK7+yeSvU+dAN7zgv
iQKUUtosu1SDtj2H3LG3r7PMKuLiFZfo3jDoBPhwIhFMXtgN2Aw6YzFGlVWYq7kL
Cc+UUi6ZOx3rP5mM6SfWC4jLYEZHoi0Xh5B3d4TzWfbQFGPHo7QfsybnHBalssVr
gz5ZajqeXpenBM24m09ewWLD6byyRaYvlk+4ffvLV9r9+2yR3BsTxho1uRj18bJ5
o0la0yrpb8hmOIfiR7nFRf7QzGUjO5+LqrJj7KDmeb6eyRDU83uwH4uim1NXfTVD
TouS2VH9QFDUEhAYHCJmgKR4I8zKLWJBP6xH7FKR1CuCsEwIxqAqZUfeqX3CoW1s
7vDQc+g1uxqCefijZEdbwjz/+SeQXBHCq6e4O8fi4I+PbkDv+c/bijY2GkFsO8YO
IeBXyKHsLsomW8NEjmSUeo9Un0nA4LecxDd8JGR5DDoeXXLOD4W6oD+6IaGuwEhA
IbGP2lQDKi1B+aJdXDH8JwZ6+HtvuPBdtBakHFVXfOLu4nv6X2p4eI+KfMIAPpE3
F5ubMOcbM/av38taUsdGfsKNhIj7n+1sHgzxxZpto3bRmH2UmuO1BL205EUXQGak
E1pe5V7sfE22N6IXH75cA7CuuyOTRDBdYey+VajMNNgaoqQ2voooxoY6dYUSriPU
j1yu/odnkvuS/ubp6kOw4bMFeVD8jnkSjxfaiT/kpYdqXvif9V6w5tzgqnj009Oj
mFOEZXj9l+bj8HWZUguOw+JN4gzf38cmkbJpGA5XTtXvx4M0+aoqWEDM2bXFtAuf
XUlbbhW3UK2Y5Ne2pN6DKZ0aXaFi3J5Be2tjwwI1fjUt9+RMJODK0KlGt7G/AgX6
e5nvDClX4ndHqbE6BEkcszmO5cYRzdw8EgnMp418xWqacxYtHXeqzZTWcMSJ9BIV
8TrLsxOElS2BIGB79dNd56tuu/F/2Ap/ms30DSMDa9uFLp/yGFt7LWJgOhDDZMqc
M8h7XjX3++4NxCmWVHkUmUEfn5QPgIj/Cv8MB9yO6zp/gxtScr2jmUv3OZF2C3Se
QMR70oFtwV6rlz1cUIHtYSBLFeGPob6LhIvhBLWH81C0BhC1pIhWk0vpj4WSTYVd
89TVYn+BBuYdu/K8TYTft5c1Hgb9lULFYK2yRDpVJYKJUArNlD4xY5Z+cRKZYhmX
Qw/oIWDb3jiAiRoJxs8Mln/CngUYUSCroT2vhqcN/lJyWET/gq1Sykj/uC6vxr6U
0pTDnr83U24HWPEnBnESzZe+IxNgvXOrNHRB8PHXFrzWo8G0tE3Y3eWGqxMjX28q
/V9F0DVJ58H0XB+KA5lCJ3nG+sKpBrL8AVV8Pq8MfXHxlPa8fjQN2wX/L3g1lK04
iTKjolxIOdjkySQCKDfWy6hks4nii5y1D7WWdAC8AbU5QWXWjV0JVYejBlWZubUp
dzG+KwQCbQnGYVaKsQcvSkMe7T1KQv0EhdN/z6+SbTfHIMoqORUvaHY0HXTo3BB7
lvsfp5TMrgQzfjeSfJ8RCffz41y3lKfV74NM0bcsV2HZM2Tn7BMLFE3uUk4lNhii
Xzh5W2+JiC2VjgPRWiMdAhAdri/eHKSvO0N+7nY8uykdv28yxW/AP0yICAeyDsfC
qnXrH2FPw5TXPDOIgWIJ0j0VsKM8Kg1IkbBYBtX2ECTHIkwLNZfooU9gUNEMtm2+
czzgcKPSfwul7Kgt7L/15ARvIPLseIBFus/Ts/FOvrDMjPHU7sYqEOY7BlqVgC61
z2LKgK5WccHDWJpSCecZuZS+KZjATSMPdca6ngf8uA/0nSnRnl7AWreY2pjlf5eb
5SOMvEL4PUPKBfcyjkWfDOFwOA+H82hJoFTrydI6Ov4jcGZfX72y97D2b+wTmlyT
Uf2yJ8Ke/nbJ+5O8plj4jgu/Jqw+t422T4G755FEpSv429Af7GLf/IpYVwoEFIv+
wkGFFGoF1V0ppkxAjLAxkenCs+IFhCO+a46BkAfTd8IXkbPWp4urDo1AHoSlmXla
B8k3UiYvxOw/pj1RavXJj1tYmKXwzSLMWOo6+8JcgYDOiKrCk/vufBEIJ15hFgJK
dJ7l9/YyCVTzsHirWtmf5V5DQv34K52ly2iLW7jLlfTA1GR9qTviL6jS21JmWTCl
WAZkF9zxkSeEkdx1eRX112RcVHPzjBONB9mzyYv2559+ENCm8ebLSIiWq9MLJ1zZ
Fmbuu0PF1VAqtfNDP83BxhJs/BF7OdB64Md06YYV2Q9XTNYFcY/b6xGgmyEek8PO
fdrgJzxlLRxDuX6SDV3q3xCKGsM+j7t06qAgVkXeyHxg+NHKczGA2DIXiPf+PR+A
VR00+pp2mKgm3bCVYXNP4CEPr2L6KyoRQUBpONFe4eQ517nOht4aHu1aZrgTmAC1
3Vg/sE1OTm7bjmB2//eFEN6o59nlezw+svTfuQmGk7+iCgauhcAgWe74GmCkjOsF
tHufg6aHkkKT6eR4dDJiOFmU1F0veZupV5L+9CoESkoswhvrGrorEuc0FP8SyILQ
O5Ganqc50RxAAOyYgl0jGhi7/LuqGwUHsCAG8RFyEN0JP6C/ZlyW/GzAm5N4/0ws
p2xn23OGTbxn+AIN7zE+//LY+rEBPp4s/KIoOYD55apmyIqBX8ZUd9FNMddn3b3u
NPD2re7xmkDKujr1Yxa2LVNbFdBBbFGWOAEkZXU20TX5+jfN2PJjMu5WsO5h0v0l
Z0fRYXZvyVYjKNS7w6ZoZ0N7qh62onyeaJ60y+NqyjJerj302vTfDv/si9h/tkDK
eZ3TCJdwjY2zSibxosBLkcC15PGXI5FCZUu3B5uWA6/fM9Y5Tf5ELVFZPfkWrr9n
FmZlq3f5WOqxKl7dT+9O9qrcouKFbpEQ8N0rFZVrHdbZVrSxEAjVcxYb1514Zg5k
gye3xDF9ckzb2RhZPBLq0YO1wU7LOu4OJFvytNC8Fp6FGnQGWFQrJtKEj4hTf5LI
pt5b1sbozyljo/535AremR6mZW/KG8y/j4LWMScKKeBdxF2XQ8WoKCAZKw0EAsU1
Zx9pe4aQLQ2ir2a4jmvdy/8PumOztVCD3wU8UGp/yT4a3GQuA9twHMpZcqbJ9g0D
g9/4ebQa4reUBCleASHcKnzp/uzTxUW9W19sQcLp+OxI+7Rto2AdVWFNUiB90+Tz
zh69OdurTdckowH5DaDNi5MnZd7FACAymySdEJQGXqjlDe3ZaYDmGhdwzubBLrB+
DD67Oqeog/41n5TGrsgleqvAZtg4THKCZlcF4kOHnUr9UtWSSp5w6W5GICUQS44D
F0ixTi89BcuPrh7+hvP8+4WH2kTKA8LiTLjjm+kR5Ws5Rr3Piywgpcm6UlN7w8Cm
VOjFafNfXNOFOFfeZG1WBfF14pfsnjqPWIlkCvQp+gKhaWSHcAH9aH23s5KY9Xbe
CALOUfh0BWQXs90hpTLUUFWL3x6XK6iBcGbuqVhgPzsATv4OndcyGce7p6TixB6O
Erf/IENfBx54QvicMsk1jGh78NfpGSPyN45denHLUDcOevoHBagorfeZH25eHjBX
d6YhsLCFMkPvITK5DSJr3ntuB0LoauhIzPL490OfQM2VUMGZNPY32ZG3LbszoBTz
ASjjJfCRb1Ts2HwvpGfCkOf6rqgnaZlU9R0TWPJzwhjyuAIPNMwvIkhFKdvJV5Xc
0hVCgLieVI8Wgbe/hd9B2jivLwcAHwSXqgg/cMy1oeJB6JK2XeYU72qocsDPPeNW
Ug/5ng/5RwFKRFmPaz8McL6njGRA7hXUrzMxmSgt7RXJf2aeA50qI+eRggKMtiZU
f0tX+MGiVfzCTJ4eCP/1BdMkYg3siDImjfPCGYCUCWg8p/vHzhAT77z5laAFdOzb
9P17DeG6MH+nw8v6pjh9aTzJtO2hJHEFNNJR9ZeWKjFmsNwrn7aqoCIyVMNlJUF5
Pp/jOUTXHTuuub1PiN0X7XX5mi6fDf+HlPi2QHf0PV84hp9E2w6azpjXaRqHzDaW
XtEsRZ5h44WODb70Nerbs65tWHdo9/w5WFnNSUxs4Ja0+UAReSfKHq6hbDmFMO17
HaryQjgdAGbgcGX9F16R5VWLQOwsqfrUA2pDReHY6gkvHnf6CEYKfonBaObp+20j
o13A8bEbyX3ZSGI0CMoG9TcpNRBmQOqhrLNHZSfXdIIcJIBYZQdvrTC6VEc9atva
ipLZR4GIxvi5Kp1IZCbUj4Tk6NxIbcvWm77TePAcCQol2gOUz7jQs6aWxjWxJTrw
kF8KYeSyW1+KwtvWeGxPcQRe+28+I1w9N9dCuWfh0Cd9pCib+xHeaegkD1aD19s9
+iYeq9noJkMd0dyH19iFXvMLy26itlUucSi8fH4bq6pvlgG6yHyquBsUdcvP589m
ADA1qBS465fPYaey+hHwbishXuQ7DpcFwsPlb4SqZO3z5PAQMPYdPPE/lrSkCvmx
hpJQrCHd9Psp1jFaATUmSNQZ6bq3j1ro/4qncNTWd9ofpLrcgtslebCWXW62rj8j
q2ybiww3SuzofjzQf0qCISY8bsdk1yfNCYXKrqAn+8UTb81UHu/HOyyC6UF/N7rW
af6QLiMfMt80ZRgS6fvuFiF4Je1wiQ5swV/BacqkRCntAikkJmXNOzwcBk5Nj1l4
Dfru5dDd7qhlgF5e1an+fHbhapfE2NlB7Z0XOimcC2hIsh44vbvT0Z6uDfGGI/2j
d5zRRAq5s/ITBgO1LrJQy1mvwkMD+R5SA0dnDnCO5eKDmaD90WKeld4Uiu3NCEOy
zCieMMFhtRxHLvUK8oCO5Kczw4+xyk9WOK9xJJV6bpBgrYuOWHEdxc9KBWtzFsyH
UGoguOK59rVC56CbiOkqJUcttgd2kOKqHLo8dUKpT3MQdBvxUUT/ybMpSWrs/gqK
sfU34y0H1/JFkHT7PKP+4UqFaFby2qsCuMUszZZFfQkxUDeIXjjhf8ze27OBAGWf
5xBZDn+/kAwk5WXHYkg0u9oUZ69CAOCS1uIpny/TkMSVV3hFemXfuuA7rw3bH4Uh
YvwcdWVLqIT7SVaQiB5vzW7Ka4rh4YchqWNS5JBklhQqSjzwopWRSbeMFfHLlFOB
h2U6bt/zuDWcbc7umnf1Z5CXBc2XlMWekhBOZhEkC27nkhzFkJ2oTNCShfXUYmsX
yyrRj97ztsnOK+GqcOTx/OFlcF2cwwOBMf+d99quQKX5kB3qXgjIvnhkh2PwEZOm
i6kKVZgRGXVs32RvMborawKWxAQSnEO1aezoIxbMyLKUil6ygLUVkRZXKeHmxs+Y
YlbZ/EMAmKV+JV3iNbQ9ME4kuuEbcuc982yRyctbe21BgwVP9EeJIS52JH/RTsAW
zqpd00lIPqwwLdGEVYZRLB1TmCR6eQj6zcqwOmO2AFExGHJSkPUmrLY6yt41Jg9I
YrVopdZDsS1A0pBQPNudKpoWn/4uKn3QNkt0s4A22vGnbRhp2wSa9rtwOM4yMBpH
af2a1+HQ/RQJy/Lw8+mzNWAJAdX6aug7YOxO4+5ETZI1lNVoTVaNSPj+RjJipGP7
NiUz7fytzRejoh6+ex0BU/x9kzJ+KPnBJ2tEMk0pHsHvMznV9Y2da8TuJU00Yfal
NVxU11qPaI8NNO/ieqX2ORunTJfNTPtJd5ez021lzkC7pi/gdDX6zIvUcty5I+zA
rpnL/f9G9sRGh7V7ZXizV8lBEtv5poecw4istGpovTP3Z8p74Pasyg1Gm57883gq
gH27EXfHMhCirlmasHykSuoj/k1VWsDgd+ObdG74PPfHtutash7t5FSQShYyrT65
PUA18PsOwPj7N71F5wJreKkoUENfLGmCELlbb3EIwWAWhrZIUiXYQX6SL1NyXl0p
nbXKkfB2Uy4wMr1TRv3dyOCe2tehYfbLRHSk4LQgyrm8efixADaMOhEdfgf6m/t7
OrnegGkng852Hy/nrpv2kVpfp0EVenc/eUSnoRMb3EF10reAAKS+c89Uh12sQZxC
D4gadMV+J+SlgngsE5KRiSouojKkiCBo/HwUnfi2NgjNURpCYmeBxrs4pI+lAMT7
dptgGtxQc7Loe3gX7pvv55AHvcvsy+yo6s7YHsrNv3JCHzzmFAkn80DARGX2o93x
7fF5y2J4eDvRmEbfhM6jkp23DMJeab1jURF8zhpwbHbk7kOz1DkW2/1HlgCoMOmC
up/e6FbdbXZYL4/0h1MGUHYKG6QcUj7xbREoRkF8AyB6zNkLN/qRqzB2jNHoI26f
zq1KjQwykY+q68VHIpZ3Ni1np+MFdeQm3nFMZEBvR17MEOn3/6fn5aIh9fSGajTh
z/IBG9yz5VDXzwzjVqOj+kYhO3PJxLTXdTUqbIFpfesCpfCCKC4FJucs1nRYunVc
JfL8byg7tfuqodL10Wv/ZnemOYVApMb8caQFJjYapjLAMqWVOm2ldkvq1NYV80Nm
9K0+WO4huV5MQCqOmJ8s8tLBjpIOUjyJq+rVOE0MVntP8A5MfqrUsLQNx4VHzHzH
7CdwdhcH4SxHTZRypDRN6yZe1waGwdpOYGbrZF7Cmmxo1sLKi/ZKqBpxm7k1E74d
H8P6X3GmTxfvxA2cBC3QyJ2xA5TY8WS55ykT62sF9kfgKBqj43aG+Qnq+YasEO3P
/zxwivoQZKnq5ByAIWc8S52DA8U5MinavFp5NU2WHB2g0aAHu8m6F3bzJ8lpkEzm
K4U0bWPjXBl3eH84XRzr2uA8Q7jbLG3BTjlUkpEOpau6+mIriALfZiYgVjSPFXbV
qkQu7KA8vzECGdo7ehnZTCXYHXQGdNsMyGyzlR6yJ3DpFGplXmZjDt3FkBHGQxtx
LfitXGa763BtbhRGRu6Y94nhrIbw25tmuTnButbSP2pR4F14dly/ub02sYETj/Ta
GXMo70QlT+itBWTGVSC+hc5XFnWcPELrP3jtcEtl8nFTjYKd1TmgXLtJDdRhg0Ot
zrtDEqdhd3K+hFsqpyvtndky0goSRndcukKVTMvp2DFgsGiYinh9QkDaN4IWQJQE
8vGDalnp4KQp4uC4gdz5CD/cXV4rcL/x3B0WmjTNepmoF6lX2Hpxv2E8Hh7h3MUD
csjwIoeNOND+ALF/SwCMLjxy3iqcCEnQwxOqL9Pz9vJvV2DQQ4JBDHKMmpYQqTIm
voj/Obnkm4qv0wN8X6a7rOnPZi23dAd7xU3i66nbM0JPgkvjs6yG8sEUpJfBXpcj
+OpdjJLc1lU27twUlclrypqF2GDZAxmcob02hGCxZjYqD8tJ7maghQEeOo4phpaM
CroPCy2+XyargBjsLJ/o3aF4MbGjf4Y2fL5R5sX+Sjq8mtuaLD0f5A84tTRso4gM
uX/R9hHg3KUjLZIJAT0eCVgrSFCz0WdyL0mvoWZUxQtWA601xx+4xOTOtHhmMlHD
Yu4ZO5cyXjM9d7MmZGMOR5XPgrkxE8+uKgAI7qEZUQaZk4vmw3rq/fcflF9I+us2
YUnrgiIkt/Q4tmR29NXT5D0it58qcLKOuPhEsnl9htbp745oEn8D/QqsQqUmkgHk
CjRfA9meuWkOrmth6LWiiK4aa/NOP3KRd49KhiiBqCo7pfdLq8YIpsoidzOMxFQY
2tyvrvUl1NU9SdUySK8OXQEfoiR/wi1anQwQ5gBb7VXFYUNF1cIKFD1DgiMtXflT
qtfC3JzwnukCMSerOR5h1zs9NAzW74/l58cpG+OTwFZ2EC3tsjAxI0ykpaDGDufA
p/u+XuIdGVHjJR7DZpaS7+c8gfFFjPkbB4oQV5fYmpOm930hMKJbejB6zyAroDeN
VT11L8EpsAkIKt7Rn6SUsPTwyLnytTdo9x21qvbG+pBrbyKNqP6vLQODoF7RtN5Q
yHiBr07EJlhcijidpZ8kyRr7XKCy1Uoel35MdBEmr8YeLKuXRrnYwUu5BF12setQ
Di3COnhLhQPoOdboABAzO/Va5hBmWa1VLZya0krTqe0/CqaW/qVGdq1fJq+cRb1P
7oAiNqI6yPAwTmbykL653drAaCLsFl+4FKg0i5EPAQuvvgMa8ns8vbx6DVDSbnPP
UUlwCDQ/ccYAo3/QrKBrM9wTJPZ/hqPuk/ULc0R6iDWBK6El3meIFsJfnKhZ0s/Q
ogThq4YlOZv+m1h81PbNn/PKPynzybo3dQd+T/wye1Ob1TGk2P0UfnxbnoVgQTtp
a9euP7/iOGXrw6IwLvswojkbQYDb5I6l4voC5TgooLImH+OzBV5EPlEbqpioIY6o
PWzX4Fuqk9Y25nNudrm/vLnW7dtw+tqbSiDjRXI91JaVDoyaMbbyvOXGwoWzbTSy
sxcdnwrjFQcH6+7qHYA3efUnkBLMRV9hxGumnNUt7TM0P+LaKKuKTr7YDH+6280E
yNN3EiMKWU32ADqSO/Bzq3X7+CwVp9fpAdoJoa76Xe2cBxliIObXk+8at0VZjvti
xuuH0PK1CcH2CRFxvN3klOyu9RDdy9ey4HXumzojHvrGnW3iJUNzkJ9iTehUTyez
Q5tYfUetyKalqDfEjDmKgNXZQNgleRmN2BXj9XP1fF6LQPmCStCRN9OKoenOG7lp
4XiIu9RIhhRQkKT+WWIp/T6Shy+BKp7yLteozvRfO5Y30dRXbRRVQn8SPe3aKEKS
vo3U24pFIsmbZ4guuhCpsYolr/8GU5etuJhIJwrYv5AY7AQ31DoYvYiZd5NfEmfr
SxN4/XeM4XakILHzvPUwKFpHZvEyZGV+/bhuFF4VR2fVlZUpxBIkg3AjTdI5WOxG
QHmS4MyNfGCS2X8e2hGMHKtA5SPjq7D/ZD474o7amt7CY9xIc0vXLzzHeUzU5Tur
h9jJiMmQgqYRxVv87/LSRBdIdpeTs/0uL8yfR8LY63Dv/SItwQs9PmKjW0jmQixC
GArrWT2zXMbMOBFVMTI1x0wueFEMFnAFCSBzfOAI0WWkpkUI7hg2nFLDCX88wcjj
9ANj2vwt8xQ+guejg4KTvrJXc45XU6BmSl+l+dQ8WVro21YXeRVXo2gODIYSbLN8
ixZfSCYjwHkrCSQs4X/t0ozSlyALP/1Cr3Zpok8/pgvPIcRPgTg2OR7qM4TsiGaX
qNu6bC4d8Z2ZiXCRyVdA610WjdoeBNlqZRjlO+0BrvGbVg0xBd35nxWOwaeAHPg2
3QeQTi4l/7/Os914SvDiCi0kAXlkPaHPhNoJ31VLSflDGLRqDndJbFXbsNjKjzJE
eGy1tyPg2xekEwDVESHfU+GAY7iPyMfCBmFyiGp+GfGHGA5pdNjfbxzjO0tXDcHQ
DrZ6qTI2TxEIlp1x5n2hukZvsmPwhdWmvGZCLsEPrKUYb4vfjwWMopLRwr4I7u1S
A8dQyX/WIxiGmLBkhkHSTuPVcSJ2a8QTGR0I15/zabsT5KRfmjxefQvUSxdrwiz1
64lCcQtpIDjJYbJ6ZYU02W/3jNcvT9l4GUuPd2rwd02of8Ap7QQ5n4QxKOAP+aZP
hBX0HGEbmryccfINM5qgX6QULfrETwxmObOrRmHpvu70sh0WQ6FMMERgkvhujgPW
F7UZjdsgp+qcwX3dQjTbAEKi9gmWiCI7Ljjg/nAUOZCVU5joe1C/wVf3qUFOoxr4
vGYykJeISn5Kuf4KW/TXRY92rJkUZqRlXIka3z9e5v3L72YOzhtyTjhOjlJN/8De
xbeNiAFCOsZNnNDST5uSxRsyDUgj2opF2doWeR2dY2CEzjLjoh7WbK+UIMBDa2U2
dE+kJ09pwREmQB6DgKJSbn4P6QrDIHwBk87pdxtGLwcFZDiG9dz8vxUfU9ZUEeRk
W+7eDmA7g0JYQfYy+77bjoHIK8SIaok3zZMagsRKcfJFZiz0sDScPL2a1+MWj13S
vEB5cAsn7pKRKhZ5ygLtnFaZijyRXke6181DG/Lp0IohurqHVtSDPi7P8oecyES4
8XzwSentBW5PDbMJ+RAsn75knI3aR2c5rnuizgiYZ2nfJ57h5t3uodXFFT1ET3Rs
FBoYkMcagJfoPIcg7H75Vns0Vz1b4PrzHdlndIAdaqcGx433AO31U5kxquJr8TdB
PuIQOiJ2VCs98Qwv5V3WfizhwDYHA8rtvXPebpSXXPtErJUJ+FKGHNXLiggFshst
gZoZC2s/5omKebj9EgI4KvTefvsBy3aOP7CA3oDGWZIwyn0Sl+hqvF0H3kvWKM17
V/qQBM+QS3Ldjf8hPW4OQbQ709uLMpXX7sPh3Ta4TZleDE3yQS4SvN6QTd99Uc/F
R9Hb2MW4VfLdEsMwJ+zifK62/dLPmK2vy+PC5MLL5YERnlfqWDBW3nGFew5uxZY3
27BeVW/Uras1i5YVVSONfPnX0a5oXof4CPPe3aWeJLMc9incv0tH0WNlUsyolQK2
ONV9I2elgf2uAv56WDtxk8woJGJaZbK6rCpBdKEH+RYLwsBQXLeeo/tkKDJHNwmX
27pVWlL4pfnaLZVHPUcLSQTtLPq+0zWT5zuxQ8nzXsPUSfV2NKbUyErKkSp28ei5
5JOYlfpBmdLPJfHqu3jDhR8TECoTjji/wPz8sWNA191OqmQ65FyVXhAfBHGD/qJW
R2BPlLq9P9Qfb8OHPFPJ2UrWoYnQotFu0PIx1dJ+MdzsdEVnVE2dVYS1qAR05n+K
s9FsJ737JuFwtNdKhBfxM8cm0kTsGTFlJP0cojBU8HbpsaS18BO+xNrRX/aiCGMx
ev3JClr6TQDSbeN7B+CjPOO30cYs27qb6yzF3eXsBMY/hVrz+a+dyDif7BBLHlRw
VbYD0PZ8OEZrleHHEuc9TaA62V6ehKwgFqD8lAoGctfnZ1cNYmhaCCfgUvHNU4c5
gAtmta0tTshXHZ/e0VzI2mSlfFYAHVm58kNVjCq20BBA9jxCmCuALkiMgxahnByf
9iL3uVIHZSF9FOrjO5B8uzuWRnGEUMrGxNutejGAwXvu+lNpmYvngw2PFpCr/0/5
tufjvxS7JC+Be2fJm65ibAMAag4+2BQQfHExHFF+A9qZLfu4N99tsGnuLZ2VG/kh
pZ5Cwvr3MLC3kUyip87Eu753yy+vig6PUK0zJeNVI/PXdi2A67e7lqtqhL1dWg+L
HCbq/ZGhDhyEVeqg2fVZf1Z91yZeXo2HxPwR4mGVf6izax4mtwuHcCxX5VIQtmgf
LtdLoBi8Q3akghuUCOKPJN4zpKw3sNfN7g6PMfyh+LKgeRtwld0p6K4OnpD/3S1t
xSrEfNekDe7IZra8s39dDH0oG+6QyQYfErw7IvvGQCGr24BnCYNwrFYeGc4I1HWm
9TIybxxm8QKjzzEIS/OlTM0D8OeSDPB5U/TOGznwHodURuIO/khv5ypCwY33wkwv
VnO6djX1VHq/AVYqtHOK07EmG1P4ifRKJxCxgMOS6rVmgwqnoORt4gqyCg65njKQ
z4mt7ugtyy34FZQdW7/5mHIkNNpDdQDgmwJcyr3v6cHCaZuxvIMQqNWbprvcuwyw
+c1ZFSitMtmS955k8v6xGpasCfWaisIN2pSUCMFN8yYBxdW3FjRpbKWkRAWJLzXK
5uIgM8Fn8rwpBh7CO7Hr+xbwx7W3DSDtLvMppOGAKvtMCUCIwsanFYpj/GgyXv1R
XjZSDlaneRbaeyYj3kpRtOKVSk8vyVurU2IY5QAWVGQmwXC1AvqhRxo7zg3+kK1b
XVV8aTD7BEIYGL4H/eN7qXZAGyEJD82yq8aDCrdMiVKvMzB4v6X+88jRU3/hwyxY
VtSoHqaPNhb12jCrDBwhQrK/+UlExlss0KSN9DrQBIM+dcO+CWvXE+HFDxfuV//N
ho9aUgOPcvsLXMxV54SoGuq1cEIIzU5N3OTGrDQmIvYIx9LzY/REGBSJD/OE4t8a
wAHXz3rec9W3K7tYGBTijn0rhOjhjh5EHZk5cw/xNaBJehoDAcGT4Y3+g/Vp1Z1m
HhXw4Bkh+SuZL/1Rh+mjr+QZB+OUY053ll+aTxRa9XbP/u6yFZZ6RGuBTebuM0bD
QhFCWQsfNCZxZWaiJ0JMkrWVXgfMzQCxgBeLGsLK3v6MFbr18cz9LMEzmnZZ4ckO
JCnEC2fyXBBHzaotfk6MimnOZ54iDDX9MP+irUFqFWIeuq8IGyUg/1o+SkwxyUrS
lehYDZ2MypUzxYEuGZfT2nlD9f2eL/IQD0OzTQ0ZSeusrx5TbcZsEFrHH1Q01yoN
r0F6ua3FRQKmfr3fbpL4zXURwIEhEMZA/uG6M8Z7nbvPiRz1pSYN2vTuPIZHnJZh
e71X1qQgfZpEA0iTxbuqi55AnPAArQKM9snd2H86lEZ0K7lUcksQLVys694+GmbM
Kuh7t4aaQP+Dp+tPES49ppFwLnSK2ruRnCXWNeNjrFYrnbqM7vhAElon30Q5ELIW
Xxcfv8sa60h4Q9pwO17I+yIvqFe1L86BxhDAIzBUTG/mWRB8I0q1s0tfDIcMfDQa
9ebTpWLMibgplS9aflNNDjeJV3LokREYLYBKPgZhZAh9L+XeD9o58A4Q26aN1yPg
Yrm2QWUdl4SslJ9jHETn8oIUg1EokD+LxXbKLVgIhJ5yYUZHIe3VBdwc/0cizrft
NT5SliY6x6d8SxhAfu1sOH1uOQP6NF/fXZOiOPBKjl/pCBP96KxB3ohvSHfqHi5Z
ut9J1l9A/Dfm1IMJJivsr+T+j/sqyFWIytXK0DVWQUM40b2RA/fkOwtu4EnXnzsP
5iUYRFnRcv9s9GlzhT1XLjn+KOEbDmfWzv5wcPlzUg1gmCvmgwVSc2KdhqLus6nl
Cz15w5MpDiRZbmlTJC3Zb76aYRUVaS4og6tDr4VioDFBo3lSTpcTl7ATXpTmFzOK
O8AvUSZRPhDn/0dh92PPOdlUwngoI9r99LcolQ7ITZWSxBIsVEWQMd2U4F+/3JUL
VPvyQL3oQCRJJQO7pt+MozLz5dFH2wRml5pa60Qyi3bQox1mUEZfUvSHMZj5SEdj
LhPYYCvr6n1WXlNDwGPjUTI454C828JF5D0RvncfyI2bGOx/+TOs8HXJbDDfIv6z
lbsDeGdc3SLIB4uDuSeBOu4jjDzMWpU3JS13mLP5GpbPjYiAPTINVILz1tBhepKO
RHQebXMzd9EPYigk//kJjlc7ocBHM+icM3GPa9Qg17+c6la3GiaI6IYFGo2xpZKg
SaWs3+LQlYnp9PNub0UTpg3vSnkkwakkvntJE7zpCGoStY4sFV7giFG9CVlLqLYS
dunLU7oIFjJo5EbW0y2zt4r3gUWEuhBrB7pt2T3w7BMgrnsxa75pchpM9ygJnP8K
eo505slfT4VUYr2XN0GddQiM15B3Dh0euVfj+Ow/vkhxEpy1M+PxJh1ddltBi57M
GkhYnnhhLysHD0RnB17CDz4hIl3IsxWHptD2bcMhyHmFd/luh1iE0HjkvKJBagFk
1Nzu/FRZ5zTZW9ZCPu5qjh6n7G9cPLnWnQkAQFqbPTmI8pFd51Ts2+ozAGpY7Qdh
HiJGT0BgbN4qyMpxBDd/StH0IPM9OmJKc8w/7b6rAaECfzu9BDN+zU8yA1Eme+Ei
JB3HCyY5P3/g0pEv+tPIKjYHe+H2VMBNx2j18y3EVCsVUq8yBqdbaV1KJxKa2Jk1
D1ahYU0l2tMPcUl/e6n+uQKDbWVmKfWIIGg7U0gnuINT1NQLPNx2EYirmkQaESns
Sko3Q2e7O84lBD8WPfNKCBOyJdke3llwYsG8pKXY5O4BNA03t+aF7GEdcPYoFaZf
TT8MZodYTXCQi39jzuE9rJDmwA3AKa6F0jFjUs4V0AkS6uWsqB1x9D5R3kDwKl8X
yMkJPInUwWusNrK9ml72FEZaSjEyfKSQqEwxqQJ3nZ0hPACTegBUfrV82sM8IdOV
Pe3/vk5GnXBzklJUF2SEHEXd5kjJUOy0yd4/Rd5uUxhMF0c9c21pgRzgqiT7kCCr
oO48r13wcOziRqpo32Q0n45cpfWKCmyPsRyfX/CDWSd/RPH/bTRLHB4pZpJB/FbH
TyXgedwkySAB5Tcno4R92bUqpec/tVObJl7JJVDWgirLmjpkzkG/10i9KJjayWK+
WXnAEMT2mvLvi5PlnUH/1qtA/6aSzq6vM2IX3tuJllVOj+g9yozS9HHcUCipzUfH
8C1TI5I2dMfvSX6ILk6ZqwEfC9rYehJL6LgTog8txA91qWFjIhW3OuEOp2+bK7vE
saSemAw59H3THbaeHmdchX8swqX5DfR0uo6FLrMnKpKRj45kVcaC3hGTt9SBz2kC
zzL93z101D8je+LsTjnEIt2pVmazR0RnRpi4RZ09uqpuhoEnQJwQYtSMatOgYbLY
a0eYswmlo2Q99dPu/z0sW80kJCqmIv+RSu8ajjuaqgNEtAYn4+3CaMDuyN/oSdX9
lGZjn9c7BTFqBbpm0PnHtVrmqETnLBOiD6hjIAYbde8q2C1n4T1d0r/TxleSTzYB
1Vyosw8nsg6FsmYziDlsaTe75VQylKDIB3oPny7bvqIkpm0zRtQzvBJ9SPWniPTv
c3lmB6oOdLQH3fUkQvMeVR4C7jgpJMpr/ljVVDDe2+6+oy6/VVdB25jX7KZ+O8/i
SbHny8i9gODOeSoZPmO2MkZY6JJYIuwjjPTIuqce88crwQse+EcXju1xXyoV7AeH
xAn4ERFxRPbR4p8meNA4QLZLtEpTzoCjhZZwPurGKpN2UhcXazwrpZ31bG4FrUiV
4YAWh1tvCewUaqTVv5gwhoHq0PJ75eRqMoHqauA2t5/P1B9s/gyCoGccT3heAFbw
rS/C4yeHbp818dkdAdcOPo8X4WbM4UK+c9bEqAexqV0289FO7NpZ1WLpxN0dei3z
cNwIRCpeF/+XGgEU2FnDF4lD1kvxFk4aDYYGHxBRJZrxTfkMmUMzunZkdY8Ypb2d
+nMfH6TutAE+VB5T2ps82rdfvYQVtBdzQdC0poB8SLHSF6NJPHkaLZ5APMFoElXy
Euc7wI0HDC6/bTlS6aPg3dlUjemcRhVmoynQ/iLABT944G1dgbOJnKPcV4I49MoR
YTizNgXF7286lk8YrcwpeMW28Ea2tyO+9UL03HWMpuM9OWvnPr+Dj/u+OxhOYJ4a
ZHGqkWfoz9oy5aSP6We9MZPyYpPVYTx1y/KWhWK23J8Ggp8TKNDdlp+SAJFxAwz4
IYkn68XCKWmp0dQ71uel7MRtDlH1jWECVz8SEzFgPf0/s7OtZqfL4Au4+HUBPJcR
xSspceleU0dfBawpiimIjbOk5q8umgLHiyPLfFGCeR4+kMWMmpt8uoWQFft0EF6F
BQydBtlH/nEWq1FOVn4xxJPz8Lg1BMuUG0NSgFG6XCGuVnHeXH/ftJV/Yhpc8NNF
BmG538tz5LWbIdk6oA8h8sLhMy4G/W4G4EkQuR2pJ0+JQvHo13T3Xmtbf/UAyU3j
iXKEs+cuSvV5Zg5iErKE2E/3FIoZOWiIv1zCkS+jR1z2sVGFpJxTlfYiMXWDzcd8
gqdy8B4y+nUjluFEaGUXTzNJfU0Bhezidt1v0nM30mclrgQ5e5+fBYxy3JNmsrFC
Nf+9KhTpl2EHOdyGo6jytCptOAwfNJPxbnL43Mkg1jzLoDxgo0s9on35BXJ9DqSn
GETYb9CtFD+ph7ay/VXF4+V29D5ZyBmdewZ6uH9p0fYJc3JKHIiypzTJbVJ9wlEX
6tVY34n2rFQJNK7EPeGsFxD7T3AAMWjYB7YHqUvpF6WDiTEF58h78LNWiox+3gzs
Y3mBqqmCZ7YDWR1DhgMapL8QoYPiUbPoda0esC0GuekHAWG9ekLrNxA7HaDw6C5G
eYmxsYXzP1gDsfRRLljdn8fufRlrZbFA6Kza+IbdXU83GvuCo64yqZeAsKXxI5Ol
6ECpSVtuiZHGsO+DxQG+0ynC0sqyn5OMwxwa71eutgT1HMp0UQPFa6HS2nwSxG9M
m6fuP2/aldopbAQORXRIE/RU1xsnln7WwCKb++1Und5BYSDIGIgQgVb+jrFNqHY4
ORlThNsxx1O9pbfmIrW2pDbEfwNMMghcyqgcJMi+t7I/uUnKYFgyfT7LnV6Eyt1z
hLLus9SCZlulN6p7wBPlZG+Tn+GsMo5MmHyr22LSeBmfBf7ZAcNq0R7fAKHqz/69
Z0hD6qVxCVLIwy9LE+PLQg1fhWOCwymPWl46Mlv3VwGCnCun87D0hcXzrr2zJyOH
82r4lgp2eZjsZ/laLO8WBWanqaglW71f9OwGP8i8UA9MbcMwnT5jchBZ+HSpran4
+Pxppf0L3/WqKCBYIkUfSKm/iUU5FuLanj1JXfSgQgTRlGpTRpm25TkMFd0sS+bC
SwXE+dLmX+9rna9xFvzMoPoYKRVv7QNUONqNXobdlH2WkXRbBL2NK9OXDF3YoG0n
yBUSs2dQlvl9UWuV+7DzVAsw8CGf/maRZWYlkTd4PCPGAboe+6Bwtzj4WuUz3eEc
ckHQd7K7iZXcR85FnRAju9ZggjJe23rrkkzaEvGA2wjS/OmYCnivyLdF1t19AILw
NeaAUEM42p0Im5uq96hquCoVxBlK7a7UkujA1Ig56uophAq6x8aB+vlt9GSK/MAr
TpgYgrpZg1FXXzDpbBu3539lpfUaNYnoEwR2O3UDGMdSBtsszAWAWjaeNBuRJZJx
/DPEdeFaZnd9SMKU5qIEhmBURn/AZAESjAvq5wEoyc6KBj+7lByD/Tvu9ERaHuyA
9X6X35IbIqjGQ3eFURPD33kB73QJnRdUcERQzAp1TgwTZE0p/pi9CMJEkhs4qfF7
0T56yIUgM9E+DVjMeRgc0KYkEIMFCMjVVLObfKnTtN5Tkj0hTHR/4lwTLCx0v4hH
eE1lJRf9ty5yvjDnDhYSDKoexgsy4I7PpwEwk2gSPONnOaunYH4IjOOOoPBhwQOC
RRxKMVbkBxzv+40GwyWwq8w8ejrQGZ4VpU+K6xpr3Qt+kApXL6om32335CuvE/Uu
jvcpxjy6jDFM+ftSQpGzCkHZYa5j9rcEsdzhzRw18uDlUOCTJ2MNsKIxKtK22X5h
rkSCBQE/kdHmwu8Tb1F9sTjKqZYJlCeszoOZ6fVK3EJacD0b4IIfwzZT/u8KFCGt
RNb/Aq8y282jskoDoaKFVhiYyqx0Ceba8xcAgeOr3FxQafasHHA2xXQyU6foxfgp
MrqXTXNJpNlCQSFRUPVPzk43rV2Gx1xioqBQs8HNUQdTGTgaq+BF/IGIEQlhvF/5
MORM4GcuEjaMstLUyy2jiWyibfihuPHrgBCO2jM/gJ2Q6HRCoPMoPR6r3zX4ZcMJ
42AOptmsqYfjsn8/BIASj7YMFAe7TU0ZUWj2ssExEbNY0viCYtU6nkkEKjUr+BrA
8mIL8GgJdyvXpwe86LJwZClJipvp00QYq1LvjRSbkcknpyd3CD/cSm/47Bq/yOKT
cod3OBaGw5LBMpdkCASwZbswkRfRl3jZIsDkg+nlr3BZ7mog911pkjBV/Dho6UBo
fwZHhmJbU1/7NhdmnYWIrkpbxedN9rPXcNyidcpNmtZKXWlhYw9ABpxJHyNCYOjN
ZaH4e8b5wVB904qvPgFNYrTCFb9NX5fdP4nUuA5o0q1+48hK1zXlosgE8icvwJmL
h9THU9YZ7ExqKAnWs5jKqEkCdaCbunh1Gr15NuWR5hazJH2zjAC6ZwL7jg7qwYXi
a1mK5Y2pVzFufMjU880zjK9FdNOfxwi+J3rAwrldo36w14N61rO3y8R+oMXz1xm7
KnmwWEZD7OxNW1GdF0kiM2qU8vbPxTcMzoFIEjsdjAGT7pRJm1WEo3taV+xA6uhS
3CnDflaikKmbTtJIuVGEfVaA0CYtR2d4SiZxP9KsyNZ4iclUX/AjJVSij8jpfria
XmtjprtKlqlJMyAm+9IpYHnm1ONLAVCpf2yiO2JMqeWsagsJY4sTIeigkhgFi9Xe
iSLByiE+pGyKsH7/GcwoD672VYCP6bS9sy4PMdzCktqC2B3l1PnHCmPkHGjFaRjy
NRcN6xOcMuoQXl2XAIzDYYV7UXNXIJa3rpSre5aslSz7aDindxlBDQq/k+kC6Wk8
jtOkYz34Qifqec9nwRssB8qsRvfNWVkgM9mJkL0fiOvwuFFKqeF8Fo7PxRXl2fD1
VWDSC8PPRqIxB0HiLRhrz48nQp0XM/RkauzTUgKaSNG5KtSE+OBvanamFrZTVK2s
mA4Q5ehQ1Vd/eUS0fOKhSQ8i+dIqj3uK22YWXwNL2yqyg5GP+BwUGdcpHLoJ+wFJ
Cc4qt5uRCxaO3MJNNPtKhYeL052U7ZN0rHQDjQSj27O0tzkju7O8WUerquvVN4Eq
zk14aCr7yMzQpBFHQlEYCC7q8KZ6AsePeuApklhzEBlj0Ez6xJotXGX3HZ/o5XFR
Z5k7Lax3leUt3yA5LY4mzvEkaaUf22sUmj4M9K5EbfBVIT0Vub7HianLLsIDPjZD
48pDa43GUrQsPmKITQV0iKYqmhY9z75lodOV0YRH2lQVJ/uRNh5zyjbo+XKKRuTk
BQTOonmgKnHFTc61zp3RMovsQVKKNEUImEMoR+3PgrPdvRFe1yzDiQ9zoD3ZWIuL
JqeyUfRsm2bb0q5jCgHdn4yjfrIg55dgZYCcFsse97bMf5DAIUzg/2v1I8XhBT8H
HBfFS4cwiKu+XFvw3iEUk/o7tDhCTcTlyCbK21bYNSFILM827CL7C0ZUJECMT6T2
s493NtI+220tJ7VkicMvECvFeyw6sLYZ+O+od5jqnFK+GWyvX8E3kcRplY4ft9WC
TBlOogkm2bjf30tPdG50/UUtaeG5SznWrpkJ6Et8Yphr+phID8dK9uPD6gzIsqNo
e7zhvr95SbubdSk8UR0rwh0shCYyFLfxTOza31En17zlVu+iTlK2mDPxhmklaCLR
b7UJ1RhzQZqjCV+lRHGvZvnXBZSOkxdLmTLxQq5CgZ8yfFr+PU/E9yXuGGUD4udH
p7AOdkMLHfaPeAgjLPQeHR37fuA+MxlyiPQ/+fGcVLei6BlSoOimqsISqbOgYSYs
uNRKDgkmYuuRbyLbvPfae/nm1P5S1wOMDiSXWweHsbkDDbS5gKud4GTNkSuPjp3Y
eAMcah/0spBMIjOttK71xbuh64lvdWA9oNhUiA+bFJRYffPLwTffvH9vzJZhJEKY
1RXBuDprEzJN/Q1IfUUvIH4sELQmOZ79/D7135NqTKo5RF3FowEev4gjplaxSWzn
NgSjAcbOpdZ8e7tgDQmTGuy1t3SoD14GA8vcVfPWENP9g2qMojs0NZIrxNABjJY5
vZuDlHFw676R62gBbYSyIQK2R3BfmWyRxl137XiX1KJymLyeX7LnJxsmDIBCsgg3
KdmSY95513ko6PXBO3kgr1sCHj1Ztd0btdw0Dda0Ztp5Yk3UE5cptKnasaKQU8iB
+PwwQGUVqPgbB9LxDAIqL5s6nZQbSZZeU3VUAkmnL/tsWt6x2NLLaz9b3WnJ2Zs5
OMzk3xsxrVSKroLqh9zWl+hgYakEEx7uenwgRUjbOSlmpPf3ydHJwD7iDFTG/JNk
tst+qkvLDKPqniSGGt0yUA3CXJK9SzdMx0duim7bsYL01relbqUGeDA4FcRHAJs9
QUrI9MYn1zYJATBRg/Dp21H6at/p//ioQgoCEseB+JvQGwYstubexs6voKcEffoX
uOQnY+AJl41+gbts3+sHErga4cjMIRrXTmt1CME5a5sqqwvcRVGe7ldcibFXoQki
vJJonsDQr1Z7Bx3TyIEvZZR4XdB+fRBd7reAUJREBrx9I0RQtJDNRNZnjMtPSC3W
4mzPnFwyyD/0pLngluPmAmY4dPC+p45BooXt4rJLtLRiwV4yELB6MD/DvMGClCoa
ZLorCESwAT6mF+QA1Rvo+l0W2d/SSQmNMI8yJ8/McJuderew+bx7YUnTXvvIeZzg
3PjHA3qhrspXR4jWAE1QONpKXTu63Br0HNk0ZobnGya8EOo//CnU6+BLONgc0Fhf
/ip5l4fYRcN6MFfxNGEcsk4pnlJZb1t5/3yRfo/L56g1VtQtMceSq9Icrfu3h22e
56sH9yrhfYzHVi56PMikYlr8wVCVxuhQl9XpIyLIp1jtXlFCFmacKo6RAwsBsfCh
VIbC9RCQ89vIG/DO2NG4uWf9di6Alr0RQ3vqye61GOSbdp9ONXQYVFBfIb1j+z6e
NT8JitHvNxOi1GDvnBiqFRuj3JuRGFyxwsirq4cURdEGMBeiIHFyexe9/dwFQEx8
iobGzO8Xm/h5i/YpB1NEoEooR5gc7/ZTSqufwoYAvWsttuAbj5erQzPh7l3ynEw5
HhPreM57yxQudIubiCqHeBLAEOTeORY4sZWeZeZa5tEJAgjA2j8VnPu2Y1eXNkeM
g9eZvV1XhBI3Xp7LBfEePuj5RGIxvebOO5xVFNJDkQu5gFx6+o4NyvVxnW8WOM/4
P28JtrBQKIwO02MnJrCGx8PYgCfSA3zuXKezGxOdUaAOBC/wugeMXgsNQ6hYMLbC
QB9bOnpDZj/Tv1SWldrbvcwI58kUvZcL+7nmYd5bdfptcryQERzyoFTvC7KKTviP
ouy2YWEG1E0AWuc4PQFGpNgk3gv5BJh9N9MPrLvVbiPV7R8HDxNRgQgJeAoFDUvg
GEZofM7wNyShAJFANnCWh3jc2ZfMWKHdCLTp5p4UV0+xNO3a6mjeWWBqTyAp/4Ew
JrtYC6bwPhcHThkOy6puYk+bIiqz/OgpTkWqye4eSLmQZyILrFIiVAiPQYiz+cCj
MimQVV+Cc+lSBZdrZtoH9MFEA5NhY6TSmy5hwseP+RBvfl40uOTsk3ibCJ6il+zH
LCET2uYq7oMPIeJBD7/peIzZLAOMZCL8FAvL3KPNdLXAMf+eSZQCoXtrMDl6Utwc
8A9zuTtVVOtKwefWn4Ogn9qkMEPDwoGx9/Gf2NScFA8Q2TotIk+8pS6rO/OQfhGG
31x+RYKeUxzJt0XPkrTqSxpxq83d/LXkvT6bL7qTXYV5T9Z5Q65vDLNN7Wz9Cm1z
b9t67nV0EKV4MMYe0fDBSb0VQ2HpXyQjUVe+5EYVGBw/stGGkSSiNg9BfRadguMe
PcxXOJ+1TM2jyViQZJLij6MPKouzJsYsq42yMpW/Vu5bCEzRi7tuHnhMz9jmMgEF
ElN7WReoaGlbnF5l7JgBM5lAXUZmcu8KnGgbmislRPzIHYGUcPucyBnCXA6yEgRY
44iPmAgySGcAVY5TE0DCIA5ub+tzAomN9BamD/w4kwNtQGzOe4S3OBmJMvER30J4
qRYQbl019AFQVvXHgs6dKUkTU9IRWfSvWCv9N6fC/q/MxMcg6cOTt0nVfflJ9RGn
mKywlCYkBEyOZxDduzPJABY7mCnvjZ/A3y2rOO4mq7FSuOaPffRoC8k73u4gz4O5
M5ZAyL7pYFgs0aBQ7MNVhDNGnLy5G0rnrjFQDeM8TLZTvef/90QKpBUrHI+HrWYB
jjhk0PXZoD+7D0t22qTjp+0Ldo3KZo0wpnOY31HsP1TULSFVrAY7hzmwieZ8VKm2
5G4cB8SufCaISrjzlbkxJKYzlwEaSaChtnrD2MKEc2EceDLYiM8GSOJVLPk09Jpq
RCQyinarUzypMmeOGHS+VTSbExwsuYZyukE7Ami7j//BeW9f8W9Z5uGFLUwi3gso
uo36emfyXW+YTwxerCS59fkmRQG7pYssYPiRWwTH5h/zy47IpFDmhp8OtLUHWbHP
t2/Hby50dCyhlaQP96yED/WtE9rUBz9rn67/eDpB38WNyvqbtl6/LH1c45r9vCgT
BhXUAeuqDY2x8kT4mkrsB2FVITcDX1+gIThtpKySD7YklaViwj/0tNEh5RkzIowU
y/HEa2JxB0oOZqD9gvUUDT4IVUloopEfM/4aaFfUaec2xVNBpSlB8odyMjgzUJS/
EFZmNSPafX4V/+QLQZMBsdkg2555HrS9xa8BQxDFZcq2VDOlYoF07LG4+7z0VBKa
uS1UcBijUAMaDiT3djKrfkjFK09JJoILcPXL1BK0fkdKcjtDA2EJD1/7O5OOyMDq
c2FadCaiXNw0AaJdYZ5hVosabAV28olmNPkQvXYt/6Xrwf2uFOxoobPm9/X16mih
l7QpH3LJmlxyBpgoL7QaQ3u2ABVz/EhA6Z/sjDz/xo+qda7WfWTWD3LmxZoeubXK
FG3GdEB/wt7PBCe6RorLl2k7WRktgmVNRChKqul4vRiN5Q7j7DUu8by8xQMF858V
H1Fde45McM+qzUCh4eOV9likzp9OcNbPR63+JisxFKrh3xarLsxXiOFXzTWVt/Yo
+WDoykJ4CpEYT7s/L4Mlm4Cy6l6qLbLkKXgqG8Lic0f4GtYf49SjuwPITxvM9mjy
/cX4T56z128W6wuUFHrpEPE6GCu3WxUIHHf/V0ExXGRJ5/XJ16NcHr+/LU8Hr86c
rcYqbRtEZFDliZpl0NzPqqeIOE4UllWLQL+1msJc2RTINmpPt0HHzb554Cq5niH3
f/GTECkEek/P4rYk2IML/5WGG/u1FCTIttB67NpBp1tQAq93hPsuacROmM0mcRfM
qIQ+NE3W4HUmIxzKlwSX3a2w3/VhT7MG2BAO5lIrIJxqTse4aaHli7VhG2bMYtUi
7qcMXa4lUUFLbdDPwuMDuf05/QzC9GlqHvPDNEs5ViECBwXc3uia3wuUYIrOJobP
PomNk8+bOOFDYtJxCQMXcRsbHzJP2iFEoQQMQNxkebRD8BFwN3t6/jiZDjNA13+G
GF0gWIF4NwsSMWNNcDPrWf7Erp7DI6JvDIzB0QQlDv9ZDyoqZX5BXRQbCnckhL/3
GIiZaTGU8ABMsQuc9Gak5a+/6OotGd5OH+2LuP3+VuqtlXHXMQAvoX0Qg94kYDxJ
ggzHK6FuEUtgiWweK77gYrmtziW4T86YXtrJAKQ39abK+cSoIEkuOhEYJcgrDxqM
8wlefhDrayVV+tzpfKk44lg2wrYu72zV4zWsNAHdIYVnu/LbbzBnCHqIF23rOdF+
GPRdpOx7zRnuw2TgQFRidlZOlQ0BII7eUGEIK1WMOMgIELiEAmLKGU0hQYgqCDfM
Y+KsTi/2y6Yu97mosMM5DC6/ZdjoN68ORRfHylv10ptrz5D8Mpy/uBhXDekIwE2X
2EhX3QG5lMdl07/3PssKiYq34pr6+AB7s3cdvDPrjPB78uXggM91rSj/UgSXUrEr
Ks1rMCEC70Uvdi9BvUyCjmsusUtv/NB+hgKO/jxN1of93gPyxsdb95O8egPSZV7o
Npf+7J208HNpblPCE1UUBrFlPldQ2Iuc3RVAx7vO4cWPA7m1y6vkDPDKwhHyS8kT
V8hvP6oWpveOoQ61TkCQvRTql4Q7VtYYwi+kAahEtJraFPVs7IJb2bj2O2dbM2yl
wtRWpN921QCAWwuO/puEOCXtPzl8B3LXugryQGXnU3Z3XlPU6KWVTZf1EoHNAhYq
US1kZaK4acRfeBGJ1/eYie3e7XKkbjQPH2b50OXp1S8sAX+MRO97Uc+hlpkOEGwe
XxiZpruNFFmuwOqGH98g+69O0w/cY6ddJvWbQfJNLyRVzNKazcM29fkJiYTulad+
GiFfGlyzqNrgiREwWdcmK1dr8j9hmgkGzE80gtYs+4+toxeU4U8OGibIpRYzEoBG
yI2zhiCvULa7GRa64LxiB0q8JET2fjqUbzwN/G5wXwqA9GqjC4iWPBc8fKKGsHdt
j2nm4Ep/AgYMd5uq+O+PovPT4GHl9DB77hCjcobs2lGq4t9RiayQgzfqYJ/bKHQU
8lnKQxPRhW2YD3Nxkk3vxQcY+LqK558oca24gPaV4MaMuEZXCxpdc/uCphgbSiaM
oanWxl1ihowuEwI1PZbTuDmBdh4pYL5jp1qcvQaKVdqS2gZ5evSXUmqW7hToAZuY
Qk6ipkDVHoQ5OVP4Tas0APAJsDLG2lJcxwYFJdIznJgV7mCtTWqgy1UD33xqDNsv
DgvgH3IDceh98063x7F5VjOXLFBQpnkFhyxQNp6QYcpgsNThgNrJfY71IA4OlIN6
rIMRWakyinL8JHzC4keHxxNWgrlILa6ktZWRx8TFxhL0JIjVFyr7E44uuJ6zUAJO
Jit4CV0qL/DvE4EqyBFCflGuIpuLOrHrn8aYJFg3IA6ndy+UvEniXnK7dG3bH3mh
TL5EC7Kc8uOTqjZk1FYInXdA4Sz6Pf5LaPai+pR08aNcyUYOOTrozfh9ukUXp72i
6SlTDbSCYlCXJb5KDhl90qvTtbsEf+7OSq9dUCsYMDsJOTxpUBu7O503ObROhgEV
E6a5l1lVUEnQoenhFnnA7rKKK3Gwo3nF8eguGfceLGUhPRwdjx9FHdy9kNhnFdYh
Ur2oSf4W/62jDXCYyZzw+wY02/iOKBFcaLNHlzFW5pGN0OLsDg5Jc9fffE485XkN
VFEM8pAPX4ktUMcvxZpsD0CcA+HfdiZDO8BYkVswgistV2DSrg4t/pUJkOUEc+B6
nkgj5E8UZ6tcaaWooloT8xEmj6XNWLgHm2BPbsjiZAX0Qc+pbxCDDkIAVH/8ghnA
Eh7i20KcdqRgAu2RtASGisdad5oLLvE5M2S7kJ/TfV61ncLcbHgzXyHlfjK39Wa0
WewYWr33J1570TQg3g0jO2TZStUNU4po4Q7FzI8VY0Ko0UF5C+4qKmbJpqLT/AsJ
pq8D4emRgHZosA+Lh5n636tjZCZgr03hstgCu2lWbbsWr7wTf3f7atU8+XpfwePb
HjCA8rg6WhO7gJHMNhW+mCWTn7rIdjH15LLnHUSwKxSUzfnO1MlgPPVW9ays6del
z5/fDTL5hieCDPXjfU4pKPLiC25TZ/MsyUpiOYDYJWNgpntganVKJVW+qQnaLwoj
ceOTTxjeytCq0hCLqiyZYoRyL10TckL4e4ZagQa05ck73MWzQE9bC7C8m/zW1JUY
WtOEDjAON3Epi0TWYVNhCwdl0IWOvyvUgKYEtK526fuVmWcAbL/Xjq5MZsrWZ6w9
gAmcUofVRxOhgdEP8hDCDpFrWx2obS2yLAP48BpN1ZeYdveb/rUzzO8P1JK8SFeM
cz9+SCWjnuu/bZR5eZBDo/vJoo69RIEnKVo4a9gjkiQeOlrkaeoY2FDYPUfKBU6T
SXfVhB7ZUJIP0cDKUPSvh/Zi7Hx1e2wDCdAmh5AKocEsmaycgOKdKgEP7a2CmiTy
HwNx/mIj0Vk62ge7s4lH0Xc5Tf/gIwY5mMVR/ro5zyDnw0x08cvyurNJEz425RlF
+9a27ZEFdFPcopP9L/TnDl9dcpMe4kGFZ6TKGtby1AMjWjJWkY/PZGqFofdOuVn+
vBKhcRE04ATstyJzhmZMSynktvnbsNQnnzk8J0tzxxNdIGdh4wMvxtR9b6ccdFiq
rLBwOnJgv3vcEhPvNOpBi5RJ4QYdOrVl5Mb5QRRxQd43T6NQ1PRLuIr0KadOdquT
YGAhS0Uq3HXLRBx5dG0JN7DVrjiz+Bl97z9jI6X43qY55tZRySFjiljFXR/KzvTv
CS9hu880Zs0MXQCdt6gH17OHKGIQCam3AYi2JtHqZnOwCx3ylZYMrsZhYWfj7lO2
IOar0A1mBcPTNjoMSFpQ8MT8qERPNjFdupQxiAOnKY+3Zcx4WIPVaWPdmZXdk5Wd
EKtwpjwXis5rpP9IEVlOzfmzDtxpt2W6oMxxF27AaSTa12O90toFUOncIBiScUb2
APk/BUv1zAPJmiUOTIaMgxdRaeFpAmu+8djS487w3ujovr0pcP+qsJmYqkwUupTI
CQ+mQwoF4YfOJ2y4AqZoVB3/LRg8zVqza5IZzLdl7eOLLJruB4HOWLPRn5KLIELB
w2fLQGMeZBHyS6OTFWvU/vluz4lQfCCSkdgSubFFqd9aiD7294V6ERoQx4PDvCpW
ozdKg855FgKupoee5mRDR5CxEPCGdgF8xaU5G6i0JE0EnWD/5KMNhEAIBnLqT5GE
UEXIoc6F6IcHwvg6loqZi7IofOGkSSjDCKeaX/P0Z+XBxK2QYmkd53Fuep44BX1O
ypmBFmLZeihdsJXlvIMAbYg17mfk2SP8CuYtqDlzD2hpfjk8v7QNaVZWCYZa+6Mt
ng8qnOtcHBrOM+HD28o6l2cg3wEF4M06PeaY8gorrBeXN1WE/8t8UWbC/GEqldE/
4AZkFm7zzKumyosktZST7uKRt3/32J+PwNxeAlJ/hfetX5CKwrpIZAQIh3AadAQ8
+nGXTKBVwaJ4XOt7jJVQJIiXBiC7+/XbHtMs691irw7WFV3G9JPSPpUOCPYgsuCh
UMQD7QRRMeX6GrECYK5huemo8/wcsqqF4XoWEpNeJvL1hNw8aI68IxFzcLcByDGL
YJ1c9yxR4gbm+5BNa4VdZlx935Z3HI7EXSNnUWUEFB5/HsXHARU1m9R+UBx63B0G
TH4UnpTSOagPApX2vyZdzpsWMjhK5DWO6va5ZkcSXVkH89t/F99PvUorHPqGBLku
AC7olsmb4Raym1yme3Bt5MsYqCjfKZ3NuOKiDxvt81gjFI+79A5AfkY1pcb7wjnB
ASZNw2yB72P0ZuJMo98pF9hYYs9hu/fQuaw0TWzonqXKxDsXo3Q6CY+VGPeLx6e/
iZGmL4UbKGRxJfCsGUSf58DgIC2ME/uzN6g55ZE3DDfYyAr3THC+lyUy1tCIq17k
xQCmgDdyf7LvsG7te+1ZsogCYJvrsIel2OC6mqkF3KF6VhYQ4Olendyppy5096ed
dw6s2VV0kOs6qIb2yLffHsUCNq8QXF7iAZAv3aVbnqVrBoznwq+7e96QPXrjpSp2
ZUohrU7l50okz31AT2T2vc4MVRzK1LOaylBNgk7f1zZYCJLygJCqUBvU35XE2VhP
EDSflGWsTtrxIbjz+V2LUFoyulPNxKDmfH68MdAoB3BFVPxiOlHiv3PcbatXEgEY
K4Xlbu8jh4eBTW9+K7fg68g96GksLzeSw4J6iVskhglTjz2IEgi+SoLxNBAFQMmS
UsJQGWSu8wa3e+uYio4o7DmJwFARsnQWbf6htEiysUna/9mIxcH3VR3ALiO4g0dx
VoCV9o3bLiM7HQEy0o/LdAfLmv0OwWGFQUaPyCdOevKZefGTNdUA0eOkaEKAgVdL
y2UQFqSxgq4NubasioWsJoaYqNtkHo1f1bQngYOwvpqUqW13sxzmiqqJXAITLB9G
eLNsYUKZkqWgTjYbBwj3gXkvYhW2kv+1+/6MyZHiINN2nz0eW2pjZd9ZK21A8U2c
88eUS8bnvMHE6U9yRJUEoQUHz4o87oyXb8psywawSSwXrMOPtMEKkcgwcK/8KREh
fMBxfGbZCi7Ad2tJchb21hge4/OQsA3Butt8TGJP3AI44PVxN+Y9ZyYy/MrlaAeK
3Dd/ih263sokjqWv2yo2sglHnPlxXFNpvrKzXs0k/Vs3qWNtB2FY4TpEZc0ZsxmV
LK5+K6uJdFJ+cpAI3TSms3VKk9nBvEwO6Z0mCQ3Sfhlvf1Mm9DG2tQt+iYEWs4od
b9SoV7tgucI3wxKt9CUxmdqjIkcmvPmg29UvFodHWzYvCbIm04vkcVaDWelsz+SV
fYguG8HQfGDkwMpZTb25tko4lFtVOrRr0qpEDqFbKQqFgOcmJkXz42ZQq5kQWA3D
b0arCOm0fZ4dwfzXp6oy1iymRxDTCvR8qrdNj/VP/avwhLZZoMUyIqVdv4VyzvQ5
mxEn9pvN0awTHXAWLmDaBZUOyJND5Zo2Q6eGLTYPfWNl8F3hHirukwyMfFzHs9FP
NXLe3iog+90wq4OrDUSe8gmGaSa2cTPgAwb5fLUGHDwTDCwqIsCYzjYtVm8fMz9B
2KGVeAD0GWr8Mrvg7UCDFk9d7DjzpwC6VxUBQXIlivPdskloe0dRbStgDPaF5jaD
PxmPZXEw1HJnUhuXJBZmfGpSYN1JlMIONFB27FdMX9nBelggLkTR5vd4nmZcZZsv
ZxXbzROyI0A1mYCmOP/wDoeqPWgPvI80JwpRxIlx7VIGfBZU5rD/jL9BvnzN3fKt
MNflwdg09aQUIi9BN+uIyfp49xJH+sY9VA2CJAtrdAPP6N2hLAMno95sfjC7ypN2
Ahl8YcP8EbK5E5JqxirLjLxrFW0u3BZ5+xeEoyudW7XKi8nuvent/wdoWL0t0ohl
llPfj1rbGpw5Nm1H21JLxWBoVwIoCu22B+o1T7dp0Q4nMDas0DZA69Y46Xqde1XL
tRT8MHKQHDHt6Bj/Z/vvkmR3YjWkuSpMOXeiNuta90JcMOCNbmixnqMOtBkfSEG6
qAyagipQCX9DuATayCe+Y8Fc/ZVWY0RAucEZ5T7NoAoHKIH/k5Hw/3IPKzm+2VCs
/YMPX+TSvSnhLhMvbgzZhMBnbUGm6X/S6xFiIJZpqcqPI3tHlR64VmKZGXJesUDe
z58FXEy3IU+0w+meijlGyzxe9E5/VmZ0gOyyoydxh+Yyxd7ghFWRX4elPSw3ccKF
zLaUraP7wInQga2iS3aPo9uEmIpRrS8ljvpVlqxNrJma7kc47RtfsBlPmYy6SnlA
rN1hphC6CHVL5clfhJ/zS360ftXgglt6rKiM4rlSjpo+rq5VSwXGCryIhptQic+L
mWD7as5EkaJI6bVNJLql8CyuNtMm18mNi8xNrcNKjO/JJ1LMe+z3IknTOciFJC/R
GYHSFqpADk6Y7fz7tqELpUR+dCpb9q+JOe8jPr1ZiMq7xXhV6sFzPBeNhxXYglGY
4nIKXh7odCD8XwwzIlEqfQ3hiJntnk0ix/sXzFBHZANbyb2fqS9NjkCTs6N+dW5d
FrzEIXd0zi9ZCwqEn8uEMUeuo4pcTtMBaNk8cwPHI5pPLpcTOyJtninFad/0HKwc
nKKxHG9p/SF2ZcE/j8j17xCOfwcA82eNUJs7TzfvGeLH7PSRbrvKU2pEzDKuxOIm
rXZhh5QDJkN0OKRTT8RSGNuY51P6o9YFEWiE0I7lhE/C2IqFQJd4FllQopSjej+a
z+rOPjqjjA5V0L6WHeTWS0QJ1rM2jTDB62fADnRdl+nSUevWtUZwobkXdI1ZpJRy
A4XxabmJLY/7JJ1/QTsGAUJG2bVquouxhB8VLM98KqwlN4zzP6Np9Uuy9H0sgTqu
aGHJlPFnuj12jzkQV97xqRpu4ekhC7NWGu6nK6s4Ta/02ijyuN/gPuTSbzG2sZSf
+S/Z6SYWRCLozFzSHEot+EncqKSh371CLyR+QEYbrH9tPc3WFv5n8hPBjxQUUB4j
ibKsgndAErA1SlitWcXOabDFEFAs/QHweh9ZEV797N8+w+vDFvo+o06/tvF/xsX2
T73KRaA9ktlsNp++21uYIREGWoCKot+KiMSa7mIvc1xZhqpKQjMpCq6kt4qlehlX
5rJbjkGH6e46ztvrPxOTR+RwPeDWUrC2Gv5CJjmSEqydxaC3eksEI1jkIm9aRjsc
MpQhvY9niIuH0HR/jUoG0+p3Hs0tXy7zq5BdDpFVEoncCaFQxvMnKsQiPWeHo4TU
WwBTZ9uFEZuR1pZc9STJToWs+74eXFm1ijYeVt42DBH2qvCdCDBJ42PAU+ujrdA+
BYAD6A1rpmUTM8nLK8H6cvzCgYMqNNksrLismXvfZlCYwZPDMmdc+PLNrrfiTt9q
VhdHt7JU9PU7h1qywN4j7dCyTjuBicOoffmZqxA7jHp/cXk18KvAQG4ZCHJcgaZO
rB5VSiMQXUlq+60HMSGvnkdS6oAOw/BPhnK1lVv8QPOn4ME6GN/zPa3/oGo+pzu7
TNEPDOnaz70RMkLm/gfy4V+jygcr4rKzroRtyPhDamJgDvJRqQQJymtvLSbgZuxp
6K9ttcXAmaUMomTRPqvgbTeFOBkZAMX1PzzZQ9Y3J9bjKMXOK/KJCoAv7zSZzTt0
P0wwF307reTdkZaE9xEL5pzGGZgv0gEZ0xSn5zVrx9kHGOk1vxec/yOg23SAqNK6
tRGBjC1dhPcwaa567drMj2W9zhNdm6HQscO8FCf224ZlCt8nspdCNTbtLMq3sDnG
3dAxEF/l9fDEs58bZ+rKsQMkvFrWvqhvnCUxdXxSjJava2NqkjNnk10jfk5KQ6O3
5apQm1BYn2lnvNjamt0ahtgwQMvz517El8XIhWf8jesDyIJs352632gJoe0dgNG4
qP2mUC0L2YHwlLLa37ckY3v4Nf7ws1ySasKvzoHQNP1EQmjK7LVJBWa8qSNSmRce
3+pHC8YtmfGl3jgA/gaZYnQlbnWKbiMKKGC8EbV4Pq8S86R3m8d0rJqjuWmparTs
QusdUYi7OHrPQrhjcu8JJ7OgMc+Wnql7zyml/kUEiqzzd69D0C3DD2coKDrN1Ble
jrcYVa9SE2rIRfU25zlXWtYbky6w9eG8jhAJgBH/b0iCFon96j37W8iNctMVcLl0
hUwuegG+v6cMs2bl8iaSzC5ReM1LUrzCOR5KrrcgbAj8A6lLywVXMwZjDcE+1Rsu
uYj20KgKn5Snfq37VRFNn946uJRvVsuP0EaB7igV1TpD0xdD5JhhjDPe/ATeW48W
dT8HwOWlc+DVr/ViFvLX0+SDx3/QNeTtW8T0UTEi1lM0YMYJ5EQDjF00hfQbWrCa
K6ysxLQTUagRbKuIv9wPuNFCsAOlsNOUYbQBr64eln9aAvpbgmpFoDrjRX/W90KI
+OUGQbSmxHRH31LY5McojUgvT6scu/P0LrzeeftZ0NU20u+oH25DHTBSQmq03l/C
qnL6cKhP58CPsDyQi8vxnpDfN7rMoNr9qc4dfe0SIL13FvKpFXkaZ/Qa+4qDPjk0
f7S4OSlQcx9VAhaSsrUBsckhz4YKGjZ/lzKlo6cTWTT0a9/Nu1kWZwzHHcDE7+cA
otKI6JNYPQ2uU7oPvxwcBrGq50DYNkRbCq+M6iPyv+Dxn3UoLTu9uikNpmZJvk6i
itZGJGNLClqkWQV5FDuaySmf4yK+XUPNNlDA9nVnI/ZIhCT9g3CvuYLQADk9WMA5
rt1lrNuaRf8P2KjsPGdWmh9V9T419hzm1oF4DOrxCW1vyHp8gyhsFYXmRbT7xtv9
BTMfCgqnMEwSyyUUfOB1MbLJn0Xbv2JfStoH7qaCMDiUN3xhXKgOanPIfeLwwcnA
avQ6exKA+KMhR+Iu/m+P9pMqIZGDc09HXesEcGGf6TPId7jb68yBvCAiUOG/Ll+v
lESubcC5Ps+V0drw8vMvS/VUSZ9G4rIm7S9sWqckbdl4NoN9w/REI9EsM5ck3GcM
ZdUwsR4cj0Un3TK0HzLigtN7GghonNDCvVo1o59eTc5xJ/1YlmHGc8uuNba/mPbt
6dMfS6dQ6lIIP1vQz5ESyG0wU0nF1jA85Y0SRXFEtPfZNzj5rryTAM0cXNNdOIif
an0PGZiUdCoxAWdgPicQ3J22Ty2xIadJKgEkYFrqGEXkSKIfhx13uGaZ8gDljO3Q
ornnNHgXg55N487KRk/0UFXTFbJEhb7fZQuH/d9e5osKv3UPy3dsmTeYlJS1qrep
7WJNe6M/gZGMUSVBCE4ESA4GYomxmlJYVb0tDwomYhDWAQv5vKmicGIvH7tKYYKl
oNenHZJItcIHwu5T9YJG6zxpkkQw2Fgon57c6Tg7hl7WZbbje5PFfSmZRHJzb3dF
Wku1+ZlpPg++olmsZ42QS/YGZSsdwnlZA/Q9E7BT4GHlrzxoCWBUcmDmmP9eXrTU
7KuoSBq6xUJ2RRXqbeAYJ6Rfsf+cgJ9MgQv6YvBlEd+k2ysLRe60VUSZPGe90pX8
MA5jJd3JQyg1DUIMJUTpj+ZYTzekL1G1AKB2M3nAGpcvhUqkemcaW90g6rb967MS
X0qkdDYeGjEwXFSrgUw8JmkIamuXVh5pkv4C2XJcNL+JhG2B5xTgBYSZ++r2bXI1
ButJRBU5pbjonvMdMH63CHXHNyNesjuxeC9xAt4KfoG/nCjJOyV6Hj1lD4PXy6kH
BSSoC28fOfBF8o3vw5I9WsACJ8dkL31AKEDVCiZ67HcjVd7lu5pp2pMs2+N9kmOD
En7Ekj4m4Lv1aptITXA4I7hlsFTqfqi+cj/cuJYPq9jnadWkUYEepLL3JYO3nE6k
Nc3Eo634t3grPQB7uBx8j5CgITYTezZn7Za/9U8spft7THgEz8SlehgsZhh48Bq/
Teke4mtMtdm3pe7ibzrwO3D9LDRJMYbSiU8FPY6LQdOqkTPYf0yoVs7YRcYM4ZqG
cPEA9lB5cuyfY74iCD4go1yg4F+0VMk9hXogkbwRmOExw3qDDhVL7xRAkIaHOybF
o1Brf2SiVD8pAYF54L/hSdGbnSsmlxYU0ME/+/pjeHqY9l3DGmdTTJP63G2UPxMD
HfRBclFyQK/aw6Q2A4X6xhy4oSBkrxdgQbUTCJbnmcA90qkMbCzyWkpW0ltk0M4v
1j9yX+Alr8Ouh/dI452uyYyJnNXR7XAKRHrIrKqlBd8qTJ1JZeGZGejpIKhY21Uv
2zudiB5F3vLmSXuY1JmAW/r2fzC/pl0W2g0086jkH/6C4RDD+JKHCgO0znauiB2L
66J1TYo4SqBFr0U896qp07ISZSHGD5GTgFO3v21X6SBiCdalFRbGK1hHvsLGxtHp
A6Je3lDM7zzO9361MclYgs/MFhOsbCvLUsz/tKghUje9dnv4/U49qoNc2u6xJHTH
HxIBqYKfjjFhbJ0A7qyzAftMVPpIZhGtNr8b1/Cy2vHOa2mGL+/4Z7uUXY2ZA+8c
vTLuFLh4p+b1i38gnvBpFq7QTyPI1B8Je5aX7PJIgwS0ovNE9v5o25CE02V5v0ax
/gL93mwEpayWQaDHyubXt5XD+MQcoXCjfMsFLS/U45hwtaxu0F1Tz1dY6BBRMp8d
A0ifk6XGr9lCaM4QTha3Wda2OKbaMN5hSez2iLaKft2tILaM9ifHNm75eVrPLazV
6C9V3oSWKQ3qabWqxYAMw+tiNzxLIQuWRdQxnt/TRq7jpaHR/Uxm1v0BSF7daY9F
mbz3WRjMcedcUlIGZ8vM0SO9O3ynof82APNn6b+jIz66imxWGMFK1J9FY0iOBg0e
FYod0OZY+a1dm4Lexd4KgzIYZlVNFe8vp5CcNexyo6vQStjSzmVCtNPHMXlrGXk+
tGHR6wsPQmYP5rENRcTaUms9rRwLIa3HHBs78+4orgS5tvsY6CN4voVDqcGhj2Zx
Ps4Da6OrWozyWN5swTv9zREJUCNJtTXfxhH20pr5zEoaZQeWxFe4WraFsva81vls
RMSiqXIi7l3rAL+p0kV08i66jHR4flRtEQrnJLlgrwyL1HXzry8PO6QnmNArHBzM
zwEv1sNWaOX3zqqK/zcW5cfS3XDhxj1bn0HmcZayo2G2yNcmodNUzHisDvUXlPdl
gFugY844rw6VdcJd9oGQ77kVQGhr9ohJsbelHjQlTRMhQ4E3UleDL25kZ2HOap+W
QFzDLRDBdLXzpNeTRu+SGXJJXFZl99SMHcyUWoM1NzPX5ihmcwIyB2rGIRa2k9QI
IjFJuoZd4TBGykhZ2lEYqpMlKd2s4K8+uh0wCUySBDxLLVQuppzVEJ73RWOn3PB7
3yJmf2cc36PzCJ838Zi2W36/0wh6V8Ca0yLv8Qv6ozT0Z8cE6yE0tqg2SC4pkFSz
tuLrCFs9e9Ihq8hEAM6xqKUcrfwB2L5IZMPu3FC1t+3gWHNwcGADae/Iz687si+4
QGKTR1xNV9SH+giufmUU++iDtTwuhK2B+DX2rQ/2/sAmt+JfBsfyNnY8wlT37C7H
T6YlVubB30DNMiW0Y8MqHwdl9rFGlGTkJZGfK0dpysLyjueENQfa33yEljc475MK
tj9icZ+ackF3uOdnB3s6aOH2/47xj+hobrA4xVOZXZGumDF/wfMiCh//DBK8uX1Y
UJ8Fl43WjasqTree+QHSmBDDqj6NsLEqLUcDC2ha7uqwBWQPSHj+IAXF/DWGLMg0
9AuPpWviMRBY1nbyeBSLgrb3SJmaTeVS4szLonvydHZvTq0c0eyYXXei7Fx8reTx
w5Pz2hBoyUUthcVFLt4LXz+0A22JUI6U4frkAewsDyJcK29y+1ysAbXWPYg5rvYY
Uf3gqDsmbdQ1wvT4rFEABsIdA36yH2VGubVWOLstCU12xced3Pedv59+4C1DuxKd
5SNyG6fkEcuJls33Fue4o+SVoac7uEKd/esU0HuL/DamSiwpy1G4A/nkxDnemMNa
tAvnf+asdsAQ2IFwqNsqlv+Rn578vaN8O5R0BJapnGhGhNEOUWlIXzfRUmrm8hgY
dXYmVS8e4To0DbNDpjhwm/5jXiT76qFSPv/1YgAFAB1elWZL+nXOfapd45Cktal/
Ow6FFRB5NAaO29ZnJAInwazF9rLaqgu+i4cY4CFwdeYpgzKpBsvtSFbv1DKu7AjY
yp7DE+0d+YhnFick+Sez3Np5j2mfV1OtDU9As4SSpxqWFK/2FgmokyLj+JmCW2ql
yZ7cCT8O/YN6pQaR4e/DqoianX3pqGFjeuDCiKq5ImFbKGFM7yTdexKV06uQJ4jy
LKpDcSFhJXGe9O3nl88JVSeHQNA3jfwec/Qss/BIjJ8B5xwkikB591oAfmmHR75d
80pohtq33PRCVwcu4D+Vk3n/7RiO+0p4Z9saUhVDoerCbI+09SMKsYIIoIcAatWZ
AMAoEup+Q0KhUuZHuVxxXt3c56AI42Z12ReNj3LQrocGAR+rR+mhYTLMpUmhajet
MGNyklEYeOoPwepxw2ozHRwRHp8CNlXRv+WaZkG3eqIgfdq3bD8hayfpio9bcZEn
jI6FV3ZOWZ94LHNzezfCT8/C+J7GwC8hKrkGwrXVUTApw0cVuyjxSNvBoyC35Xbo
dH81lWhru0WdFKxM5vQkU4a31gfWWhebFlmf+5qfY5igE5KzMw/DAgdX1UBDzlBU
1NwLrxfzO9MupxBSS3+agxl16+lEeYrJ4kDoRhHoXinybVBKKMBv2CEF/VeCtckj
VTKyjrY+xvQkMtglQaJvERqHWS/lr0LPkR5OvEN55xsAxlEtkZlH75yBdlKWLTUw
pE8CnIWCg+KZENf21jGH6fAPTNaLHLinuZ9leHR8mwNYuW0+puggDQ6/mPeRWhXF
qpC+r/rn2mn+vptmBQ7UC5eX+6SJNE2/ui57tTgeXTyBlociVe/szXX0l1Kvs8ys
TNLoiY3gNiG9iwvPjvB+z6yJx+oBnfS0/W/v2BncRH+Mm47NvWV2hadlT+EErwqQ
w93TmaB7RrYqkecIinwgE4CDk8yvvv+XuEwWKrt9gWMTrrBYL6a0VHPe4hsafsYI
q+KOXQRgKjJtoE/o9xwHeUudyvWDjJLZorrQ3HhW9qYDbTYjhhnkCfBK31X+9VsO
GTz9sJ8LICoV1Vj65bY63/c0FE6BqYR0JUCU6ryAJy2WjEJB6U4lFELp+vu9Mk2k
H+UMrqQbNKw19dasXO1Ia2+ID9L3yTdxVGJZhULLh/xuhrFktwKZPclojItwllZe
zXWZ865ecPTDjjYHb9pZFADZGQQDYEOgXfdvqasxl4sf40fJFLfCLfpeYZoQ0qM3
6XAX7GtImsv72bfa1zAFzoqwRfWw3MBMHOJD4O8CDPSjjw+45WqvpFuwJT7WyJ7Y
GykIvW0sjcqpmsasfe/2ukc1bfAFRXE20X+nZfdCx9xARl3Z9Jgs89sQaffEUrD5
2kq7f1/phJtXIdlDQD9+7JfIdIlUAIInWk0C3yexyEnN6Srhb2KnE6HbbLTs5YMP
/8AHL2mLa5ej6Qoc/oieoyP3RgzqNybdZdtfdh/X0/vuiRhHaFVnpfe6LpF7NMSR
4kuQr3JeP4FHVT4LLZcp6ZCFb7N8ftQXiFVKztIFKnDVJV0idwZIIf3NnQk/3Ga6
Lw57GsIQ8kwDWwKI3oWIZKcMO8jhpNbgz0BnzvNGxyrTPAt/Ma17t2RyaDG2cLLd
TTEFRcO6zO1xrHFK7JMuA6E1/rcG7/oi7R6FEoM9bs5cxCABar4b7XEUjdLjJQ++
DyHa6jsyhvydjbrUoSem8MvxOPqXboknOJQcCnDXTt5KIrxPo2oOu8RSbJrgcoG4
YsHkoEzdLLQAqOs8DMDh3WNaoPlqZzA5eytKmJNv4rlVCWXsGe9BS5vHYuvGGJZL
0Ex6LNtr0w1LBDRri4wa/nQbO7TbeelguWNDGuLVvGkbUnH+QGNERyvAN9fwzCwV
0a+Fmhn+qPgmU52U1yjKp7xHUNro80fX+Zre1Vpn+JP3AfhbBYJZzS386MkjH9Fi
VXL81MlthLLINvq29KBTPUnBqm/r4ORz0s0Ka01FRI18BOPf/5Tpjc/dVXk5O8US
EyvaPu00t8s2+g39BqX+13AdNe1hOvTtZyyXm6+ifn2rXUwvhkuCjaT+zxqUd5OE
OUblPL2T+aIXJ2tpjqCnJtjFQuUzWsSN/o5xwVB9a3NLduEj2HhArFqZBejgw/QI
YoZSe9Jyz++ykV+G5Y+x5m4VfSGmuz2N2PRWj4tY8bgxBQ8XP37FujX02VeWgHpJ
a9uQ0RZ2Y+1VbjUK8S7WyfaFH2yBS10Ij8v7ZSFYGcIJ5an4JnrVzS3GHQIjp9AR
6xsT6Xy3j8Um06LeEV4VB1e5WqEIGFizvibrjUsd1AWBIc/sR7nvCufEQbgdFZih
ux1gDxtYMVM3QnQidBrTWmwTOrbONGS3VzDN5+4crPRFDOJEWeAdwQtG5Tg51ciQ
LDfFwB7ccw2T0vW5627dTx5GMye6KkpYK82kmpwoT9sQ51VIP4uJk/OLuDX8aoEP
/s/i5DOGNP/6xHwEJNbZcCQOfp3PzKi5VxUxfnFdBt6+wKbOtFMU/56jXi8U2+MT
uPeOiMWM8NMG3xaXbTKX8mvEXfGwXtKZAa+KdygeVF05AnsIY/X7X8WmomFGcfrd
CcJ8AyFA+WokhqL9sYboo1+cxN1To4pmulc6gJ5vio0mqvxbaXdS06JhlzxxkbYq
sN13U24PX2cK9M9AC2YFksP57DJYD5tlr2GyjNWRSBOfZPX9LLW3Hbf/liq4Yy1O
6XfCDXjRMZLTeML2c7ZfZ2bxPqQNh2m1wvPUzoPwbky2m3ujUCz+rsDo7w4UWtez
s1MPPGi0X/GaCbbPRpVDQ8R/zxaX4VjBy5tBWwsTLh/IgIro1OER9I95Vm+l0I6T
X3k4tvj4lTcT6D+oSVr+ZfMUKbO6OgV9ISdSRSceIL36KD10GeNW9vTeyFzB9skQ
VCuLREZnSZ63rDRiQYyJyHEEkfqqtYAdFLDaplGsnp1Lk4VdN3hham6WyXxR70Xa
CW1efMNwNGzEpONeZUp77VKi0k+1rjalsdjLplWgMqyTY7eZ+9YfFFcTh7PDaUYf
X9eUPujvpD6jp+gOyGR6Z80dwIPfdt9uq0kFtwgL6nVJQrkN/2OFn2YM4MDpOjH2
KYKNsNp63nBVaa0IU8r0/WS9prEgj3b+mGQnu2d/kGMDGNg0dOw0zmCIwul0wA0s
fqWT7FpxNY1/NdYCU9EgkR9t95PqxLa3NS3CsI+l+L/dflKhhhL+IOD2GcAK+RlT
1zHeCC70xTjmGjGW5TcNHMu6gEDz4cFlSjjowEIMU6IH7Njt2bQyeeKAMx/FXbaU
5CElOiEgwddmkhoZuOPrhN2uZ46FJeGhZOo1yI59yED+va/rYyrB5yl/MwRQj29H
7QzWAlavYodHmLIg40UjkjBSNPpcYlp6bqjlOp2NC7c2AQvuijzRQv6X5aeUPunK
WjK2Z7Q/DCCs1Ol0pyrVXYRUg+SuXbLtpRHfH22Nw3vVNJDqZfIG6B9tOYfKk4JT
thHCcv3psjb6I63cuuaFGlGERok9qsI3sHb5I1yK0PwLTRXUoX96vi5T9uQWXzx0
JUT3nqbZb4cegdBrNfaanozTEheIKXo0V/HBhsDd6HAMjvAlFiPK6+XhczsbuwLr
Xblvj5WsEDO+R9ldMQ9Avd7jL347NOjYt6ZXWNNiR2AZtEMzagSGBcFEHZjKNrpC
ui0Yyfcah7VnR5IbkWMqLybfrC2SYBgT7yz3ob2JPG7sO3JlkA1P10xPhX+f0lrJ
/VoUj0o/yPX+qWWmbJLt5UZSGUs3prqlRD018IgF0F4jLwZxiIay9Nn3K+wZ6Jac
0gfkOavc0S4G4T2C4f02CkIKT9JWzMhNU+gzbDeExuxNDQqPeUoduqHQpEEXx0WQ
9qxf21aUHJJpjE1qY4k9W7dBitlgt6wrznO7A/sYsIzI3lShyAKZfcsAEZyanSHf
B/pIiQTcSf3h8gpuvvmHFHpXsgd/bU3tG2Bq5895M0ppO3KfBQ3nvJ3l5hsGD+Ir
u3JjRte6Pcb//4ZgBp6HwGid4LMxRknGU1ZW7UPRTIgvB3QAGfGHmGJMZko3gyu+
fl1nC2YuqI4SCc+PCVkjNUX5Psqgl6YvUnrWjST657e39aslDCGHdazqk0ac53jG
/iHp0P30dHEm1ENzptggwFiDtHFu2QrGlDYCGgVe/zXC410BdXjyjbByD3MN4i1k
uABQeFdJXVZtkFCt3gpGH3K9nRLevEdcnp8BoAvxQeLey/J/L0Sa7np8DoRw3SE9
9DT5Kr+QurX/GI6TcxQYhB5qOalQAW9n1uEQ+doFdDHNeXQ+TgJZx0RUmxl1dR8t
6Kfdq2piVIkBzoEMlxVHzhc3x7Zu8Q8w2GHHTgtwbpbJMCDzIuZOLz5pT58D/R3u
ZWBkZWkWwucsOlSi0/z8JcSKKpXtLUw1E/3BT31zf6P2bJqrpx+Zi+aDENWwpcxb
H/JMcSqR1xdFrww9R3Fs4XGukPxnk0aADNxDX/U8yWiWfLtGaNkvOLzH8PnhyI6H
MEkdCaZmcpDVdLJVTFyWX8jMEhlUNFl8IA2PQLmtfBOk8kxC6EKisXkeKxzbad3D
ZLtHZTHGWv+LRp+5gnJ+Gb4g1LqA5zIla9Ke7nCz+ImwPnNMGz7SJb2AjmOJIFvv
H4hyX70OxPQ/2dVR8ZZxBqOwN0f2Wr9AVGRdQqJJsFcirE+wfH1ORc4e4llHUkUb
AHjcmcDjqAK044+NE7F0tMQOZHrkxhZdztedpNHgRQIhLtpsqJ9N1WK4ZCFFkE+N
0xR/nc4FwRKjOq/t9ly2ggRfYWct7L14zIAU7jKJj+m+iYWQ8hRdLrK2+DOshlKi
iPYBo2ksgI2xu2HM2GuuFzhE/ho7sQ7ZrZdZ9w0VuThg3CqfwTSyk/KIWy+PYEll
rW4uoxmtqPtMOB6q1F44RizWrAKdYmXNoDNFiWymheBVXGSSveYBzt0ZMCm3L1Vl
7qKYX0bmJWnvv0L+n/RmV35aN6v+foj12jTq0kLgw0EdroS0WhlF/TE/EVRK4+CC
W3nOFM/LQWaThiK7aSsLYzxVMVYpUxQI4IF2rGA/fGGRyT8SowerxcfZTiNjpGjw
QgUdV+w+fS5sXSsDG1p+b8iMEU8hiaEGKQX9RhyeENyRWnAeEI2yyeLUAAhZbi2K
7TwqrCCocOQnF4EOn5kfI3SBwcV57eMV51YzIch5NmPzTxbapGL9gim51QHp3Gu8
HrvPWzWtlQkYxNsX9Kw1/AiZXoSh3YOF9LBLo1tgOq3l0isvzzFu8KwNV4uqIWPS
38RLUXgpgB6mahlAXcOLZmPB8uL8Jm2bxxyK+ftjuj1WQGfkPsphCsiTx/ibEmGR
HB4/rCHiVg4tIkh50+gTBVbiLreXcqlpRZ6MOEn8g6fGt0OXpyawaNhg+c7eofFb
x9DezgcJSKlOotFae/oKZfdoMynilhbFW7nzXf64Ccilpk9JdwrVzBTXD/xIe6lm
j1Qm298f94a92pcb8l3Z4rNj2gxUQZIKRtBT3QjEW401HbFq3+jPwmea/tNP00d0
eves1RzAVEy8gA/JJEF46aoNr/AuJHzSp5o+/X2gMvNvN+eEOY0B4tkFz10a1UQr
tWWgpF2zTibfwbw6PpXWjKR+ZV9c1qIoyAfHJHbWZf30zZtSfnHzONrpXKB6LIj1
hlPQqupuStwkwzTgFAB7hny4hv2bRV4NHuUENuHCRiT/HakRkJUGZGUOWKUesRj9
agdYbgWcCdHzwhlMp38FpGvAJFNfUkcFoRmlGR76+X7I7bazC6jE9WxmF0DL/M03
l9mYbzp16asjwFjmwKyHMfRzES+9feraI+N3XePohFOiPaPE9DIJquZXTB05vNQj
EBSSAkYFSwP2RKxA76RMKBcfMsygenmfg3sCXvV55yMZV2l6fR6kj83MnsRP2TuX
WkgVQP06Vuwkg4rqrpBVSI22gc0ShmgsgM3KCd/j/dueS1ua6ZVrrnYUvj/uKH71
RUMcUpzF8HwsuUkLHCsJYU5DPkD0mXa1IVAuQTalDJ7BGHlTE8xKwjl80xOJrJgV
MljVVjLK6BfJ8dFv9KEZifgopzF5TyEJUxi+/7L594bhMVPOta4hWT9cTBbI4lOW
ROkUpotnHQzkCS/DTi8XPv1nQeggsukzvwb+4+FFobVnr/1jy2MrNYCIxjunQCOh
pxdUMqS3egpyppa7C7Td4/IAwQZFuS+aZFT7l0XgEyWB4D1fKx6ZVU+zjckxS8zl
rhRObHOi+5PuiFrueUStTUYul4rFkn6orp8qlUtZ8qjH6yYy+It+uuIWP2KmMY1i
SOYDHkE5jvArFPUjSSEBT68xls9OMmUYqPSvTKcg89MlfovMTVM8DVxzZ55MUqHh
7mibABVTo/tcsY4YflBSseLNjnoDhjm7TGHkyeZb9/wyqWf1VS8j9e4HZQ7+MAoA
XcEKkGb5CuGG8OO0hg11ioTROGSpPRZwx97JsM0wVugntxPBbFtVNdILV+vWx/P7
3+XlsY4cfeYu9tG2t424WX6sk5jAp8Cf9itleQGOUYSSE7rZw6oKyEdgiaY+DUtW
LOOK9MWP6tD+Bc24GeSpOvhWuYX11TgxW3sQ02bCsJxyHP6j/7D7Eep3lety/OhG
rF6688UnNLMH0BQRclBHAI4UOGCxKwgOtXi69lYOH9HsROCNKcxehywAU0R6qbG1
E4rI1Iw0DaYxysVxWyvh6EgJGAaCZgL7IJqQqLzBRTG8R4gl5V7rM/1gbt/ntzTd
mJ0zFmXI3xMwZUWzBNJqb3Ypnrt9b/i5LuvpPTDPzru/q63oPvqOW8hEtV+VE1T/
k+hVwdt1B8n3d9lBwVlwXEx4RfcLtXUhB3didOFLaaIWKGT+9zSYGzXlKJryFz/f
CiTGxoidbSmZr/E5Gbl3IWQu/G7G0LBq5J4if4D0VeqwPRRo+OJpcb3KkVCxgafk
KFk8Jwu7SzYG+689VvR4pXRk0mw4QNWWx0RzJZPpwK70aB2CrL7d9ZaYE8a9FDEY
Tx5NaAkKdBrkRO6R6M0VcXGubhEVaHhOwHedkkA/cH5bcDXPSqgF/5DzbD7Y/nKV
0OR1L/rpQrk7xkFwORKDAvhbaevD1Q3fsV2xK/Bg6PxF9tYTjqWVxbfvydjNFchz
etE6L6DDPcEq7VP1pChHP9EztKP7Yqu32Bnr+Sejmswsjbct5uIjhHtDaXUTYwTe
uqZkB3al4fVK+JUO+Kh+24DPpX9w6AjnbHxLO9SC5ypKv3JK8DPIK3RvK57oABdw
P5Nq70qG2k/Dp2OzHIGE89dWFiaeAHkzcJc0Njgty9WqSaBHYYtPoaoSFWtfrVpp
T/0V5JwflXik1x+Be9nW5w1NCyX0KT+0JzuKk2WiHRs5FhHTRypb//Mz/2+GS8x6
bggbrcU5qQzKMNWe3rt5keywjz8z/ESfRrrqBunvp5bqYYce6X/pUjbbLuYkknap
80IUPiABX1bI4ySgvq5Ze3SCNopq9ySDUipVRPCn/uuMPGlaKkdEGsdVgBcTSNI7
f51/EXWGZgTG59q7uQNJ0Fcr6joMrrKgEaYbAE6pNpMmc7dR00jL5pr0MwSrmt26
LpfkSL4UiKN9IlA9pwK8w9jlTR7nZe/mzDiZyoa8zIW97DLZO5d6jr5bmFz3Xgxv
PZoseNfROvB/+q4GaR782Uhq1YnxiPY+B6U8DTjwqYMQ4lmfmHLocfPjD9+90PXY
kWP9LMcB7eCwWuAa3xDOgwivfX7KBAACuGGEZ5T6Ss9S0slQ+dklgq1NAza4vzgH
gwz6A5zx72AbVNsKFrC6CioS/ZMPw5ZTANPnwfVpgyZxQXvxW9fycqkVda40vXeW
jtL9wS1zlBHOK8qQby+Ob0Diw0g19xQRRwaIocNKPiptKsVULo5/HTNGz4kRY8ei
yzlKtWfJsZHpdm268KEAqBxlSGlxckeP1h/0msgl+iCHQA2QIymDDdOnO0ZSQs55
9QE272fHfOF5dQr1aNorLFC4qIo6pM/L3fFOh5be20c6nzcSNpkYjJ5dcnlB7Wbn
hgg8wvi627RgqljvkIc9j3L/JYVUWMXr5hgSR36X4H+XSKmFy5kHfxd8bngIjTkU
sT89zv7/e9yBHWWfLwfRaS9IQpx8N5NZdB57mepx4gTxrNvgQbyvARhjdWzlU0kq
AsIvjHEVuHjamMtxPWUaeHnoLEt02oElnEER8qWNKjreGfL8mvAFQs7FROIzhmnO
R0fAS6IA/+DB7xQv6ud0MQXL/267AgrCCAxQPiJdwN0Ajrk5Wdg2CawFJU1Wmset
jaj6GEfRazBPDyuSR4z0byIRbByKCGy1X3Bfe3CRPOQbEAMgTAzQGm122CKg49fh
0mkeVNrq+9Cee6XQdoB9+2PlNNfvWkw/nq82VwDB5TFhjIMsgDqIDsn0MClVsIYn
wkHt9nVkTJgzaKBy+OrfbPiWg9QPoRZvm0C0G1Yteisz6yBUjO2JgC1JgTPx3TEG
C2h7Bhg6eFhIevkUUdjp1O9GPFYqGjsjN5QnwZBIYDsb9KboQD/oOX7lLhTwcisB
HjQzg92mUnsKvSF81xFCsBOfcdGUl5XT5qKN5LFRYgS33q8ASKenDcFlA4foM4D/
R8+4k5DqOCSpJU5u06OQR+l0xfbVeIbvz5twWqQhAoZlk2/Gy1heP11ijAOLnOFV
hlpvdvyQmgBkoP3qU/fLuDMIDpHg8Yx50cs71UY5qx7KEbUVvwQc/BngPd0hRJrv
YGQaqBFxcLcCtBrxfDpNnwVVZm89fhxuQOZTHHBxTBJcgRjhai0vv9rmMCf6bAJN
erVvfaMsdWeLjWZzrUQFq+WRGdD+UiydrMQacys40jswpQUlAC+MFP+DqohMW1cT
okJRQ314Lsg8/QQDj6q80bHanbfxnrgF5P0rkq28kVwkXljnppdXbyqvFBAohAfZ
fE3mGgZACMWrLyaM7gS07h6E7MZNM3MALOy596CflzRoRCvFpZxhu8OMR280mgRl
0YIsZkkAyor/CnKiNF6BPWXIOHQOOEYYA1mY0bHlRznrcXH3MOR2bUcD7hTR9Ap0
rc1/D04thaUM0HICl0Ox3vRrptp1nmZNk4m1H+p2w2QF3q4kk6iXxQRDcVYKJoGr
Ij5UNrToi0SQmFW+kSbDvHXklQAYaoiNYRQmGBBOG5929lyucbjyNbVRXTxMvliT
Cq65oejNFV9lFMD2eTgy1X0r8G6WUN9Pt1CmQZkzL5cDrP/uS4bsb+7b01+XDcPF
orpSWFMDFs9B5Qq6EJuqcloHmLQTf90HtdUGQxqX/RuCIkeKTjvXa84YGZc0W/Z/
hlxLoh3B4+9VeyiANn2BkDoheK9aIYEmfiP7kstr8lFIRk16xnhOILtk9NAGOZ5F
v3XWiLTQnA9fr5cM9gYN6qV2r7UyHj2QWN/1oBNfJlvbuGZuMluDYEEYB0dPOnCl
qHlj7OOZz5umnOjRl2LONjg0euhNclD5CCrmD2KwdZhlTaUI3i8uOrU5Dt5HDaM1
2mNjQJE3XbY+e1nyBu73tfatdFFzMhMOnFCqlRFlHohSDlBRBCSqTIDTlzqZ96U1
IEg2NgV966eolDSZV/3CgGfmLO+cL24/Ta775a7B5H9fxXK3mrqaccQy4Kv6oMx+
yLbj7/IAv8b0H8hL3oenxf1XZIseUTUJgoS4m8VtU0yHdx7xiRwugbt0R8XB418C
s05L+KR0oKBRKB0wvaxwnqt4FtMARTbkfUFt/zPZ821zVlftRHMNHccd97asWLOT
K/2B1ARlCCflkPtXZDRgsK+sMw+zMxfKj9jKiSDQExptW0vHBKvAGInPXT0+0VG2
Z1BfiNF1DzWCcsOV2rsIhMRnmix405o7/MkhKJSh6x2AxjYK0L9qVtwX+v00UMgo
Ivgy7i4MySzK9MlXscGxSnY/vf48lz9Ox5GLlJHDR6FUhVidWfmnj78Pb9PJ1ghu
9a4NGbsw5AhVhZ7usMBqvokKYQEXu98UZ9mgmtOauJKXlXBHRdbPetNTvSXssTR6
f0MGwDElK/sNi6ohfb+goRuEx4yMNFYx2k+ck07OnLym92blto5QcEOe7D1en1ia
veZgrYeTLhoHA26sXzcymHjPUTKHUqhrcgtUErx+bUfE1u4eYVN1eq5f9bLwyrN8
IRyUiQ4b0LD4CqBP+4WB5qMSoim/3GcywJrXxrLZjTfBrLvlq2FwxzaYT8LOI7Oy
AYaAn3EcebPXJWeuuzQBQm811ne0KYIgQbrhjW+rcCbkuE3GSdgwa3kurasFznPw
nmwPRtlAVWysWYYGLUYRroQ5+VsCNSPt8F/pYyRGAVfSFKcUQWRHF8N1429ZHmjL
bphtaWtjyFSZKSDnsAv+Mj7nFB78Y/UmvWSSlz/ff0JwoP/r8TujJytnLhEJjRPj
S1TI1z/ZrWkEVqo/eXjRTXpfExeLeGkFydgf/ZHPm3OVqLRR6MPtsSZMu+CLhPj1
sEOkcy7c3dG4A2sfWBLPXu0avc62yOO5M9FrK6/+UmCwcGk/20uZLBfznJ2qKRS+
YKFh3JmvOxZYeQM6X9lF9FO2G+kDHIypJDk0g1s6xOQNRwHF8uDsMbWsA1OEWHLV
3s56VD9mKbQI5xeG60/vlGLxAxljhBawCMgrtRM0WQLeP7vhZH1zsAntY1OXMdQm
4LTrzJ8QdlEp/TChezTrG5wdOuVC4TQlMW4QsliMMnlKU0SosrjgDPwBDxtzhGDL
WBLf+b2lcuRYTsrEu67CXf7T3xj/qlEk8OF/gO8aB/cozoQJSsx8iRORDbXMBm33
gaMRQ2+U/tFQPmw5I98KDjnJQgE9sNh2RwlfmEmzUxhHiq9k9Jc1Lz0KUVi6RRrX
NGldY+LwB8fc6yQ34KstRzM2uJMA/uOGV/EgvpLK/iQ4/fcv44FVZgOHwF+ddQeo
jo1iyg6Q+RClJw4l93H75yWS3ubNVqASNgeAJrQBfHHiHZtLz1X7Jcw5r7/kouy6
uavfiOvoyk81/oQWtXr/RNzrzrmJWwxWeTIp3v+0eUyhKDrIBUE/XCRCTD3ZTdDh
xwZWb2U6U+/DOCxABF9itWKTk40/rVRBXltGOoMhYiqPZZMnWjqnYsk1oXY26u6+
54daL+mr5H57jGBoHf/j4wGJZg/JaEmMUiMkYEIIk7gTrxy1qPii1r8T6mzU+4+I
CP8kgqATscP63nia3ui6rHXM88KrGuxnu19LVyQOKK99mdcDh3V+C9hJdBq0lh6/
UnLdnOgXFHsG2ePBUq5Wz0K7BmGs2FffX49RG9ElGiMajxIyYUgiLDG1BZcbG+/O
ftOlMeKVhcZDLWmktzExbzwfTpS4GR61zPvx2G5DDJQVEs4qXMqKU/788Xcr1fiX
h3c1szOVSRe0FLfq5y3U5m/Fbmp2tZjX0x1U3DWuf+AHvtNPyZ2gCJrDnl+ph7FP
slLbBYsNY4KJ73qhGccvxK1b++t+smgAY9I3vB4Adqzca2Y9ZLO7Q53is0FFiHmu
2bIpn57xou9FzwIOYIVEYbBUXcq2J2HK9FYuzIynoA0mCBn94q1EP+2HX7O1Xz5R
ysvjForD33/ZNzM3FTaeMMoIvjj7k2C807jAIM7qfs37VoWZxuEmWU+HQbBpeOTO
2zGEY/36YaYrJhy+xhwu2f9dxAtWpjhNGXbDMLddjX7TzoqqOQCPx9YBz7KUiIia
suVjk/f09G8vxYWmRJFNH0mcmcSkzfSikAcaSI/2dklNXTUah5STSL0HakQZspBN
uE3N1Vf5LoDFCxh+lzs6AstqyAkWUz9/ns48EI7plu77evcoHVRjOpwq7EFRpla/
8WWJeI/Y2W0yTrhzyi7kS8Z3dw2lS44QOfsQ2jmgpQJyQCXaA+YLWoth7bztYaMx
AAHVnxvN9zPdtbZeTeCUbyTHJ+UXjlQdf6Y7qDSliHcz5oOifiS3VKmJKEr+FM3H
ImxJl3btKkAgwXevcATDOEyPIr4V8LyOcz8hnA2EtwQUoAoJvNzOJC9h/tm3xPu8
xjB2Q2SASMAl1+5y8qeQZYCb7uYB73tT1C1hA++RLPQLTTwA/Z3HpKfJySYuL3zB
pd7CL2U9+yJls3ji4gOdBXborc0r/R648cyamzkpeDOxOhW1fNLiPYj8sUwQOgki
6yBCYMbpy2ydV5DmDLx3XsH+bp8i+ZtxWgCVPrtDytw5edINkQHQKDxDfMnxoxvH
EIXEoQUUO/BwTGs+Dr+M0/b4C6IZznAbunYBJKNL9bPfBwNRLX81M5/jzr3dHt2+
LPUFW1UNWT4YOOTU0usNdSvZkyLW0N4aU8nh5uqQ5lCqVu16WZ8bEqWw2kqzYQat
FJOs5pvswqG4ZM+sEWypFqNq0NZ5gCDu46w2a10oacqx6ZzScKWfx+EBjr7rMCCP
jyi9SiFWgQsrgSe4oBA5ZaA/paYnOcu1DIBIsfuN58RRkIcIVL3RZwuTNV/G8ksR
1u5GEbweAWOUmYquSAKy44/hTg2RLFwLhulnZodEOoHixFfF4Fz7NyMIFaq+vrAz
fkJwPFOwqjhhTDAljwGWWl+bb6RHCH8IKQcv/mDQ+QFja+SqqFVdCmhadIh/fN/q
IhMCIdQbo/d+D8n5k/bBYSsmLZ4OjZAvQ1gnsMTrFOsI5YYDzrdoQZwXQEc2U/Q0
g1lvo0F/JYZf8WuGLThTXpCRm9SuXOGnODMFQ9nqKKE+5Y1msLfSRxc6x7Ldwp2o
09wmn+fMnyaQs7e0n4/vVZjn6oeap0EauLMsZlux9TPjkE0erhmK6tPvFd9W6qgZ
9topiu3wau7Q2ycfnKv02sPqO8y9JsyxJ0ARRqdCk7QLeZ3TM/aE2J0dlbTh95JT
qykRRlPfuitsqWXgom7k494YRqynwP6D6cy6Sp4sI53DTXy1X3VndGEergyBqntC
WRv+mpN5S97RRRxgLSVipdvEuZYAky/g8jPgL4weok0GIm3hLz9eT97sfNLvSsi2
aC60m5Tn3lxcx9eu9fCrZPHBK7PDY4b0JuWsUDMlJ14DhNuXalaXrEYF4+3duhvF
/iOBU/pnAayhue5uv4HkowxglLK2+wo+J5wKJYtP7WXEsZ1otAYtEzBSKyNHOXFP
C6ETlyp9jMf+EKbOGJyVA1/R3vLM/T088Bg/s9BPbZDulYM7IefFcByBxOd7exCz
ZZSI1m+BOGM0KWyc1rqWPMQLoiIixSOtGNCuSZ+2HCRDA9H5oH+845KMTrmFdvEx
Wja/jGLzZ/w7OPLtUADet9d1ba3KKO5Id5tu/VFSt0sQvTDrrvRpRZIV4AYYXEVN
vKpo5eM9n1xFO+C3CM2CavlKoc3wswtGZnOZZ2XTsNg1elmn3IZZZ+9j5Sk6Nhwr
y+S7XxKyk57JEYArpWz7P2wvv0Qytj8BkP4Sd/bIUCmAEOWuplPG4/tup1OPex44
G6s90W1TVpm9CghKYtAZ/O5PvJtyB9pLbhV6ZFN73hb9o8L16qAt9zFllcE32WwJ
9/N44F8nYb4Udg32scEIZM/cq2juI1Fq+f6H+a3db2BPumSiQxNOedc6m9J6VVVk
1DwzDsDsFmxJFwsvpcUW6dmlR3OJwQ/Odlv7CNbXAx0ee6jfhHlaPcenyf7ZrY5s
tqRdFpi7bwfAzVPniki+OuZ8W/NEBnDG+6U23fnJSN07Xic2tn6hT93sI36Nf3HF
fpk+aWTApO145G6Q3BTzFEGITf62hOtPQ/MmSxXjQ+9tBubuTptAV4nDBS0J+mFh
KjhNEs0sNeThE+QvC02ioLQPVQD0RrmfQ+62KfHSubF5TrTza3LELPgwVtaCFji6
bbYddtEHIoEKDNutSDfDmu7+VWr12qUlbDmPPK89bqmGUDg/auZXotgTe9Ri7YYw
j8QhvHQjbQ4SqBB0DvPi7kfM0LlCnogNd7Oq/TFRU55h26u80c971aDfXPwxV9Ci
43wwuZhN0CUvyLBOljVpj32Q5xguPPIqUTsY69XbyO5BN/aGZjAePkLSAKWjjHsb
kN9X9lqFC2vXKDyvLxK3vDm8RlFTjC3pgRzPmc5u1IqBDJ2Cnto1T+u3cTQpCOtv
4LLcnp6XkLHRk0KRiPRsCfKueMZeUu9ELp+EfhTSs4vquvNEBhku3Yz9pic33iYR
KxZadcAeWLz655oUDd9Las6G0+qHjhJFFo7ztemEJMEKZIySzgUSH7Wd4FMIhV44
mT9b610zYaZ8fm+vEvcmf1UmayFi5eEnFDPZr+oDiZ/4KezL3+V4Sq71TDDPuvQB
iI9NeQOYrPJJhvb2ZpMbApkUEe2N/YAx5ma47dxoLRPKgQ8rP6C1iPcMasOl+S15
XKSFgMbt6KSfL8X9b0QlsRHk5D6yx4eYUX+FLlhcUxDTFsmivOzVtnteyx3hUWIj
gZqj7jta9atWj9jH13fr4J/PWveD5MJTcW0ieYkqv77Nu3D3uOvETV5kdTnB8p2C
5YExGzNXrVILoRyk2gkd2HWmBq5PCa0eVU6+FpY5P/2qnERSZnkDwe35GDShOPLl
DKQzaHpxcIoeIMg0y/USXTGYuOHuDYa6WlcjyMtMP/ewRoupNK6ZSacAwVX/slj0
jFngSrk0quivUtlBg03p5H1pgROcTc3cJ88Il1uddjQgsb4PMZ/sYbzCNngrDeSH
tOEVrMB1ZTdiYTNUfl6PFvoDU84rGF9Dg6WT7x4oL+cjv7+iFmOC08dM9l9Bi/py
FYizJnlrwDDimNrAnhqOM2k4g9kOY3V8hE5bxc5SQeQS6MVBMq8+81QmYOzg5YQl
CMm6Bem+M2jIWNj9JFvBqpRyY3WJ8KRFKIbhB96ukiKc5vH8n646ek7wWEzC/Pn/
gRk+bihGnbsidVjmPlvUwdrMLGvTJ052bS7D2s4oFCMvI5KkUufu1JHydYREmHzp
hbuWJaMo6RXImvSyF8U3r7LY5o6XkJkCMyAIArYc09BCfw+kGbL7a/zrNFtJh7m3
jyEhaUy29Yc8qS3skl8DFY5a2U1ZNwG2dqfCLsx8uZertedCBj5irkt8B8jRBZsb
mobdB94eRqu5bnkpqs4H+3gLi5YDFrmc6Yuzr941ncZkh74aVRGnwjLA9L7BtNu5
UuE3E6aP2ZceE5l8U9mxTseAur07y0oufpHRr8/e1fSDLJ5OuBplfpdSVjZ7vJn/
RjypoWSV5OhsSy2dc+TSmRU5U7slLEfgs8EuOpVtwub69lgPzsf/WaIVBaF1dDbW
CxKIbUofKwHFE7uNw9SguunNjsAI2CE9pRW3dtVuBhRzj6xu1RlbWhG0u3ZAqMs5
9RvZyOucH/5BaHefaJJC6QvqObdFyaThH8HCojJCq2AceeqjsWysskoIc39LG+xx
SQGDB9hvySBtR9ko5GdliPTO7zfhjfvneb2oDfbYjHYJ9FPGWylQIu/GBDi5m+S/
tlsmIljXNtMoIZ6tXwiRtneTIlcmA8pNtpw4w97pEdaMGKKQ8cFXF2DLQt17nMTk
wVQdzcAxoI5FMSkbI3n7edInpg3c25SolT5Js4RjYZS7CE8Rddux8qHfV84B0hPH
086NzE+E0t4vCOG0XP64X5xSV0gmqsgNFXjfGMg5r8kIgLU4dqD2wJTWJDo77XkS
eBtTJwo3XO/l1gI+pKM8Moj/5KRIgJdNuDfk81m2RlHC6vvLtrmP7tKvF64DTxyk
uIQQOrxgCMPSQ3yx42JwErqPYCApl63aw9BSil8KbS8gBLIfC/CemQh+20BiSDaP
ciDNQv0D1MpOkn+IQkLtjdPKCaRui+YwFlr2X7wuYNe1lv6hBn3qkjNJJTuOaCpE
WVPneKpJ4Q8ChAGQ3AVznd1Zbx3Ug3t6goMA4n7BGk/jM/ArHbVbz6do22AZ9vR2
Oasg6sOnTbjpnPdEu9yeZLnPUDacw2qeL1ZZ1RmPIOipGz8KLOkYW9oUTNacfAG4
flVe74rww1T8AOdUlpeoOR8yndcZh830nLZvOYoEG6efhdmliMzyZCadqUVWkIa3
/NkIC4Mj91GKaisrO5ynr6HS3AnLAsKHiQthfHtuJc7ft/gAVSR89W9KK2xT4Qik
aHt/tYRem2KoFhPB7edLRqDytZdFLwJLAIJQNeThT+w+q/YQ7f254VOLI4twYV4D
zRNDAa4NK+60Jksjgr7A4gntlxUMwssJvO/bTn+ULyyRFaTcNsk9O6XN7aN7Grv1
N8w++Fa1D9eb79vSMRwepwfYETZL43vRp8Bfx+dGXi5sunLDEBw7j3wnsP/eaoUn
2OOZ+lCSlbF+l9uGcCLyE99x/U015RYdhVPb/pQvQ7chSSJI1fmTgvhAOP/5Sbm3
KFnYv+EBTBNjVT1L7nGNUxGw5TvJSB/f4EU9qqSmFGOEqmMdFIv1eJUx9Io2YBlf
Fkq60LCgrBV0Bnu0apnZrFdm9n/XOwLbR86/Kp2NFjtrWiNrXzWfHI51ERYqtMRf
RJJLk3/XA/+YSxe6qv2Ie2ORAIMmxcJXrHw/VEw4YCJydZ2ek3axcj8FKsJu4mGt
TS80lTS+iRO95jnzTObcjSful2vU+QReURSHyAu0zs4YiLjI1ncxh6QYifG072KS
90IcsO5Sk7LmojUyE41yFlqBZcgakHTb3awV9iF1STq65z6FfOlK+LoSyNSkQShi
3csct6lOxds1YsFU6fMRD8riUb95LnmyUPOToCdV2J03ccveEbDur/N9F7/uV3xh
mmBlT+jCV/g5s9cakYm5EY/xy1Z1h0mdhthtVZysZqPHz0rowbtNtjBWKlGO672/
+M31v3MGBrbZSsIfkXPu5PrnlIblGgFt9nQq/BoCtvkZx2EUaNzeS7ibPFUvdOIm
/+uWkupBsOVO/fTlIRbMei3RPFu4efyB/REkegOOq/TwSd9hgVa3BWqYJg1z3Znk
y0hnaFtmqJ1L64X97EA+wCRg80SENTe03Hzh8vxIh0UkzH5CNNwaSnDnyAGYthGX
Z13Ah7FV8ojNHV0sWTFE2SZL129GilIFV5gyHEWESVU0Fmpl5sR8kcxk/3AL/un1
0SU6cYu57uiKYaR7CInhNze2IWyVUXfK0oX0mJpUXZHK4MVivfgsktYucAHd7if8
TfNgqKrxCpT/2NcRfvHCP+mW4sqDNqm1gtUV7X6QmuboootK+9YzioGmqi8N4Mt2
tporilziJ/NYS5mYhTYv23667gmPm5xk37Ez/nsRvLguA7++bgSxyLWPGPaQeD3D
7U/upOeCI4nXWuNpoldiaIJZ8Ju+gRLA895akiQBN289eHCAwjhGBzRfynnn1d1O
fnVtFMARQ+E93da0CRPKxUOgqRsm01WPu1ABlAO9E/XOYZOctL7wfvlOiUi9ljbk
VzicCLPs5bwUd/DRO5eAmHA1O+O+p63j0mN5M6tGZwCwjIYbFrDlKKlozOvcm5iW
H+A9e/3p1eBD++ygzVS5lTvofmUBr+dPbjQTif9wlx1hbV00V+urnCvF+lEvDzbr
xtu1r8ADEC4vtgplzKOo3rQivVqsKpldsKfQEaEChuCkdf4SeOXPjnXFIVbllz3x
tK+ULez+PNaLM2CtbRc1Xt5hKs4i8DfOoTvX7j8bRV1n7oxq5EF0Z/yXXX6zv7HC
7j5mSj7LIl3/4ZvGc8g3y5mLH0eJa1KkQXCRn0/ro1V83kUu/tWWkJXTk7EkPVU2
0Tux5oxNhxh3WBMeV+dBR5ddDnACbzgypSMtjWcIa5VkkB361euN0Fx+Y9tYpWCh
RoQDVZwzp+luW2KWK/kOk/atfYj1qaurEQ+90wb8YMbs5y1c2yrfEdzMHVBAMziq
Ebp3NCCg1y69BLENbPVuJdXNwu43o5ULHBPVWZYP2HKTSZpsqfxWGBQY0ZrumwCe
5Gr5Gql+C/FNY/Lg443g+D/qFdQG4JKHM1IH3Kt4ydvQiYAqzNRBZQfWaj/0Uu3s
2yRk4sEtSABIRN76J330Y3FPO1KO2N86f7YqOzZHqO7xSntMo4ZGCsm0uGji6lwq
Wit5VaBev1bDWoD3pDFXpfX7Guz5K22rFbylIWI61DeEPB+EVS6oESlVxolvlwRc
hOJD5bDpmTCQQz4V0wd8sYYvNrZ+IzkkqrQKxdGGxtvxgfpyEKEEQGPlmFiwFry2
kSvRb3PI6sc0eQcaj28UTSjQmPO6GzfnH2LRan4CBqJzW5/NHz0/j2JvcoJMaUzz
FLM3XeyhYjEqD/4koPBDe7TU/B/OfeD68oicyGuMRgV/XY3dB0nXp1ggR9K2yYba
OSve9QLfnE0EvtZ1btFQUzbveCXr5BDDqbAtAuPgjJ00E6C+60rzFwK1Iz8r2KYR
bN6YbGNsY1raWoJmbTsSyO4cR3+rsbA+zoB2Hr8TfIMoi5Zj9/xwg9mxZBK7sqa+
7gb4hUBgZqSrPRxyVUcKR+kDlYS6gX2tRU8KXJJ+tf7ZXz34AIuprUI4X61JKjvA
nbIPMXzB664hFkI6Uu+RisLSHPUTSXzkJYf6yXCZSJbrE6kQg1hfQch5ozUkYXzo
nHf6ivyDiyROPk+xcxlpnsx3aK+sQ3f9oZVe+fBZg+p2tthkTo4AVl/xxaCpTOq1
5sCPTFm31hYe/M/M0GNZBZAvUtT+eJP+M/1yLnr1G60lgZDN42sjQtaZAcCG9moX
GOXs4r2yBgMwxcyoKVF5qfLY9p4CLOJpTdWReiKvS0t37KRz5pCe4vzURsVFVEca
bMe7EgTDc479zssWklU+3N+8YzzDBRCUr37j/z8wIJLBmlsc4ML86EjMmePRblI6
8XkBqhR40SMeRzlWD4pONLZ+IFvxxvaeiZ+GEI+IEGBLqt2ZK1FXk0DPqFsYNEDd
XsreySFCZv8sDQJAC7h/no4eknBmHh0cPdwNqfdzwu0lYZ2YOwVjy+V1iP0M4PzE
b0KsgwWkbcbrgv96xAbD4xw47pt1Co5rNOq7i3N8uUTWy69w1RVVYC1Wjr/8iL6M
ky51lLgcGUo9VDUu2ulieBbcPg2NvjSfD1YK7WOrOTteH7EuGbyvJtvEoRFI0t+n
y+bbx7SdGiD08O6KlWD1n91c06BhUAiKCgWc7kRo8ivxmQHwbvqGc1EgyCevmod8
nwJ+b3k0AFGT684qFNiJ1/Q5YxPo4SxrWjXfcCJYmd+mZGZcQHsIO9AYXAvOYTrP
iBiCMspboa6ANOALI0hcqMh0PUXoZ11i0edR5o2ACgDVXp4SZ5eoHphBQEpxTiSb
fkOkF2Bqaf4zrxUhDKaYXJSnF6JYhSlFcBd+aeFbuxRJoy4FrIpLp1D7hWDnUMfE
6nk2wth5fR4khOYvAXcTAlAOsRkWMcHbNsmTe6d9x/L2k5tNXDZsM3HV5fVoHzlv
dF09RNkktfyvT7aKxQSQXxR5oy4IT8ZRmPEt0tUcgmSspmTeGzwG+WXJ7Du8/3rt
6iUmNk8XWhHmFwzxYuUML+xUwJUgoYYlHZ62EkunQV8v8EeEwoc263HfoKZEKUdC
Z1wQP27CcdUOB1REnpmVx+YPdLfVkwMT/HFDc5BIsh/MZemqg706Hla8g0cQ/vBR
K4d656/TCJJ9P0F3snBABs2cZsrNtmFw//lcmaBdFOZrH9Y5A2vfa2E7E8RSb2rh
DqiLMUCc250pNkSrNZ8nMCidywnG9ew8q7kyhlnRQzJ2ttSPdfeA7RQJwRUx2TzH
PdubvS/VwsLyaJHft/O8El4ixPqldrpHV5s1pOcw0NafrdKMkfRQE8BVOCl5MTJn
843667zO3AQDT0QpOF3EV/t0sxWsM3EuMu2uC93ciAq67rCp9epRSTfklRIDSVhS
qmS+4qnfe5HMHHWsxovZdGfhL1SN7XqIizhgda8GqvpzapWQKWo1FeCVVJICW/lt
98pGowZFgkpzL1Nejph5J1NTDEM1o04A4sT2UsY4K5nk7ekHVbE5Puh0sDicPII0
9fwj+PY2TsqPA2vGbPNjMYIro5VcrBy1XsBNNIZZ/dRwQ/FcPohDWph8Eu9acbNz
OieJGFFTKhnCw5vVwQ2sF1WxhdEWOZLMim2xkz/j83yKJshLBuDepR9xz3neLIHN
e3CT8PjOseV7uB7j2/C4DfIhRpc95CrDyir8bHmHU2Tdtm3PfBGTVpkygqkc917P
5NiwLBJR40yd1Vo1ckaEv12CNijCzzUFCfnT4leAWeK4nCWZH/xA1ZiFX1hyDOlN
TfjSvW+qHSUyafAwbYS5vDD6rbhVbupZBm5iJ2I5R2yZHlTvFv8c+q/QrCL4oG5v
YeXKLEFxfDSabvFfB6YJe1qMcU2kaiSl9k4sP0URZtg20sjmzOfeKlpp0e8wiiJ9
xU3gJJQDqV+Ifg3brOKUEhiKpN+6vlPq3BT2KcWQxl3gKxCY+xL/4ZznysNodbKO
FkwQBcrv10lXWKmU5UfOYQaS0DdPKp+hQ7iSjKY7Bu3j9hIMu3inUFVR0r0DGEla
FbHH2jIUi1znqkE3ht4pPoLFET8KbxJ2vKTgOXN/hOe+uMzxEroV7CEIomQyofGe
krK1wuhh+djsZ5WE93cjTlEB/aW89H/d0a1X0+PGyXlcW339AINzhfJU8irs9XsU
4BgVdf+hZU5PacJ7OeyYpep9z2z5hujRJDtxYmNeBVdYn9AKPZADa1A5P9cJxwM+
Fxq8P0CobyEA74ehnBVMX23Msm7AiXQuILQnfoLukU1Jl/s6EHpArlWrK+Wf1tNi
LzA5Qs9DW2XE9U4d+JFPnpYYmcQ3FLl97Wbv/b1eBhebZrlHah8juGIncZzFSzJc
xbnCQVgSWSeCwdu9hzROcgRFpsHfrSDfjDYTAVLXO0l0hROsXhETgfJowQyKGesc
mMxzNDHT+l8UM8DMrk+qtfJqpYfYxyM5/QRB+le/6+rxXZQyGYXuIQPLv807v8xO
9yLhj8ibJoFWFw5BnEH+Ru09bNoZYM9zKp+4DKlClHmd0ZQNGg7ZYLaOzFJtCyVK
r6tHXlG6OYGM2TvTbcknufshun8skkknbLyatXpyj8+djs7n3nNwnkDGN1MzZIfH
QuUXkcGVe5tJB8kO+OJsFrQpfDo35Ne/B+aACuzE8YQ2mFm0H22RuTstbJBi2BvJ
Hi3fB25imKcTotd/D0Hh2seBNo5c4euFOtMh3b5q6UM0xtxRe8usOfYd5qlnrc/l
lqTZUyWiTH9XC/2WrV3C/opP3drPZqFZuCk2c504n6djYcdEQQVkTQcLa1QzlBuQ
IHvpRtwpuR2/t3WFAbuKKILW3Yqe1RYulQ6M9uiWhfU+BipX5WNYOHj21xLMT5+s
p02QQTV0sZWpyaKyc9qd9GKLLFCkNutAnViddF44+ZdFLJepc5bqpWekrRd5etj2
zAPFuPqHljFrLtfRkhsBPpZRDnlue87sC7SZP348vOn8t8YOYv6VeBmI80dwiUZE
gUyZm5b7oeamfkcmhur3MKXfuZ3AFsPJtv6ArB/G+YoQ1gqvY7lrs2x4yFmlA3wp
JGYRKr6PtbTg0cVsXxKDW7bCH8XNZQSL8XszeTBpm+WZLjqGD5aKTVEeWHtwE2RP
ABE3/NzoaSI0igeRyw4h4HG/ucpySBEBBvRY0l/RBDnKdsKKC8xz63KMaoVEMIzl
QR0G7vzGBKzW487rWIx3QTFSYhLfpQ37HSh9NI+TN6Mm776wujJ+k5bZAbl5ywVC
kj0+Clhzc3R4oQcPze5Uqf6OUHsr12IN8ykkJWDQY50UNHIHjLhjjhUyEYdOw8S5
A8BVqOSqR2qnR8zrlzN+BdQuDw0ZMyionp3cgLY2+2L3uU1T82i9x/PQN9VgiiJA
gU8TocQPnB06eAEj8M6he7WXjLmqG9Koblgfo99OW5jDPZjSn3ePs3aNRks5ZOhI
8F/Eg1roHIWsouYmJe1GdteJoLBbZhZytdq3GNkxblpKhpYJW+r8vQFQGLOUHb1J
hT7lT/nPM1cAhDUhJAHSltHrZmRw0KO1eKJUx3du0tDVumOscGG4A/NkDHkrHP5T
Tn5tD/cQfbhWWjHQC4i52nmFfPqtJvHZCICPy3lMGThljo99Nb37fJnL7e6Uk0o8
0UREEJYOIXwZ5vnieAm6/5TPUu8b1fscuaz2MzLoNyciSMn59D+eoPDwY0fTlkjf
B2IdqRIpbQbHb78pbykb1Hd3j2K9xzU7bP+gF+MrSvMlufAuraSHSdIynZSIUnvK
enY54IbaY/Ur1EKY0z83DLiuL3QvS+JVKPiDEAUtvUkja2ZFi6+wBOuDEAwIIGak
X04SuGrmFpGLu63zx7X2oHqTHdA8TYo9qWjgKMuhD6/3zukfWr4yOe74HOQdHWCc
zxWLgzU9PoWWVvOWsO9goiDCnBDNYYxU+ruYGxZyk+rJ0wi/+wqUVfQbJS+u4g+p
/N6vTCJX2tPH/A6D5H7TpzX3dciLyj5HQSFXd+QurrMDBtxrZEugqX9RcwEGP3IS
IeYJCWet2gCNmuuwwmFxEUU6VoQ/V36+5czhOjJHdX4FLAAhZ1sVmS5oaBj84AH3
5MKjp3d1Ob8VMCsEBHp9sTpgzNrd2dreb/LFH6jGySGKYNa3KCbOVFAJ37OU4feo
lW5CHNND2k3UOpaO1cz3yH3vY4petkokHUAbu4Oa9Jjrxk/2dAFdDvAFt3v5t6B+
5Nk/N5yrrWDG6KqOVdJPaKCnjenX/6vVu10wCQgx0fA1TSIWOYV1I2gPvzzr7/Qt
3Web9Zmsnd7YazIKJNkl7y9yGAJytfw3f9a0FEyj6iRWmeS/ifaj0q3u0EA2uqS2
0B7/4tUrqz7iAlDlMGyxT8EygOltaFIQXFZ0ishvRKBrFp6JCh8jDcB6kNcdkn/l
BHkPcSOKc40VWgqMPM+25Z0N9nDTxo6y1NSilCEUlqW9qTCzL4Klslrv7haF4mZb
Ss7mwBGoDm3stKW0gl050FzTpguxidSvod+AkvsdlMxqSLV9QfLoDXzIMFBsOwkA
FFttsE+Ryl2z25xJow5uNFFi6BpZm/FirEQN86wTP0g2LR31MdAkf2of1Xp/zzW4
6Aq8hxuY5ohl3qWAkDFHvatd3P331kOx6jToSV7hilbbGjW2jR6allbafm5PJ6Gt
CWgVHrmPVySlEbsO23oeD+K/VsJ0DBwVDkJSu1Nnh8lLDG/s89hN6NY7VGs1L5at
ZbNTTPzAB1/HV/bUgZf/6xmMt3kL1Vd68wU24uLX3pDoNzs9urESZSkbP5DXJjhN
r5TcnJs1WUQ5g5nHtCRLOCVMNBRTr8fT933Lbu1a4UBBxve709/rV+LtinNE2eOP
dhV5nz5VQnYlhnLkb9JKnlNZoYqcfRgyvCvTi9SVxrpI6tHKf1XXF/Rojw6V4gn7
nHb1Kue/QlGfiCxrqHEX5b96zeIEIir2KaUZ6d4GZNLLqoCnxzvsSUBN4YJtpbz+
tgoxb/qFU00joPvVIcE3CKmfyffFXyjaDpaXsTLdRINfnkUuGFX7q+cYUT+kEy7m
/XERu6u4ICSvllqcTRUoTjr8Nl81Y/A1bMt9WSIFW55MVG0gKPwms5AUeGAAe1ju
Wgdw/xgQAlCCwpHeoE983rQJY32soXxVCotT/R6UtnQW7lcrVZ22rWUwqfL1BWDh
fH4enCCOd0mUXgj+m3tl7h0NgyDuLOkp3AihOBkI1cKqLuRFbvmTP+c/sNjGarj3
Y9gbltMl/oKlt0kT8FuqTN3I7nSr6OaoXJwsVjc4E++RkN7XjjEX5T9qJmOusfgY
UROnWeBbgcExX9mqHrtC8i5xv7sJska+ILPYDWQNZJHiXfuxo5xcKrGC+mvdT0/t
bhNylxEzdjSlQDzK8A8fWGWRIBFVMMjsWo8SyNhotMJQ8wc0zeyCjWudu6I6PhUN
McIfYshacKU7V8qvjHXtFp35xNb/KZQKDndZZKmVfO1i4JkZ8LM6aDDYDH50dnfe
sY2izbeEd31jQYaYFnn07iMfYIL+H/hLeglQMrZa2zSpIytn4FH8vZxpxdIvPnI9
F3H7TqX13boq4siB+UKKBR1YX2A7SAOc8sAUijN8OkxkkoerdPyuQLTH8x0V+1eg
MLF7W8RmYNTGz4LXD0rzlXl2IzACLXu/c3ZD5VoKSjQvOBjsgUyvk/5D3CF2Bi1l
L9N8uSg2EThMl86J7lYnzUInKjxOl6/GamNATodsKHQHzeZV1WWaG98KOtsgpuIz
Xva64nKzGt1+mBEHkDXQwubTvgE3uXUx+LEkLE8FS8StKjCWD8Vv0AsYlLD3TRBO
5aZpPzNagD9G9II2S0n7D5vVVyRsP8tboHXkgOdv3mT6jHs9Bqd7Fi64cfPFmH+U
ZnKqtmaTiWMUziYtXmme8WVPECpgKJQZ2LQlmpr8KNQ0PJ/SytAPU3lb0iTBTcl/
vuYljM2+xyW58xzW15jROG7f/GSffgewt7KuC6ELj9AFIGIEqlfQEh/2t71THW6p
ZVLMJahaA4T3fMw5efHVnVQvfkZo0cgek537+rjog2eRCYygac3XaLWfRLEs4mmM
Eph5/v/BN0pGxraDAyrOikJkCh/b1mPJZxGsbFA4jr3ZaVtEh+4TNAByr5i/Us1C
SYap93I1IiAoR0aD6y8Ex3367OhwLHCz0VVZl/fH1f4vUQ3e2CbSMJ/1kAp/3xlm
add1Dj3BUF4WnQySb/Yb2dJTQ3SxzjwTp8tpZlZa8z2UZeZ0IlQx2sYSV78453UR
3+ct2Z/yfNX+z0ms0k0qQRGpO56Wp3JABrdNFrQ1aDNg/s1YG+7lQcMJ5gYAp7FM
+/Nq48JWslc1I37r+HqlfMpE3/Z2VMxhNu45o0UmciT155R66IEjZRHcCTRgzrG9
eKUQnPNb66L0MHXAKuGQnLabXeYq6DbGZB/+NGrzbP7Gzfr2wSdAI16w4KAFJ1yE
Q6AjS7AbiAvkwNtw++z020AvgTnVGXw1yjnjRQtgRD8RkfwxNdw8GtDEtu9go9nu
rgVQMdXdIeQPG0wiDeOwlrO2HZ+ChiZVnKjOQzBMiTUCpEnRS8hqbVwcV+/tYZ2Y
u83Pfy1Qg9ymjuah9gkuiRAfHeSkNuXR1iW5O41NXmxIqgaNotTAX82sDczndaIa
NVD+EUyWWgb/7QfNAvP7jJwfd3C7NXVdeXvCgjWQ9JeGn3pw4FvgXTbED1BsHiab
uW8uEFSLX68Lsbon8SM1QPWmHtnCGC+DxoDP/TwrEpitGGcH+LnXXPMqG6BpTGZV
MYVBSL4Qs6pDN+durpEvip9Cp3FUMVynpkWdgMIj75gYUc+Fuz1/K8lq8WrvRdcc
H5apTwzgH7vcoAdNL3IehjmhKffxlwzrv2MMEltPHKG4EherZ5f1RVMwPQMV3ogk
H02jK67xkRFWtWOaSBQGZ2dyQHPC+8pZerKaRnyB826YJSRN598Q9DuglVnABu0h
tJYWf2pmyBzyOXAzBe7pzedtoHp2W2QwjidKTBnQizuSJx+uOq9sMIgruYrhl/0q
r2MFXjVx96GXK57hJNCy8auNAxILuvygOoMaWd+1B3Scgzn4gPjJwqBY0LhBrgQV
/PjNULt4keApefop2DEd7XJW45xcwIMjdsf63blzPXIYn1cxzHdHyzRJ+RtXLtPv
hngibXA6yBJZHwWoexPlBDZjl66/Y/Csyn7cZVuLSt1nlkyfqFxUXVDTAZ8AoGjB
M5KkD8HakMbDUHC8yodOdActoV/LQhw8AEaBqxR5Z+AsfxpFobIVgFvAeVvzD4TE
tig7x0d1GuCPTeuMhkZLmmQqOX4RmqZbERW6WseyaRnpa054GELzh13b6WgRDl0+
vKIIphVzBOzIalLopujQT4O0eUITS6V4couok0qoB9zpka1sa4lMQPojW/3fwIUh
LDzekIHvSH0YkFMqxaXkz3n/Gxa68znya5xwB2z2TlTpzctL/eLORQWpHl6LbrSb
s6Ghwh/2ydnnYwepofaUHc1vzoNBC0kcNZ688PySlYOt2KqdD1bWm70NtPpEWyBP
OKTYRCqgimn8qdJwPVbKx3N4B5mkVO4niNgP4kSR3FpV8fFfC0+L48AsryEIMXaS
QTol5uH5pi42UafePeCuC3xdRk1qvMz6OEbGACB7hS96jR9ukZLoPPXTc8qcF6Tc
7r5PR7Y/MGxnSHaRGvnU2jI2qOXD7HTCuxZaqK/xKOPteCSmmS459u2xPUV345N8
oMw6DB4m64nl1da9SNBqPVGJ+cBGXC/NqePl9LWqwNfEFwKKMo4qrkWp49hXOWM8
Xj+U5yhRnvh11RVtkNGMTnP2iGQH40PWNeYrWqzI4Qu1DfsGx10tWh46QMuYAka1
SuQi0NY/c2y0qi3zkVgZ73Hz+76dyqbqbT8WAYKBcAwnZnKI/SJ5MEpa6flGVwF3
2L0Jg1SxupFjKjVlLHLpwdkmSbbaHfwagvUZk9R8kPZPEyBz1Nai5TTaXfQXvON9
S4pGsZ4dVKOpHlad4cbms7AYa8NvVVw+eeAunLjkCff+ZDokK5DeUsGZpDCJyOCb
Q9MNpZPttToo7ZdjtopUE+DdnmKCEMGXHGQrOil9TdKxDBLW0JTdSxKWTXGE6jTh
DROoy1Ko9f8S3TX626W0NbOudzurtuZUJGuLvkZx/tP5n4DEQ9ccBVJyzq2tXgOH
HhPoPvWdKT+OrSOLkZ4nCL5uqZhXvAx94VJwdTh5J67J8N6nS5q/dn2E5RFM8Bk4
ktILKR+kpukXqdl0uB77NmTMOYXaZ98bhJTJ7tNAnq7OUjegLu0CqhGs/kpi5UB3
MWCLmKazuxayKVGwFe1L6daSSSpshiPIshR2J/gkCcuSvvcAdB4hm4pGav3re61x
YdvMzAB4RePJPDsmfiIvcaz7w99Kb3YS9XxR4mygXct6wS2yD0mD5aIcMlJgg6/S
HCHbIEVtPCmWSab3nba2agrBZvuiEExXU1AOf+3JuWHAEDOlvMndCPF6nvTPWxtd
JuIQER1ml2u6C7KenEIT6ktQliLxYIkpu3w2bihXUfInTLA8OCncSwkr0mQzdlLd
GXeDSG3KQiFQYNOVphs32KlbsPmitKWgr0G30Ddbt4dXRR6rYf5twr3qHLp1eVsN
RPT4QdLPlpov9CpE+hwfli1l8GU494SrFFUE2IN5L50y8QxMg0Ju90Rbs4XXxR4X
2iH2IJUxjVPyWH0bUJoGXYbsk9MZ8+8/aDHwgoXadmhFcY30uCyJTHZvgs1utk9N
Qs1cjK9vGHwr5ws0tonhQkqhMU6Q9g7cTuPiqjrcsOv1MrSub3akXehXq1oK3MMC
EjE+1Ke5iv2s767QueayX9CokchOd+psrhCBd2YrqspshL/Veb+ypWDzxVKHP6Yz
GETgI3HoN9WP999k7S9dKS047jHtAvFaeThYJen3fx0wKVBBzPL1r80RDli4JldO
QndAiQwo/Hei1NEW9yyosVki5ZQwWWemhhX1fdsdIxTUt1n4RIzsnmG7+QNjMWPF
N8YZPyqp5OxkC2bvHE42IFfiZdUWXEF4Qc4ToIVquc8/hLjSSQ2VaO5Cv56hFlj2
kGaCLtGIoBBXDWpC+luytdoIm8DW55aYRJZ60nI+vtaefH4b44jgNWDUrmjiLU1+
9Km5vDJQL/cQNz+hAxJlE+RoNY8mHd7hmsIvRGm4BiyF7hPvQaz7X+K4HAMNcxGl
POmpxCNd35BMowCqX2He8QAWlelWy8R5qtZyMsVQHJcKb59nTplUd+HvM3E2G45C
MGlTH3ri63PrJmq9algsCutQz+7bB7CfNKbSTZi4ioSWNl3snyzpw4uI3Qm8jL0v
xJN5J9UG0y7wrmlroBmdTFg0KPnmXvZnR4AWgq7VbFb7m+DRWLK75b/ZRxpjplTN
F3H2hijlBVhiQouOoDNxv9BvOAQ8jUUO0sTRcJ1nC5M1hGrMAfnn1MlHNM1FcbHd
yWZbxo9bjG8yTcL/N/cReT2Hu22kHW5WO9AZ1zgKELUlyoOkliDOwfPwIinMhI6P
LBXTlgrLmzSUuuS8WvwGMagDZ0gr/ZsS5HILeueP3YU9Oz7tkucIcGYb+oz6J+zO
HbOW/dw3QLgB1w/PojNQl8c7WxcHrXnURo0SX7E+nFfpNUFI/fFiS6Zbvz/d/Tjb
S6xx05+mB87pzsxYW3XUG6d6+UMfqPeAiFc455+Z1sPbqgegfhZ0gMOjqSQvoOIR
Yu7TpY77tqvG8ZEqF+mjesS4x0P9i0W3lB22TuNkno8f2tImWYhOUQhSOI+Pww+L
mDHc98AFUFTiun7VflfKmoyEvx/Rr6HIfz9oOjAEVtNaGEZ3w/uYytXmkdjryu2u
L1GjdjjXlbPuUJwNkljYb89zNf/rGEWTn7rb/y6adWeHKEiPi8qu9Jqj5qGE69ln
JLVkbyd0vUz2nvgWnnxR151FrjfX+iq7JQsiTlBsJmMSnzhYWZd+DKCeRYmaSYS/
f3uwainCthzHy6O/lc2HXqNQB+2XdQUPAKyzAKkVzW4ulnhEcc32HxR00v87Giex
Msyeh9yQFO3lVTFt44PolJwRKPw+NgUlO2ouruWyre3VyoZaeuy9kTwiUn64fu5Y
Mzv4w/bDlKGm5vii9XGaAaKqpASE3uDdsRaN+Mebk7CThdtGwfQLSmhu3JTDR5ZS
Ei5+gD+nbT8O7jLshfnY+Vt6meqHZTt8YH5zRVWoDTpILNMiHvJ8tYXkJc3+4qOJ
ARbA2uRr36J7LfLZ6OEO7DBJH3chaEjbaEqfhG1CkRjxSi0C5Y7VufiT/zU0PH+z
NAZnqJV38mY/jSdJf21AaiO5wPK+10JhDHCOEc8+JzrvyDEXUAA0Zh+4c0j7kpoE
6yP8/C4AXwDOBgdQgfmhLwK8Bb1S6utDCIl2jWxaVYBL56aVMKU7OFh7Rk1H9itR
g0hjGxzKwx0HDukPXy7ds0Plva7JA1NdspmGpi490cjI27K5W/mov4iHjrwtCimv
/fl9jy8CUjbAI8y93wG8NOHAiBKg7i1/KhLb2+I5fPNIy4zC52UAN+kR2mNPTs7G
38L0OZLvWW515NX3C3r+n64R02VfyClb/GMNSe2IbNA1pl3Y2SYJukJEwBStVSpb
UsB3PIkFmd1X9wMaYaxsZV6ErRIlZhx+hMoCzEYv2lzk8JrpcNRIgtXQEgp0AHdy
hYG2MKs7xQ72f7MSPxbZsJFV68lCFhtljz8P+WwoRbap5SLBY53QeO5ze/Uc7tLB
/Hr5DRWUGy1Uv3TN2ta42sVDwvNfav5g3MWgJUQ/cy7qhl0HHWOu2YOUUzgmbEcF
F0ZAR7PLfEFyE/jnLwmDbJK4zLTnbKJ00MZFkye3LqBsK01FSjwhFdrD+cuQ/VBa
z+5j7Mtkbs5kRYrSeZQvbXeycB2y9pPJgd0z8HWR8p/iBTsPa2ObCBeeEgwHfE3Z
XOSivmp9VBVDPE6iwuimZDlS5WaQQTo0qu3IN8qFCk4vFAWQV3sSxTVi0w3A28E5
IF356EIwKEx2BJ5mnEYfPW7V6H07UZ9oPZM4w32odyD1JxMdvAR/jJDKEZs9iSD2
/esTmvyPcJYczJBA8Z2b/qZ4Oz1DIoMXWlAk/biAsBg8mEx2+l8T7wYn/le9LIte
/aXLfUyLNsayBmSSb7QUzz2SSS8zXzTHPM0usQxQgyNA9EC4qKaPYnDPNAx15ZOC
v72WAqQ5EXSY/Qb/O0p68wRuU8ZJCnzgxU9NEkLr7TSWDIptknY/ZkTKjnq8kN27
BD3Na1kUIznE8lJr25KieeEflybj083fA90QAgLUJISlzuRJZdy1Hm/O0azm6W/B
CGqTmLQNVKZtBhBG09ezn8UEoTgK2x8hIhaXQZkhcH90IiYGUePRlvabPQPgT52l
7xqxSF+gQ697ejv79l6MkhRxTrq6n40t8DcgX0cOyeUfj+5i2yaa6pKticW0urmC
dVQbZ7MoPyFPmPcKJpAAUjnXT1hHPaxYY4+V9+dYQthnlMv81yteZi2UVIC4B07+
ugrxXkc5asMVpjZrVIMf8CXCT/DRi2ow+TgK8MiiwmNXUESWaEw9rulY1R4iO4Mf
p1ashsabQ5w/VNij3aEOMVUH5m9liunsyXRZ46nyk6A7D1vKPoJjn0UwrK2hXe5w
tzMs1gShGHTpnu4r3u9gqV+lUt83VtT5STYKwCyjW5vZYbUOuSitRLgdoO1d85F+
oUjW4wvQ3R72gF4rU9TJVSoi8JAxeDJt7L6yjhWVwxTZIsRbD5yHxYwp9yGWsoRm
4K0fGLbMEkqYypS2QOg05EMOZx3B3foX6E+gD3vWBmQNgCrxemXSG5d2of06Mbli
Y1RWE85pAenN5Fhypr3dH95r7zvitqLmyVsI3/EM6R1ekFBK675uEYWIX8AWSFuh
V1EvoeaugcaZEbqlwwqf7UHJW05uPCJ0LnCHhKQDvGFk6ztURUlSpl1V+1YXaf0f
3CuIx0yG2TmXDUDWY/2sxbKkpN2YgDCiACFeTE3fLQi5W8ptaoiFd1ISS5OFx8JJ
z7Omz1BfxSfhB0dUpp5fxuJSq3Tm4q+ZFqPsgmWFUKu3DCgMmAXVkAVWgrzAQKcb
NCZud6Il8TIlYIGVm4RGGmGFeHUIg85hqJm0/kfWUEFF1PjzJs5yrwRhlmozT9BP
D38iHJpCCs56vLh4HKcb4yhjVyZYPZaLLryvUZHrCIEu3+ZFdElHRq/VJzD6KrCv
SNgYJ+CKlRjHY9w8JiL0fFx0b+QIQoXM+Rfo2T2w8RJleHzO7uwqZGjqeqWgABbB
IR7EXWE712AshHEzVwGYpJaREmfyISgfuUPzzUbmJmyuzDvDM2e36mze5mml1maS
2DrQAzvcaGWvHIMZ9mD5XHtUxayJaqw52cSiNJ/XPWc0GGUnknm7izwnu7tWPQ6t
`protect end_protected
