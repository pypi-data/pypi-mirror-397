`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzUEZmktY2dnA64/pBJlxUQbp7JDeQyVpzbbotWqpXDOh
35SSTmG6hQa6Ysh7V4xIdocdCP7xaxluoZdSmLeqXqNbaE6ZhUdh1l3pixKGOvBF
+aEEkzB/wO0i7YevlmY4v5OQsul3U4JUP61RwjKOR8VjP+HWCDCkVb1t2N5vs8Fv
V79d7qKUGuTsrwGR4WOiKc4nmEsaPdwgAXPmap77FJrZfPucwwJIhWdXOcIbibIq
XXyRTCaCCXvliP2YkfoPu1feuFbr0+zmXdCCfcFWe39Ua1XitzwbM6MUkqYPh7S8
LPNm8CJC+ZZ1R3ZbYtmqoAkIBjpIyZ5onK40Pp3S2l/jaTZ9adibFVpzuWfM4PGE
5iky6chkjQgF2X1/fsQAgXSSE3KHvvFVNLlsE9nFXeGiYccPGg7JOB/hUIUTrg5g
Y+mz26rcOXSmwLtTnTRIE1T+OcfFrL1bx9Dv4Mp3jkNLXD037jFHuvcfLep2G1ke
kvZwrXDxcEb0ZFAZfEIsk5lKuHWqZZs15Ov0YoT20Mu1/fYeAQ+0cb7OK3k/otpA
nQxo/dLAgLfgVXxNa4d6Vj/CwWTpKnQPDBBXjI/GBo13z0yI04eSuQyalS4zUqvN
mDvVHEkXy6OVMr4n9WM7jmU71LTmviI2XelcRy0l8fkg9L298zt+wiFYx1xQ5a7/
t9cQiMSwhUMGIsDlw/FBxBVoSFNKJlZ8pxr6xjtVu2L/336FdDZt/4QtADGBSlJV
Iyp7oAW7Q6kWdz7SAdt/1Evw0bo6xT0oqWtgRxdCoV1uHc/vIy7bvOtYuSiEp5fa
RYxyRcR09++nbJTE4DevLTajnMGhFmaVRDJswkweyy1J51BWP5NI9FN3oyZOlS5e
hsmTHm2TWJk76ZsflqCrYsC4KrX8bm5cB0cd6AIiAMYHRioq5v1Z0XkVhbb8Qk/F
hSRTJ1kzRiOzHtImtdf2cfJjoaONQIX/c2VNaTCo6XzOh+4BQj/KnNc0Iq1sK3uk
dHhlSDdQ3tTdbUycg29DMMQHNIOMC6pvp+0VaBg8VuYIBEYydG+zqxYTCUmhG3TX
R7JNtMzffDqEzJLcdTHscNTvFQIR3loMgr2wCgaCEmYQmm4lptVce3Tw/IwzhXKT
wu9Kk8Ofz3cQ3Co0dg1xr7yvl9rNyRd5F7L3OI/YK6xmdK56i8SgTu55YsjZcst4
rQqfhL7ijz2Wjlg1GliXaiMfzWoFIASy0etOeczNrY1K7OEPFKqvnEJ2oEVVnRFd
YdsfLWNw4FxVPiiFhOvNCm773sa+6losVr15VmJFnm10rtC0/G8XUPk0sb5i1QEA
MPbepDK5EJhK8IHmBilnJyhLxDj+Rkt6m9qJGWIpBdkzMnK7hzVWor4WxHVL5p6S
Evbphx6bvdjBGE2EWkh/QqlVOs5LIq9J2TW2HZo22BUu4XhxkRNkbn8/YCO9lkfU
/QQHs7rt3TDjeH0D/Xslb+fuftMOXYJAzXeDoCF3J5YHoU3pG3EsqH7PXCZt8iV2
J16ykHRomoiyUY1p5K+weaZktyaqKOD0dzRQFgYLtkkdJU0I0csyyLb3lo+3hyPG
zq3lEo+5oJt/3pmYmW6G5+Vj2fURPopb9fSUcU5MvdS+HYPwddRtwq5xRTwfy/Gp
a/bM0Pv+WnRxqtYJXz82FgoHcNQ6QZF3sOFSBqV0knRkjOYLPj6lNnuOpg/hkadb
KnMtp6v7OkspiBMNt4kMrad60UHNUN9uJG1TOZ8nYlpxPZUW01g1hXu1ZVQoJ1sL
6CDSO+fkj7SYHCU0TK6YLKJb+UvmmjTrrDXAD/eBWIiLf5ctWtMK3UPv5IT9DKX5
3RQTX3LTqDo5RlzAoQX70IKTxyeTEMnjv4NPuslYaOC/xSN04HKw9fiEVEwi8Ek5
irz8qLFNtxywSBiG+Vt+4D3rt4j7VHbWY+WA77Oh8if4vxEe6rn1os//4gM4WsvZ
U/FLRALdNreKn/ghE0m6ErjoG0HklN9tkLgYWyXvhlflLPWO6f8otSTpYbwBHPXO
Wu5kdrtkE5ICSGOsfMMn3z8HeXMjInTyycvG/7BPF2YX3oMvoxxSUhIxxHERA1+1
ordhPSU6zjUPF8s4+TiQJJRgBBe7tbfWz0o0M3ESTDa0uHFjIDGJqlG0ICY2NnUK
g6TZ3pWAkjkDiFklJeO1iXibDhGfveNwNSyRNYr0fBKL1ULIqF5p8LzpjgeEw/Qr
TZrse/rezmmO7KOgVi7mrc1yEDSJSwn5weaBh2KbT2w8nWSTzeNQaKAJ8mnoHkab
T4AfayOY5gLaKTem7334Cyn13nJNLWYfRAhNMJ8hQQTUYKOGmfuwJ+NnQzM6ANWN
COqrcFpuvpAWKu7lJtKUvfMaLtNt3pMpdZBLHjRqCoyM45Vlx41vIY7xM7BIHwOz
+a7ZmdWfEWVYAEFB13g6IijPWiaTij8Zy9ohfPJF26Bqgk9tK4jD+XMCu9uIuzTn
UkxdxNfN/aXCN9coYV0jFHsSdXXTWRWnq0bUN5Svtn8s9WKMEiZIY6Lbjr/T8Dw+
74RCLjCNBC43pP/vZwcEjCrPgxyhmM6MVVRorGzinQsGHyjdmVYp1yW6xVRR2T8M
FgUL2l4zp2kUnRvuIytSqbCU/5ZbvIZ7kfLlCZN7MzFlUE1pAia6HKdytzD8lGSa
UnUvEiQZmf87wFvmOnjfM6Xl6DOBePBh+972fyCvJ1/M2dfJJTOb3wGRW75B+vZg
6eoe/M33GXBXLAJYy6HCdwVXyG0Sgo6I5bBUGp9KRQI+vQ6Q8b7T8fbBkp2eJuKb
NtDkqNUJQoKgYWHHqiHDyn0R6RoAOn1EviQNPqsH+D9PpOH8ERUmFc3YNviHBjwJ
POOLk0q046oqtDyP5Ah9B+j3OS1UKpC0FFTWTFdwiyex78mYG77OzvGnhOcAtet2
0c8w2FRGRziF4TpuNwvv33JjiwDCqwCzKLaXefnA6Ev/GCAGar0MTkFF86XeEdf1
AeP/5WkXjhGWgG5npnfUl8jFClY9KC5a+Oqwv48uJAm43Vq0rPSi2a9YL9kD3d+3
NklGRObB+zQN6zdZQoEcXLQLIlLzPNcr7O3RwTZdVdD9LRCoN6qs5oDKUMPbXXRO
IEjZeZI+E2LSXsIBx4ILv5UouIWadAVqiIhbRlx2z4xdtlRTAL+aYxNYRToutqJP
cqme56en5mr2HO715lVmbCFCzK0fWJYLfBNJRSX3KgfhRLNh7PwznKlHvFRdHl0c
1d0wMVPSKH0+zZbCKov2FfIS3qxz6+QeiaCCwGzROuKVVuAxlNbQ0w6J1Dr6uJIg
FjGFxP0pprAhQ/Zq5cwVEVFDM62TnTuyoVoPvok10EWcY8wVZbCBMa7ERjdKLd/b
td9O5YGyvoO6sVxlzEUogpBHP2pNGV1OgGJjCXGUQhyscPfmtRUV/86+e6iW4N2e
xLhPEgwtjBdEEbPochoECdawMuZjiCp3Gn+k/okAzIsynAsWqyt+M9H/XutbPKlV
LGhWknAyf9gN4cyJW+udO+Lt8PoEe4BYf9kulIXmoJ4SeLs/0ExLlgjtXYJZj/Ku
dVHEb4poCVHua5x0k9kQ75sxLqC2Tno80vT/4Emw4rS5F1uJKANMZUrJ+jAbSSC/
RzmS3SkJCc0WV7EkuahPR1/GMgywSsP5kqImEFUQMF3P3YqmYhXAknoivk0sl0Bj
WQCK9/bDaDz9aIezt6FJzYLtejgF2p+r+Tz4ObfBZUXwmlDK802aNgBrwY5a+qln
Kkf6yv96Hu8BhiFtvd+9Nb2VEzuIjIY24fEjnkorInWO0GsVkw4X6bANTPiZwuq7
JaLSOocB+zf/sD19BSW8IYB55RCNBbzh47+7oYo23fK1tOM+ee+lRg2/nTbakL3/
T6JGIhdPt0VKEEc7x1eB/vHtNVnZV9P2ABHBP6WZar577Pc0K69gAkorDrgB2YzI
P85FwqC1wevj2BJp2LguKVtMlk5TjyxUj4vYv8DaO1+37RNWf8XgIw6X0RHwppyL
0dwqwKHrQFu6CygqfM7QLBh56IyGp1tWh1Uce6B51QzMDdIOWCHt6Tf/+s5cPlkS
6MKiMBYXL0PXIvONBo0S+56fj/+4069YFB0240lum4Xt+/BaS71nc+kT4vFDipJG
1S/81ZH4Aa3cFjXbb8TpNXNC40ZUYcYlQJSCSOu1ySIDD9zTitWixDbQbG0D5BIv
ZgCPPZAmiOobruQKCyoYT1dMVMZIuQN0l56JF5s3fmBd/vY+rnBCCV7ayWl5q4SY
qWQMzyR10yVHXQZpn1mBFw==
`protect end_protected