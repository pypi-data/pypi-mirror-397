`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOHwrkQXtZIk/inau7ZD5OPd8/Xj+D+7urt2f8TgWXvYNN
2Ko20oMuUv0YZpLbEqyJlpULVa6ov1jUeiQw5WEjKG5vrRQrRJvt0FlOZH4PSe0A
RyOrZOvjFFnFapJEfMS3f8vhpFlEL53wicKbN8O6gx8WqRAmC/Nk8UkrFB6q90KM
2TuoynEeHHsXOTDvXA2DIGpgC/RAIy6C2cwAPheN96ADw83yeVlElfhhzMTSven/
esvP/8uwf1HcfYOPV8aCeEuh+8iu6jUkk6WBWTWaEtnIBPfGujJPxPV+hQPqKrgV
cFEfEbvI5wz+UjKvzJqqt3wtV3S8K7zxDsmdXLMbTYktZ4VLk2DdEl9fb/Ex9aVX
DMus6YE1h3zx0p4r3LiLU6fSw63Ra8RGNiMA2HSqJ5Yg8VUOLMMJolrKwaBuT6me
7Ci9mk0qKqjOpAs/H+gZ+scY4ekmsFgddQEy9UhC+fco49EpAZuKNXQG3yBfG058
mkaT8a5sBhWFLL4+rPXZlRW/NjsRprxWnOsP7K1Evpfa7Ijfv5o88TxgZg0/c9Fq
T5LwUArx43HaYuGvTQvZB0X/1B1E9rLoU6hk6k+2bTM2Vt6lhchAVGS/XnAw1L7A
YRggpkhnZhzR2okMETPFTgXU2IgKENS5Fv/O5NWlvtt9xJYRE+hyYYMsz+my0xCI
NuZuaoXi0yJ2Wv+H7aCNchwqtf0GmioWzte/FZy/+Vj6G/d8DU7dHBW3gMDZGjF2
aEv+VSQA3EwEwYt5F1LWrPqEHrd58pvk7CyLkwgedlOd22DgSlOSJLN7qevxoCSw
xKVpFdFsRxAH94v0L5N33EH7YlicqITSACzKeoRWlU4VAbTmYRC1Z5SjmCpGGMx8
S6tmhfnjiRfjbMXEYaTM+BMqn0N4xAYLpu+hSHBkz08VZf7xYAtDJ467MgEirIuK
mFBVKYK7R+QZTnjP2ZKXgq0FulECsG5mYzkO5mhEgEMomauQmUPHOo2FXGJ7vwOb
Xm0kbNWyUuhmW4KAJY7Bc8jb1yL9TtzkbAkojtExY6dvKfHQOdLbnsbPLzE+Dgx5
GMdNhki929J8DnONq5/bHAxr0C08lJqco5iL5OORVKrGcvp0BhrrbI10ybZVWHcc
WQ9LhuTM05NsOEhpyg6Jwd1fvniOnwEc0Uc9q57gXl9PZZBuGarydBCsirGqUZ2O
meW68gxuq56zZRR9SOmKZrTaUcur1/tZdZzVo2uzS48utkteCa9Np+6NRloMx4bD
H2NMrCMzr6MYgFcWFFnh5Ylggvco8Zm1QmgmAEqkaprsHCNaTN1OKf9G+fAhVqGr
W0R94LeSerOWqkqLCvQTBjL3AYfrWX3EiiNzVcWFeZaSjb9qQ5qXvSZS+odWIcbp
DsT2wR4/iX5LCUiQZHhzGO7QVpIzR4MmY2V5Ql3+4cFYDnQBvmkC6fL8sSOPZJ3S
ebgk9epo3pO+3zEY3t4t+gWhN4erEZm74j+9YkiXDx0+FNK1g5348gx3GPXxCewS
0cTU/6+tgK/ybRippw5fKy9m7I5bBAhVd0JMb7TpN54YuHoXYFoCkCPh13WZh3qQ
C2mgzXmmNNz4tvYKSpoLUGDrQ/a2IZbW3+iltZ9BE13YxmbXGgZtA6m6HBy5u5TR
Zn76NUX6hHrvYsKsS0oHNHR88Mi8//BW221JiwIzoepq5IfX+FCvYTHXjAbXDa4t
c5eEsUqwGnSriarKB4pwoew0ErSsS9bQv6EBf8z+LlMH1wb5G5gSTynZx9pQ/DVQ
5UpEcx+MGvTRkVsSoLl4AFBLI3Eukto4X4CKNX5aV5QMWJ7XDYrhQ5kDXrMTe1Yq
pvOBYeXrpZY2381JDvr19L29VK+xCMtc9p/KM1QFemyzu5C21+2CXh7Eg/2Tlsiv
NTpSD/6WNrOspkC9lv9ScZp7kifmVZcwXvvmzq5cMEn+0XwHkTjqW+Pe8r3l736g
UmV5O9JaLlNyhU/AfiO5Z2FryS3Kd4WbElWO0mXOeKpBrJwIXzAdAgQbwyxAUrSi
qTaqdKEZ4AoPhXzHIk2wurvEXuj2DJ7I3i4s1RyaMQga7xsWFhyYqBej2LxXb7pQ
LoR0zqaWMcJcoDXHep0bI5I5yUocxgQ/pYhzlIsZVbftIcAIPUa+3MuiwpLNpy8i
dB2kMT1af/q7mMqqwbzBPw5YdPFHjeOUP2F1/adagkJyaDu2Xn5M9YcoHuPMKfIi
8wp2HWemC0OhjHsJQoAlDX2ra5BaTO0v8G9EnjC7vMGd6A/vZamDakA98lN12cg3
mitwjkvnSAraPA1t9FJnfdCW6A+n9Hri3/kededsjPkpzCVnfaujvXf6eSHVRWQa
oy2FTmV6fXD/tDadWecSbGjPEDvm7YkKXzTZmyBfqWIiaxiJoi+CIGzb9bwt1Q9X
j+ee1NHTq2gJuMsIf/Js/wKASYsWH2HA4hpBsOaCnYEsKVlmMZTZZN8PHEBHinQ6
c81ofJMnzRtKeyY+oEYqRmDV1v14FJkD2Zu7wsr4GYJuRcEqjJEQ6RE7Nr6f2+6/
G3R1XT0sevnevC72AVxu0GFviiITaWGCcyCyq8b9S8A6FyelTQOdw09Ci2/LuYDl
5c5VdEpjtd+ag5fZSw3th3BX9KnUN8Yb/hS1+9TsM2wMUQ9XyEjqxnm2OZqZB5TS
CM0ypUn8bb1Yr67j8YUGsJdk906pualIoPZX8my4lUPKx7R2qH7JdKRIP5RWhDvf
ZAt3UxzwGTD9IwIDZwlMr2eAk4ais3eiWZQpx2YKrbw/HC08i0/g58DQqc9HgEZb
kolovbzQDoM0f2mEnHY+NMGHy3AT72d9sR9ep3N3fNShOp3LHs6rcV7WOGRUWLHC
O5PySvnTSsK3d9h4iGdTt7jfMOYZ7xWEu+c2eAYA+ByNEu3HDUHwHNN+20vK/i91
9NYf4yB4UzN5vGtlZzfSAw0WgtfCmqHdxngeTJ6UCLfi0zlLYzEHmUOB62jkOUbx
DzkZq+YdTXkSLpJjNgCtUZL6G4GMCXi3EZD8ZCpt7Mm8sGTWTxmPzzo3uCfwb4m3
wUHsLPFFY2yRzPld+Qe470tv8MQxaa/EZFJSHJ4YoGxeAESTXIUREDa6PpRvGkwS
1xwix3edd5JK1wd98LWXH3OEgPOu5YOTgDierdgFifiT6kJi81aMvkEsCLDKetaa
P8R0PcrWUhtXv0ayMhQAB0wjc9t4XPz/Fm7+mUwAZEMzHnJSm6R+yoLbbZBpC7gv
uPOATWPPdL5RDLx2UsQ99mVi9Dj3B0QM5TEW7AZ4UdU6FPZtmo1bFq18ZPjou3to
AMCaQ4FnEZXbXq9OjHnBs3JpdVSoAPTIto2B4Wqy4+7NnXytogI7EKAIDw4Sz5g0
NoC8Vn2uT1ovrkT1WeC3O0da2DWSmaGMF/jYo3MGgXRFtodHFoJt5Eo/7Bj23FEw
bFt+8Md4D6nslqNkOPkWo2yi/B+1k09PiF4+YsNO816J+DaroyW0VU+z4NVn3fnD
76l0f0P8F6/HDIzI9fiNxhaIu/YLFh4qrFz4PVGzRyhr1Z3s3Wtc1brSTouL97xl
1OJphLHqlurfiOWZ/My2dY6PKHMkBHxCv4ekCwUrl0Dd+u8y7ldZM+hAQ8WqM7f6
TeLRnyugLseEA+LD8FislSAf1E10rBQb0UN2MHvizeFPLOse4056EKgx2dj5jwvf
atTLrRt65pECSp1vF1AHJ/um7plQxbRbG2DcHGOaHgLeoCW8IJoz+GaA/TjotaIh
LqNZ1PV1j4ttv1xB3wrtVfongx6f9ptO0VvYkl75keY6eQtYwFZM7yfUsDy4BDSu
cZaQZ9Vb/+24DVRTi+DfVaRTkMjH3RdiKLjkoSP+fwf0TQbsDnROPOccUYciHlzL
nd5oZ/gzg1ZY8ByfKJ6eJ0QOsDOvKY6mHqM+w9udWXbwk/9OR42/j/IzLBZzKGZn
LBghTFgc6QN05X29c1fR0z2yeNpNvTe3e3Y6bplLmbV+2xd6MnEAQ0XphI7CTyaC
XRfenFrUbp5hnd7QZ65lBIQyOC3dUwSzcPL07veCEA4fObt3bI2He88LdMj/w5EQ
/lc5jrbBp5lBmqkf1nvXRZtt8Ar4Zip1p/vSEBEImFBMnXYDNGPbLvP0v5luUMKJ
63OlEHflo5Qab3Z/7Smg9hLVbsZjU+kmjCpIL/BB6b/bJbJ/yB9CBXZ+AO0Nkwbm
4/FMSRKddC2WHtiMhPok20DzuqtRdezbYCXcnPA0y0F+PL9RwixhJFoSmVXkYYve
ELuVz8nYYDqtSqIVpSepWDR7QrthaGG9uXKRfH3YCB4mFcbmn9tlcU2l/WLm9nKT
HL40wBM8++4IOelPdoDPa/IjTRKbLlTmMN++N7zVILLauYxHiZNZ7PzVDlaVrcUa
p9mgja8xoK3KS8sbjoUqfKQqKKm3JMjR/axxw9Gs05e5saKzm0UuZD2/n1XqkKMz
YOo7QsHn4/iUaxeZi2L5LwEbptv2SXEYfwEauP2+TRZLSXYkjcXh/zE334DxbeIv
MgbzItuxSCh7a/lm4qm18PO2l330xs4/sNC/PjhwhdZ7978crmGsM+K0UcPU71Sj
mj1SD5RyDYWhv8AIU404fJ3i+T1Agbyww+xL6EERXt0lLL5nz8MnvqYriHvDRw0E
ZeBI8N8Ftya5GzTwQqNcKmU64O/2J1f7IFW5fKnGa+a/0BIovFsUUt3j4rDLNRKw
uHh4P1PiA4RCmkcSQsst+u2xO3JibGkSj8YLhTJ7CWMyjwJ4PjqJkWqU88KNtdnN
BUiAzH/nCXDJu2yojA/h6Ib3T/OpJ+PZJ/gLc8MUFY5rCy02bmFJ4gWozvXUIqto
eYr4c4mjlYsd/OrtgbOLblNeEAf8K23sKkHjBeCl3gUcXo3Frp/cvlvRuximuFg0
L7KHhJm6VUoIPJ2W6Pw8gyDY2740/lTDhDbIzBbS0uo+3q51jc2Gil4hgCHzQ1UI
8/UPjpAhr0q+XnA4zzFOPtoAUhxM2CSMgJVtD3t86GBWrNh9qHs0KDhkU4isWhjk
yGBURJUtqhbousI1Iei7YHDE+wUFfsiEzS+R/pjxQ2KsC/FRX3Vwmm99jN+i/mI4
EGdnLYYMrLG3hxO+37FUZTRO7jtrtPsCa7V64gn2k1+zRS2gOaJfeD15nc3xJ2p+
kE/M7yo7BrH9rOZ6lo+0BXpJPQQjEOIVtKMICpSafm4VSaGdZZfdIPZh+adXqnnS
F7i1TslNfV0EMkXE3jtBbp8ekItxjFFWpn5zG+gCC8Fd4FHHxTQRdyyyZyRS9uCx
y5ttaY9CxBElAQWjTkMyh+eSoaQVFeMbPuK4NnXBiPAZhUj+oPvUgKGNT81DrGEB
aJE5XPa1LiymFSVKRqCOYaTE0VdjfZrDfrTqLy6Zygq6NAEbtgj9xigzZXYNoSL6
r2qdBs9knF4oVLwywrP4M9cTTTHKVu4A2xHprQ4iDLsfLkwPTHtp7v+uW+Rb1O3R
uUeOLteXS9C5WixlAXmsTMItpOKfWK3n/lD2tJYXLVQK4aT+4FKENEbtOygN1aEz
HS7uoGeVd6m8ADn2Whfv7AK4p0Bu4iXhBRCWOrXTKeE6HHnm3ecOsGek5JtwKpbr
fDXWkzE9QT221G/eHTvGRIQ4DAWRclCBCRlSYUWfjcs2i8EDcCW8uW45lXNlwcgo
YWX8HoH0DywLTohzgYboi2p6GSZKAdH2n/iCwDSZShf63AO7XCFm3Yd87d4dSClQ
Fv7rmzGdA0vU8FBFbB3E6GJVz/98xKVlLj2PrMRpp4SrdO8hBPQuWfdQxbzXYCRb
mtw2j5aDbQN/ija8nVqXOQZybwQenWgB6zRh6qexlWWLKl0K0rV9iGevRfoMNI6j
AJ/1E94gG6e8HTmNg6ef7ikuZxonF75/dluoUQHkjv3UvANLYqmHNEy/jFVQULDO
o4tZayr/v4BPGqWvnmVafH7wpqwYupwM4Y1rKYlq/3AF0PKkzTjOgcMM1gVWuKP+
IMv9AdMXJEkpujUedYZ45uz4JbwqX7LY4muyfGWtrY8ndE3D9TF6SDXl7lr59rAI
WcYoi0UMZmOdDs8nI/LlDHl6kMJNo2s3ZAR+Ns8ofWmdTS3Mje6bQRoipQiRg1OQ
TpJv9Gst/tjbmL8WQqznhENu7d73mM/qf3i6d4iua5h0Ar1ABXAZKTEyNXMxaM6T
XxEObGI3zNsfnxAY1/U3vSSOr68UsbkevB676fnjpQ69RD6VZi9FW06CRDpvKowB
7LzUZs1j9NnDPF3KqV94BwawGG0raJ/gU6oH7noOTkP7DNgS56wYLW9pY41idHC0
YdSVI11kSddDFSzS1oYXcgAyc6T125AS0q3AoMfY/nqT1F6Jwxy9G0E3APUJtHuD
s2kvIxv297r9u3haJzv3PayCyPwc7KMVAgfhWQ2TXf7WDd0LMoAAuTHl7P1/Ng59
DKPuVIWxj3KzZ+dbCMOPlCftpt5q1ubKRQ4u5wwI2pMKuy33kZDi6LNwggPcFuQg
gqleuJn3Pwcl931IHupiKtlAvZIDC+5Ro1d69ska8ngtBYtARwddw4BhcrjbMv4+
5/UAyYhswcawFBIfsOX79JyU2Jd8eg2r7t/Z74WpylZOoyZmA6KlCIUkPH3Mbam3
jq0h6XthFj3R3MoTXH2XFxWgIu/HrW13Q4r32Wxydc24dbVHdHsy4qlGbMfwT9E7
lT/hJDfntq/LHLYIVSEO78JM6WSVzNcBWhdH0/2D2QZp+hRldbYFp8U42gucj+Fp
Hbb7NAAEq12UTwZ7cSiSl5jbhrOrFi2Ox5nNw8oQZIzT54NpAIHddKBk8Sxh+aPU
10bxqtvtj/jnbMVOoAGfvmWMEajgCiJlwaLT9haTvlfTjthZCfSZ7bP47EjJQL6a
BozRrlNM/HamAfT3t/mI2EhfXPQ4nVoBWLNcxleph3liNfN3kFgk3QoQk4mZasR2
R7U5Gn2cVcxxVRvTUKUl+WXordb/Y80rYSD8hF//02Pe55Nvfv7bpmPQ1YEXObEN
MMTZToQktPOjV/ev9BRGa7PW4KOYSzmfT5LZNoCSHWMqhuhChrXS6nPDbrPZbl/E
7BK0q34fdu5jbzZQfqa1yNIUmmcI2G6ptVD0c35QgMlDfaJimz+GcLT9W2Iz3pcl
OMahBKKb680hXDrnuiqmYHcj+34G1ZkS0+RWvTTFlRlKcncuepOWbXty8kLd6AjK
zPD3ScmhgfHbRP6FN8g6v0JzPWV/zs0V3SIkGqe17FSzMZ4gE3KtWCyPc+quIzMy
WBMpfBt/rPAeu43OBl8AllfJonZ5Pm3TAykhqXWsHEIN0qrhpmRqaRby2cRBqfYb
op4lN4px5IZwcUSlNRVw9kE98txKjHDcBJjHYmTx+cW1AI6vl02dx8PZiygHlxUO
xU+oZro0HM9ddjfMbn2BXjX6ZnUHbHv6dX/NVpqd2MgII00jkhlIcHwb8M8+LDap
S6IZEGJJtWJVG2pac+IXEKFbdUe70PgZ6UNSDLa6erWFWi4tJzXG5+5hTqEpO7e8
bJyfiuBrIUyhTC+3OomRqr7UqBEU7iiFcbw21r0mX3Rbh7emTt3YGxyVQI50zEQF
EdTfjWot1ZVtt0M3rBWa6M02FMVWxJ3dTjbBsuMuoRLIZUI7mM140GX+vkm6nT2E
V36FXe9705blfbx3XkdqdI8U8IkHS06iTZcFx8IE4lm3a+eW9QHWtPJwphnACF71
p88FDqAKMrWvrqCnWRiaCiaqfpgADmXYM7PtOcQrJGHI7fFXOKd1Avgtgx7ihS8/
0pLaYee5fofhtjuXDlOuvGwCGQAEzmiLmVX8xPeO1ZAo1NhCmlK2JJw+OvplQK+M
pMxMjZQF5q/iZSrnxClYL4yINehtCoNrGkWMm+DRxElSCVD80BGTnMUvPzQ5uE/C
X31YIpsRIVscLY6fKInQjh4iM1xkvj/9WrnpPqcvkH0xIVgp9+SSsgjCFyaIR8pm
p9TKYTW12POuN3B4pSrAAyP+KR1HhTHqqFsz+m5FZj94r4WHg1w8TCibD84ipFys
NUjf2n8Y4XPVy4oCl5Ba2VWTvDjZRTxHDt/tGmAP/5pkpQrm7y1A9d2+hHsaj5Dm
N5rVUOTOVa+WOulMUcFyk22lYtRqIyv/Kqdc5GZPKgo/p0ftem9lJ+IPn5QdyhGR
tTN4CiXBl0sy/0UpB3NZzzZ++oP12r1E9PUsp3YcDc/Yd6aJhlaluUMNgX4ViQlF
ygfFubF9zhbz+0q//vj3xhcjvM3hFYOG7xrKAJ4w+oom+qEQAUkGF+QtzSHkot12
lyyJyIj9blSLWWgPgJ4+3s2+taILKwo+Y0zfFx7/+8T3xwrFELkVuEWbxyr7NwDn
f6zr/iQL683/TDkxsTgfyOWRSzwerWI0ANimxczSsfpcj5r69+nbKGCgS33xEiiT
lNs71JMeci6CcI7OM5uCURvAALQzLsQBoA4Wwo725/5CgsK3B11tKiA8KztEICLY
2hzErzmRRlfMzXdb/QxsxT1oNnj65LLH2cFAHDpbSPVDwtKDJL+XVlmlqq+dvTsB
K5u7yCd21fWWYMJLgFUC/bsQD0lmHUyeUm5PQpGdhVF8UGToOUXloXvmJvWN2e0t
GsWLDyIfoXQBevCOMSIdTTPWakC1c8zPlL5nN8dY3nzhhX2rYHX364xZhucCdK/U
9/+b/LqgD48mHI1AexLJRncy1zxBX9JZZYFthwbJ26UEHomp5CjSSAIs4w2EA6BZ
R9EOYTK1/jVhOP2XYmiAKFkGv10SWumfV3ILYmBDLHbqb0Jf/xbsjlj0EKNCfD8h
FqXx/H7Uw1TNhqRxSlH64ep2gTc6R7bCaTiqO0Iu+H1h0C3pNe88XHsyaxgYYT/r
ftFrsQAK4QJT0h/TOD1J8F/UO3xOrOmDB+Msr4YBjxib+/D6Kgo6FDZgf/h/iobV
LVsCXgm9lO4EIa8etFmg91MyzKMHOkSjjNLYpIDQfZwG+BWGayX/+X/sK26SOSxH
0UJIKgdEgUtbm2Bqdmxl0drNlftECZdU5YOR3Nr6j7LC5WQuza/OdtlbgOVSNPxo
KQosRp7+uGDR/Up7jAsXgF/9JTrySHVmZegRk5HgEDS4r29LQrriwggPn8CFKbrl
TryLsxzAyQdxx3adPnRDPbRjtfu3cl63MsyHjFT6cd8IEDxnupb7ulQQmTb5fqoq
KzIx5Iy0Ox4iNIihPVGX71Ulc/YV1BCD9PXnR4ov2mf6kaDuDpQiZklc0PccKx6M
hW6hXLd0e4Qxfm8oFqkFQ0NMUp6hlLV2/gpj1JvmCTFYMn1R4dOvBw4Lo3zPIGB7
aGo/lCIdXHqhLYhPWjRzDQsM3KbnNLkIfOW1nsRrEiNpIeUcW3T3aLzk6gxESL5/
VLoWXWiginGY/ps98YlRVx9r3N0DeqSaAJFk8gmnCYBPj0iJYpQrnaotE1knMoH2
b492X+xs3OqkoFkZUpS06qcIS8A0IaIEJqraARG6SXitt9reKWhxg4ugv/PFi3g3
bz21j9C9f7RHyYjPrFeUmQJPAQKXTHImYZ5IQYADCzC+Phjx9W9RRc1cMfjf09Xw
rm7OEJHZmY/Re3Ui026wF+0BSTNOeJ5gD2ioeu+ITSr0ZlxaEXOq8rg9G3wgr/fz
pi4Mdt8SMx81yfRPY7/j5mBSIk0V6QdIGZjLJtJOkQNjKqfNyv5RsEx03ia5zT72
fyOl8mNi/Z1M+7Z2/CpOzlYWGY0yCLggLsakx2nD3LBb6xrRdrGq6HA7cZYORH8+
aup20rEKplALiIeKy0ffuUn5wiO1iofTUBLjujr97qt4+LqlWHebuqqsl40S9dje
JJGZnjKkh+gPHiVe9l06A+AqyLQPcW38LjZwwXdqjczMsnKFo21smBe7LZmlqVkY
OwukbXn2uQqETFzbt2Kbr/evAgvHwaJBm7RugTaoiTT6+vHhxt17ctYUkCsB83D/
IRqT1rzIwRkv+BKH4CnlbxkReXj0x7dvqHZFrirU7sw+Vcy4NDEKejvZ6IS82AwK
YQiZWEWX2tgvCewRgju9Hc7cIURR8z+Yu66xkgqEud4BWMndOL2w51uGpYGArgVM
brkAVlEQe6xWM/tTgOE1Dx3/xWCmmYVN9qpCkLqjWxAbXX6GV2oIR6l8bX5jQNvf
/kcjUdgGMLMUD7kKALK6vnJ+PyjszhqMLcVnUR6NBcC8eWT4MrkGiD4ultsB+DE6
rVV4ddxJB+xQq2HH+Bq+K82lvKl33PjWx+jhz3zn7IICu/lKe6shgMiEx8JO5Pbk
PtGtbqilga24GUoRMcSlYtIYnYqiqAHxwb0hlvbpHO9KSHaXy8xs66Pm99BOYp7y
FyK7LTMLhr8TokQv8rXpL1yn+/Igd5ER5C1Cgu6v4vQeaPtK7HujkSNNS1TFxuc1
hmNNZFl6DboTRCGZdEHovTZxAymUqhMysFy0UgWtLy2vpKSTHxACGgwIHe/ckq+D
iYXLkDkYRgkh9Uoz1PCq4NKHn3Gvtq/Mv9m9r3n0lZgl1LC8M0viM3+jM8PFOrG5
YwItibiBUZBL8zdDLMgFieUJDVOAHN8UiBXe/pHQfto297hcRqXfEjO8yQGH/69B
BDH9Gjn3XENJEfdjuPIEJsAlmQrFqYLUO+BX3157CbXYmFpNR8KcudcxN5Cijz0J
uVF5lM9ITBReWYJ/rNu+H18nUSc4xRy92W7Yajakm0pELYATT0ZHT4qYk45Ft+Gx
JKwBWjU4IT4WaqTpN+MTUhPUr9Xx8gqWA44Bvi6qP7/h3cgymS+xSQpdYFQj1vz0
jOHvGkpozsv35YHL2fUx827DyZ9UpmCN1lpllC84SZGfRpZRg4iD67uC8YMb4UTl
FLJ6UgIPu9o765UEgi4QX9M0/RA3p9sGfDRcjMRfD6j2NskgkFL21UQ+hCeJtUgR
ExwGFMSvrszP8TXI/LiMSRa8FudKv4Ozd4P07mtuduBKFcn63/T6j7IfR45i1RKj
z+fqQ+GOLsplC/+3cQCG2gxkjDSHEby55jcoPt12Qd7kswDKWqA0nT5Jrmq/K61n
L7c2XNbODerzl0rjqdg/jmf24oLEQjmyAkHVILI39dj2jUbcstp8jSSu+5zp+e7x
xGxyx6mZsFdfPfzIbszVU/HRQat/RxypW6sHAxJcSqK7PNt3PHQK8Tb+Cvr6GCYf
/s6UEg8itouh+XJX5m8EOCzOHHK1ozK/OgZfkGttr8DadARAOG55xzdBp7Bl5G0l
jXIjsOb96Rzr3wQjketZfTdn5yEvoCAG6VJjuzh3fLWXyYHSEoMWA/fYJw+hcVnl
u/QLX9LEhdz44KLIH27vfYHv2anIWnTpYH65o8AbtO6VmUjYyBBbt2W+LrYhfoGQ
rlQWF82SvoeR21wVG+QI7/LlASUyHzRapENj0U4qO29l7lj/HcDoZbUlDgHfEStK
7OyPwb3tH7TuO63P43hMvxW20gENTpUeR8d2W/uHHw5OM9kqEBOaUa3LkaW1ZBl9
MM/UWVq4GaQX4E890RBiUqaJ5URuuThPdL9YQlng91IuQCwgemgFJvnGoju0a+04
FGqeBjAaltwTRDJFx3a3NiAUrHl+5EqeV8D+0XYkWX68DmW0zT3HWE0V7eM05Zuf
nRBW5jxm8mC4t/QVncgq3CDvKMmD33WLM5hFX1VMXPP7sIllKF4wVKI5sVqUsv0o
TCsd2kpLxlyfrqeOVtYdN9oCbvGMIOSa2uwRgEhkDfHaqYePCsx9Ck2DOV8hF/cf
x30vO9ihEOk1ED2zn/wqcuCyOPiBUShBd4vUx0PTYR+094dEbWmA4Wn69wxM1FCl
INd2uciWVg9/PjJGQfS7v6a17M/v+zsVOe+OoTF+mJoEiW0Piq4O/HtvSQ8wEzxc
EqdP0ytgYm8bf2ro2kwEHwPBBvRdotDC1GyCxKzZuY3IFyBzjfZHo73gKErPrCBL
YRhEInUa67MrakX+hsirzspasgUFkKctyj0tkJrgvE8/dnr7qymF2Jp50iHHBhiV
VEdCEXg6uIsnolqNY1/aGGf3EMezxOorsz7mizwRQVkIKdkT6vSH7wMayHxQMowp
JzEzYKTGJ9Tk2fpbqWyJAa96KcyVSgBNP9Oo2YTDXBHj8lLvcbG4LXPIMRCGZFhp
kW78Tr7D5MgPhB9TjBLRtkS9uu37BBKiN5Hw3g0ZweQocRDffN9aTijrXvsQkWeB
zpE33KyGzkXzzRIDJwTY7Hf1iTOapxNSMGVSq9h6PUbxUW5dlaioJZcm8nv2RPfx
i9kq++gLrWV01HpNVN+8SoOFDKFaFBt4HMhubKoLDmAbUvqEoghk7kqp2213B1rw
4wQzWYrrocl42tF9/QfjlNRJhLZyzHKcDoe8a5P/Cc8HPZHAlMHfCHsGkrRDGgVc
iBoyO3gyYEOGu+ZXC2jUPIqVk3/BM3rRVV+ntHuAfTLpDPigl8F8iYCfdLtboUuq
i09KokBGX8+2jo9a4XFuEEqHxWBGfut/lEvo83EK8nTA7V6MxfjQyVg9mDe1gxph
wTTL5EwQFinVMPqdSLkjsPTUEFyIaow6kgZlhdqHBjy3+egVZTGk8haM6v7W8ntV
qkVpJbEEVczzU+udfjjQHCvDzR8Lr4+CsrfP8f6Ldyr1wMpHp/nqENJirH39FeBZ
DEqt3+7tYFtP3btPAlMYGuYeDsCpIOvIsDt1KBBuU+rKtg0f0bU4wNF7JMC1cUnB
RTXHKVcii95EcoAO9FCoRCyknLzkJ+gmiJjIrZP3gnkpbEavDn6AYvAOzvUpAc3R
h9wdeDJQYIcaXF2twZhKKvCejAUQMYjLFyGevu0gLkcSvSJ6weBl1vY6E8sfhmjs
HpDMFWi4VTRLi3muxmVoi/sNHT8VorNb/MXTQvJZfXl6a3AmOTNNPX9RdgPBPvJS
MU/2jnpBjmNTYEgd2ciK5E2k0m+k4oSZYOUoFNBXW/Hmupd67HPGuyQsQ36nZ7x4
dcULlGoK477wH9n1Kq20aJ7rFelcLINoBESE4cNF78rtQjiEFJhS+cwDuxlFNWOT
zXx8JMYyLj0ghcPZfW8ry/2CCNbLWYXSYao8bvh/sAMl1jwzw8oqxaPvoXpZ/nzf
Hptp9HOMhjop7EuRTBe+lYWP6L4AbhylgMku+LzVoA6foQg+IZs9w+kZqXnlmZn+
Lwi5Dws3yEEBWIlGDiEGHvkHZrrLZrrv8Nu4rBxdzEkt2WfIrz8QxXzEZgzbMM04
/DY2bQVOd6B5WQMX3fN3OJKSjrje37eQvvT4M1Y7JRyzGwqZ6E5pHEslWDwmsDnF
B+QNlwJZ+reW3NCiNfQjQvNb06PXmPuYPPLmoACEm9r8sByOBO3hB4ZeC8L12/oM
EVc+SOqCryxvMwEcpBr/E0D0XfWjvuWT9ZNYwqiQD3SO9YRXM6IcmLJ6WJFt9Y+Y
A9PXForXqtJxdNfiZ8aTrvSDktigHvAFxGhOIpuahqSU633+6AzwvhCIv1p6m1QL
28t2vk+HPuk/h33MYhNDPY7DknUxlQURSO4WagCf5FIGTqgGuuLv05hgWxeX37Uw
ITkR+O7ZFcD/YtDX5jmI3aZ+s+gyxfpmLZVxiYvWRvSRkrJnHukeNENO+Cm4p2uE
vvwiLxkhqaCKavoB9hXc1e2e1mVmmXVI/5jepWwqSIv0dh2H7ZOyRg7VN9r7IP74
LEOZMOYFS3tMoKlNmoFNjY1COt7NQ90M9FQ5KJAwsEDCRvL/mSIcYqWrcTFDhdCq
638eNczuf7Z6kPNodSGtstD0TEMIPr5JqEoJeKS9oVHreVqIuK6unRYe5lKP4VoQ
ZuKjdKX8h7IiQAxtrLKsarQ7qEg6w+CE2WZyyyccQ/lR8rNnGL2VUeGOZJovvfuN
xTDlBDrCkIg7ag0aWrJHV8KSMXdYTpH5dw62Ap/g8tYnrlfBnlxGrKvRFBe9e7xr
tWW1zXKClH1GNGT8fCReOajoIbK0qVqLkHQtuRzvGqZ8gBZ7GvJnQ4aPLPI0uUFV
3+KtwHzWlj3XfyBekjPvVD6qsLgskBgmkG3FyinBMtnEhR2B1zk7BFFGX+VW3i1S
LknQDDElPx2/VQu93BqPWIvGjj0s3QEG9qsz4kk6mhwuJRe9TYmW7N9VPZydjSXl
U+Gh9z63MjnFaBSjCYBiI/v6vIYICwwSb8Az0/H7stkS5k1gCK4txtq4chmxw2/I
/IOhjwwsM7Pdm9BmDngjD4IARt6dF6H6fTfO0v+qWbFEEXFCXQNEf9IdCOIIhqzM
eO6xsfeLU80MAF669/XDzkGtI0H96FVklqFc8eo9/2UvUD2xdtCGetznPRQz0EA1
D/cZRK1kzMKUUFBPuwY4SJzOi5x78q55Iy78XNl3OJSbPA2lFtzCYp3eLQ+XddE2
eEECXRa1dix7MEM4f/MXL50Zfno+mCr0iXjJI9Ah1bDDg7DW8R93vZTY9bUFg/PW
3TYjVQnELoI636pPekaDNi9a7ZxIKxn41CTsURWQNFpAklyO335eJADPR1CWOTvs
s7/MHVIC+wQUZsjIpEhMLs8yBHAVv8aBVlaOZ2HfQBdmJdick/BQQFwXGCWe7PTA
FN4J5yTHQU5hlibfJ7qGCmR0D50iAfCSpZssluAqlPxILMeEjCgff+ue2ycUsxjh
G528xkJhcxE4e3lT8Yx5UnyVn97kiGotAEm7JzbhL87wUsjvG6ygQ47dKeHozNrM
h+SODYKDW4VRMpon1nD6HsLGFgxJXwIv3Zkur/uOLzgKcZzZ6X5uNdOx/PaUt7VS
mIRga30BO2oCFOmjcg00usx+MPjV9N8jrmK0yqEqBJtC8mVQ+18OdFbXUW4Wbxp+
w8zJU7ACTH4sczCw6WKcDRIH9Bjb2cczaE9y1gvR1t6i+zMOGb2nZEH0v/m/1esP
KMUm4Nz4X5d4cVpejLX145pXSZZuBpcZwrRWXEljf3vqpgomWXRp7Jaq2wL9O5Ix
MYIIyUlLzUH8zNcGQq9ftVG9+VCB1uvMJlADFUwixZFSCxYfqNRV7OBNk53ft0Ez
ZLC8grjXjM2mu8WAGNz4EkLZTuRxL1wMZmpn+ubZDu/qpL7jO85PpYi/XPlvjekU
nsFozhAWaLNyeOXkzio67eh/+6Wzk+TmnmZDdC0OFIC+RBMvxSbRB6vSpIkKySm/
8tW5wikCsPGJJAwWKeN4yFScheEh0IefccZi2VZ0LIZNLk8AJ310LW7OiwfByLdo
eT7zf06XnJtWrw/9u0Ya25n5q5hKdIHAtXJsL+ifLdpgRfQe+1/hwM1iv8RNokDf
5VSpUuJ6Lk6WUkbO+zNyG1t7lQdsGljC4xGui6YBIHpbOBg+xN3QEaKYNuEwMPoB
bjwXnfuETg9sEYUc4Jt5rgWPPudn6xoYMRK+ZKFu+af253YjCcMC8//gxvQo4/Mm
cinZ6lhnTtqDxkVO8n7B2g5yDv/xCrutryB1FG42NKByxGUmL2rlKr1ZgT5J+9Ru
dhpzTCxsnRta/QimCNjry0l4vXaveemFB1F74tniVPRVeJwGtvOIOmzexl9SiN7b
Zed48BK6uLrUkJWZWKRUCegQoNfM0BWDuZR5TSzXbJvgdisHBVMcIkW7blLazv2j
lNzVBSoyfkSy4oGTfuKtFnzagAT82GuBWJaG47WSn7WMULLjGq0vvlDbdfugLbv4
3vvuz9f9IrJPs5irBH4Ac+sKHKaQ/DBXmijoUITuYuYQzn33rxf1uAyAQndEsclM
y5bf1qKWqgeRprP1f6mBKA6Iv1N5J11xnf0RYPDa48Rh0KsnaiGs8wyPvMPJ2zGT
RXiwG0KRHoILOBozVncg2edD+AsyCdCm9ThI2kFTVhQPyGrNzdU9tGy3SQAhGtzD
gnRnfNoAf9/Bkkr5+qXcWVWsaWwK9coPUHGZbQ2uPtIu1jzuAh8o7u638/WCaZUO
RJWD9HwAXta3c3MN/0xGM10cxPehtVfCBMNjtUz4VrJE9NnXH5+2Wqk68KInIZXQ
28FtzU/t/sariTqA9LWbBQj2g8p9rf12JnR2wDWlkmaPVuS4d6lsa4HOLnWN905n
xQDStkDhgLODRbAWRT0czExg71YWQBpQFxiweP9JnB0yaLKMlGIL+hIkkbEmCq+M
9YGbd48ydlZI/Nf7pf8SRpsqW+vTBOrURbJIaEZhv7OLXsKXWsvIC+91r/c0vCfJ
FSTS7ZJrOs38NkKmeYUREyv5nBo3MLnu7hDXvWasHjx3+GUjScR8N940hTGvuwkd
rC0CGFA35oo7zNu3mhpPmoUTSU0vJguc7JT2I5MUFocCgxQZrXq57Q1vRjqBZZOd
LL6OWsegApGOifJ8/USXLwybiJsiQr9kYs7v6lifNOiElN8L21zw2cg9UoeuDaqW
XoicPsEk2eCYRVtdBLtVUXHZ2Fl5W4vlez5P3VyXSpY2L6f2QRpJbSrYn5SfHz4c
8CZOYk94chjuwh+vYnhvn2f6MaAUoVu4jaDbRptH29AznOEQNpPEljxhpeG9FfY1
4xurcBXhdkAgqw6RohKWpFIwWWnMyDWm6QzWwYvijAIS/wu9kk/fxAV8GM59zbGQ
MNIxT3jNBAeVB282a3+gsAsm3j5r5FBp2HFS7uMoRlUqsnEikzRTcPr+ulX8K3gr
SAbxocUSZgvue7URaYNW7vIlOn3T+weYr3n4uwGMr8d8TMsdeMAn1v74Zq5gtPJ2
QRrPLVzOWjJm3yqlF5PKNf73xYFqqd7jUWJaKDPzlz+66U9FcvdkwGlBF8+/MSjF
bmkKFHqHJx5t2Qf40dQzy7qg2kcyiKS4yJ2gnipnHBaJeXijqC0/LUvhxurrEEyG
8R/4Lz9o9jqTY9k2aVe1Iy8M+8EEUqmotQkhS1MoYQOg9cXEBxeMIVb25K0zibDn
PrSK+j/SyedxxDGQskdTRd7aMf6SsK46/547qz2Ex4+WR77Xp9W55LFnHi8Nk3Zr
G4qfN4iPm0BWkdSaMRrujXY0DiLJD7L20In1Kb64k3iyAdDaDPACpVXguj7zUtec
z6ZCwtl/gQOTLe4wNpjqF2liJkiMg91X3GkYqcWHKuwTSiiuWiJ3lTsaNn9rRi39
3Pw6tNYmW2S+sGOThwtbMgbLqOeLDHR8evfkZflOh426NmcyvOqzBHq8CthhI5M4
jsRzPCpEMkd87l8GpiDs+w/4pUZ7ToEEcK5o9dEY4ek/xU8TKB00TvexlAtow84e
4KrP1MHd6VriERi4OUmT1h92Wolu5tkozFEDsPxPsLRDrNgYtehMnv+A5qcSjEFp
LCpJsI6JS96l9IgT358PUBl3u5MgtsXeVWSWWr9p0tpcQ5GiYWCzwX8wRaaX+qU6
Jc7JeTauRpbCvhOz6+5buggehOERpLcQ5mNimnlQ3GDBaGeRqlWeCrtD6xYnVgdQ
N1JugxpUWfiAJil/iZwIBOG3prg3W6v5rQC5NSvIEQapdz09OiFsPnWE5sfy0vxJ
jBlTCVO0riJ/QYql63lz1uBZPmrDd446zWvJkKGRztkJAnOS65vlfsNrccLhQE/9
u7IcTDktU7BwskfYDEzT/J090stXFsk6pfyYglugwMwnc56O9lLNArPO417HNaSy
AExsSJiL4uVUl5Yfa3wk6y+jeM0EO+O/9dEvWFH+wyD8rOIfKkp0V9SFP6/gDNK5
eTwu0WkPc9BxW+AFxMZdvnSOLhOzc13EjWGDfsbE9APfxdoUqz45NiooJJlUw+rF
g/AJ3fQvmvELxVHn6X/AxhiDzKsTOcuq3Ywf+mMJsc5G/2RFJrTmkJvHr0HGvGcO
AkQET3GCW/xL+VUWS65jmARYzZI2OrX+vGix/B6UwgWlBqwNox7ARnIhREen7NSF
kBPQTDSPvABaAhIzx93K1z1iAOAeLTWlKNP/xmWezcxFLL6xfhvLKD0XuyUdhRKo
32EqH8fI8LTrv0vZ2gH+S9EjzAyWdND835+FdBwezCiGiI4Lh/5eikFEKbHi8xOK
A//vJ7cRwduu+WJZFJHeqiGw65M+u2vz7bqvXzc5KM6TNzy994aLsfC9ZBUL7uhC
tBmyhrVXT8JX9W2rrTXbFipE0nP/rpZWMLUHynDuL4VH07npv53uG1WnBtaUzySN
UL/F42nkv/+ARnMegG1CUIm7JRCPOy0+WRwX5ysmWZm55RkReozsTKhjNAW3q4cF
2A409j+fzjdq2WyBgejf1LRHOMcf9OdXx/xW6FCLfvgLckcGnR8WxmbF7n6sJ3HM
cW3Sy/L06SNYaHCyphOSqVAOELE65wXuDiTrFwcWSrK8eZ25KCmNKmkvJFus++IA
wzPeEksBsTKBzF4Ljt/8ZjQZPLBiHmR3SBfDwoyLtsdsFa5CPnrOQj3w5pkSq2rj
O3wOCnk/DRnfQRRKF7u5NoIkomCcma+DjS27Wgr6CcJB4somoGQ6xkwYGxMwVRhC
kvWMWECgHOQnej/oXUK3pDx7NG+ysqUFzYk9a0yp4tqCamP5plj5T3FIuPpIg4Mi
1/QGEcvSJZ9CO24EL4Sl+4a7FJU+0q9bOoahhwGa4EcK3oeLCNfx2A0QaWyRd0Wz
Y5v1+nqkCuudnZGmJz8XJTzNFBcbJH10n/uwNRT4y68JxbD7yJ5E+BWhLyYJK5Kf
Kfpt1ZGr+TwiDocoN58wJgiU7281uUgf87gKshO881ioDoB8VAdvxDltF21N2cRm
VjtGuqPC3Zo9yG1pUvRmS8u/yCdcrFx6o6tnH5fGNZtokSsVmFwX7KoyvrTDDLDg
xaSwerPViNNGTUUSelUAvlhyTRpJNfc380bU8m7xLxasTQX5wyLdzjuQt4pdI85/
AOW2KzPIiuZDfhmpCqLAADZ+cpeIXEd7lkHiOTxDVBzF0o04VOcjjkogQ8JaOTiX
DfUSfpj+9YA7S7GCuXvUJ3bKVPAv9KEYRsuWUrKvCO5dkg8y3SE4hYWAySGOecMx
M0N9gw/jIqf9lKNWGTnuPRdE7VJfb6vB2ajofS01ZjPvyA3li49mW//4O5oTKbKh
wsJd3+/v2Us1+fI4ryYHxZ3XVCmTmyUc/fnQ7TknGKv7NqUeZdRtBkRtog311ymw
UzQd+POouoICM2lwns16fjb6jWnffCXsl0kzl+SHRWrRmEsQTaU0VeXDZgEOlrny
6IlhaooBjsWpVeqXZ8cNTnNpeqnVsqhRht9kaBGfNzkjENhEZPCSal4WtviEbMGN
7cwTkKy06PO1BQoql3B2jm7mrSuF1je8k4MI/OPZhI0Li1DE5J2WfScujocPUY1Z
RbHuXSZC/XAmVKP4rzsht4ZGp/NJxrfG8IxHA8moOF6PcgxMjA7dAMtKiayZUaGB
Mmg1C5mgtTxIbm/SzXFjgw68ypGHfkIC1vHmv+ZwElEHLTNmuEHAUS5nciHoHIkD
yafeEfMHclWUQxd2jaB1XzLTrw0rjSMRnCc0ddLNEOenNwTGSNQmcPl2hSC8em85
kqWwCAGTWORSu3eqaSs+apD7snAmUj5UEj1e6eQsvfxecHIgwEmG/57eZvbxBHZv
6+LecdUYbL0GHIrzlPFO3kOEfBXo3opCR6HdmolnWhqkZiK2uJfXJCtEr740A2nm
d2WdQQVYwXg7nsHMCfUAgfrsaTnXnW4t+yFRBVhyNBpdzL38OdI66iN2FTPOpz5h
5KHjNVFMdBtl6H3oALvCuaT8Fov2i7Y4tC1Hj5kyFIu3Y79Gs2zNHMPdTaMJutX9
TyX08VWWMh3yCduM5BZTL1si975xT9K4cxVxTOPjydE0UrMS9YyyDSK8aMNKLATF
i+HP9HmMJtcrPTwIL6Sv0B6uyVpYiyAgChhgMUoUf8/AOcMfw1qxTlV1WzP4uzJn
AT/gEI4Yoj1WFFAi6DFTuQz6KGx/bfv6ekfR5x9D9Z24JhpLuQSeuHQnGyIG49Q2
SGm+489UB9Wg65sbUMjm0yH4ty5a086cvjhcqjTHVZeTE7OyE+n1l9Yno1JBNbtJ
+OhkmTjuBlJOJb6FLzi4SGcg1WF/Qhz6I/qFpESgDKqkBVsDEIpgY5zMo2463BY/
DYe2Se2bxWC8Iz0jV7KiM8vkQPL2MCOoEDYoKL9x6wy22QiQCqa0GgdzUlbjjImz
QDzJwORSgsZ6EmFKidYZ0b0aBCPGVQp6yoDO4E4cb6BqeAXyPVNY2tf/2DWLCbC8
EWNPZ7X6GWUAxAmTV6IXzjpJbDcjA3LQ4ln4Q2nEwN75xYWR5xn/LV2+Jg4stCcM
i8AA7UzRbd+veOXZ4iiNtR0M4AUOCgd+WtUfHQc4CipwV031BB6JHeROImTwQyI3
IkPtRJI4Q+6jtXKfTG6c0ToMkmFo4sFCQP0gZ+6/Ptb/O6clzKVDsBzr8O9Cu8HZ
2ziLn7t4mXg5DH43vIy9KHOo7LDQNFn9s8v1vip9/5bEeIEAgOc0wEwNpOs6vSvE
ajTrn93fqbUVANRAhRdcI/Rxs7p0EN9zblhqwv9et4SYfieuIYWDIm5rH+np5HRT
vLT9PODKudDfgun/xEmoavbSVsKmnM29pTSMh8b6Y/9TjomsVG7RZSxyETvt3FXk
gg8y9lmykfBqr3O3NMqzDJH29yXGruloomIAaJD1UCwWpbkNxNIjcz7n5otx9Fgs
dRFdUbqk69C53KfbmUP0HTWLUYHbf6yGoVYfKItwL3dfGY6eiQnYqrqv/i3UYyCl
ennoz+r4G33T7PIgMKgwwomIm/VvEykGoeerRrh7KT/rqX9p9wBv6r6eKIPzh+gL
9ASeGjQdmFG9JtPpYMXYgWqHBh3riK0v97dMvxEK4wh5T6SFIj8KyGv9j5GYKB5h
fSNWoQjFCYRVTxgG0WOi+8jl0zKMV3ziGNuhSodhp4XR/4CZI2X6oMpIG3Z8H88X
9FvY5Oni4ljux7fySlqml7/eRbNnkK7mdD1V0dhZVSk8QeIkPdP88J61Vipu4+qu
ZXUKt1xDLlQmkt7mgmx08STochPhTufQ9LfXwvlr2rwDPYo90Gm5WrqnbctEbjfn
vmTtifMDMQn4wI8rOTUuN/iYfhiTyI5XdaM2yFH1XdSXACYnLiqf1xk5FmnRYc9b
sKgsfhHAG4Axgw6PRlv3qIlv2iKkpMc58jsb0xFh3PPM3UU5VTQXRMh+26AQKima
HxUzbsVbE46/gjDoOj3P5R+O0erbMEGF18b+RM9Lem9YBdKlYAKVElWkTwo+N//m
T1HfE7HtjN21RI40aTYtue+2cN5rxmA/62HMfsn1eHcfae+12Dpck8krSL46hKGn
yqLtMKA+GcSgH5BbJgqfrmzh33x+utcGy0UXI8oAMNAlKQTf2IoAg6oDJUEsLQj/
axQmi1hco0IPI9URw1uRYEf2BaJMSGD2t/eQwB4rwZp3OOSEMBuquTQLA6DgHvVV
5UC1z2njOIjHUG9uarMbDuD0O76/uAJVgX9lli8C2EYbO1xQsImigSormJ1DPkA/
AbyKLaEBCcgOzyg2rpy6+XLb+S1jtIuYUQOEdteDVIl1LgDvwvrpQghVv4411l2/
mQhVpw2Hg6gCLJBqF0lmm58ydNMq5JwjLwGM2Ewja//vPX2Rp/1Vv5drrNwKSEoA
oeG8LI9TZWNvimDAbATiZO5S4p7AxbTpC1awJehpu1AhNGFdibpXNxNRZOEJv8hi
+1sVnVJB4qevbeOFk0gSsXT2rDEyRjefgET7kiMTfPSfddFL354x/TDI1QSIh39q
e7JNZKly+NIUcD0jo1Hju91viOVP2Nv+skNSgCgmvb19+FWHcX4bLdZxXhm7Xs0a
JtfANY1oZ9OkxX5clsUwhtR/PB3SDBVzLpwQ3tFuuPH/WgZNO7QHwzdlZGUqLmFr
CPHQ6Ptex1Di1w1o79Fft5juWLuHGSWpoBMXPnZOVC85240JnpvqfAWqm+dJedo7
HMkKlV2FOxT6TA/+H6WMY+cA5HkQcBBLeH3OID4AxcV1DGMMjAAc75CkUdkw0FKu
R3T9bCz6CEZjtokBpU/3NXOxQd3re8PmKv7RuUt0JJa8At4sxd6dgQGmqAgItr8l
6RClLrK2s9UDcjolwSo2IXp6aCT0pk/7+sZr340flBSF0MtzY91nKf0jSj6ZggIl
6Q8CuXeb8TRNhz2hU8M1uRw3eQXj6VZiGFWUkL59MBjKV62K8x9J5BN1qlfqx6XK
kvmVW2vNRKC0VOXyg/VXr9ATruf3uitjRJrJjPVQ0kRxlrfuGkzSdkgUwTXqzhD5
D7Y8eZNpK6tM7rXZeRs0jKEJzuRDO6lVsFYpEpT+OwCyjFIiJM+35J7Iz3ZTiPkt
W2XerQGpb4xF4FDtRG/9FuNmZujwCkZH4TRG2dEKvzJHQ+0IzVyxvgJvB58+zXdx
6cBQEj//sZ8ryXABz8i1afX4YfMF+9n0QLdykrPwhbN1vU+29rOBNiYVmnTEsbq/
EXeSRy59Jkw8W9sMlrbfYLIhM142rB9Qa7m2NS0pdLpYDu/SwfMPjVoZO+CZw0En
X3R/fPFSmSJOUhF/rJMxNmjchkXW8JtE5Wg5bLMaewJ2Sb2aKUjGQktdrMbKtc2s
1daQbYW1Ar/3vcHzRX+9DrQSGIhyNyz5B8/7lkyqpHFwgWl7hglEmtdIYOiWBmx6
Er0ME94/xueSLm/uTuVQDN81EDQlkPD1A2lAWrJqUgnATQeWKlWsnbqBNTjDE7fp
fbmGt7rf6yXAVbApcDFvPp3ppKyVegJVzWzVl2ya6tyLD6oIJqTX3ncZCMjWjH0f
9naCIc04TNfZzIbZgz4gnLVSBythxS5mWhJ/owMNzuctApnUpr2Ps9TxNBqKxtJZ
RPav4hjOc0UBSZ73hxaF1TOo64fJupLypDjahy0H5TfYOuk8K0K3F5x6JB1vF3Wo
Cj4id4+Vke1w4cdrTdKIBYTEaSLHUkv7q36EjYXInBPQWVXC1ti7e2sqfhPxsIsZ
OpT9TjZmjh/W4u4bTB7p+TC5fYiQEt0R94UozYl5iLo7eE5kJmb7KPMTG9efIB0F
zNN9zrXo4l0UNpqDxO49GWttZNXYbqjzDF1NuiFovQZqBG7pJP3tLUm/OjXgQoq5
bJVrxbGX8x2mobIbOhn1hPrU2lF1uYK0lNugIHONkHSPgzquqi0OelLMUtti4g6y
NV769lN+jg5EPoZyhSNAFVMo194Gt5VJULxTU3c30Wh/TDaJLCcTL5Ilh5aVwtwo
Z958pr6gA/aMqrXD46BE7u/fzxWyU5BRv39rvenJunPxrjKQLJiJLZr1BjB+vBq/
NLiO2p0xdSRo+6KhmyV64f/vu4AIIoGBTqtEOWjF0lcjB++VFB/P0320akiNorCK
oF1KuEpzq4hQSHujfm7uZ3a+sOJy5xR+L4QDH+4vdtk4skUp/DOOlFEHHg22trcw
UW201oSIi7xLKh8cqA0MOjXxd7B9w060XrAGGf6sxEKoEn9tr8pB7Iiz36aMtlk7
wO/q9vg0AQGYMoZp4w/mSqF2LZcMvSeYFNath5GgcsBu27/zvPZnBo+lrqlSYcrD
W1On82e9WIrJzMO1IatQkvzv+hZjl4wt5LjTAyZqptT7rvUF5sG9qU8zdTNlolba
okR7Cps9O1pBulZmwf1sBc/m3YiUsSQKuFi9WcQC78uuwb5g6JA0xvfq0jNb20x+
rzRTSupiPbrqZbmw2Qu9fqOOLDJ56TnRWEpBGIHe2fFUY/ufVFdNpbFQAeMZroU1
MKgmpX5QT9gPcac5lFAnM41rl51suhOjOp3OBNrrdRRtBfe2MQmXdIdfA9JRLZnu
kCb0h+5mSDnYwR/IadQe58Yi7laWEBwlfWphT1fE6RatdfOYzNQiObvMoe+1jRxS
Z5hB91BsYiWkDJ+3fIzfzpGcdlfnnNEth1W1lmxWK4kLDRRSCbOLpREgyahJfonr
xP69QFM60bcmA6CDJ0dhg/QGd3+mEBFExw1OfxlcrtQGdT89Wdn+fnluBEUGnFwt
+CTQ2uLydTvMOdbC3aI4jRjN2DED6LGDjeCq7Vdkizz7jJnLjtCVLotBtJLCVCM2
gRdVz+rZhxdVOs8mqGuVzBf5cObX6Nxrs07K66UG/AQGrX27YNAWsJzhwL7UHqjX
32QSdYiG6+t6kO2fO5PyVMpSqohcah90SABMFgeDkJ1/+62ToV90ZKfbjFshGPap
bA/C8QDTB8S/066yPgCD4hyor09xZtjEjtcU3ic1kZTiwhVGqTAt/zaHgfAwcuD2
nksPR0v9i1ZBXqmNr7tNdLLhjDnZOFo8oEUPc65r5sWanXfUwTWTI7kk58ZIr25r
bC0bBcUwOicgkpCHyOMUQkYVvRXCZsiqHyJjv5VW6iPM30NercKgLVV00WiB/ckx
3uTc5hOUPZdZqrU4P4SpFrY5DuS1yqaq3CPxN+mOBzdxO0JwRT1Mgm4OmOgk668H
EbDIHnP+NtE2bntsZ22V/MHQC/hFMEf7mNQX+rfu9kwW78JN4vQwCIHVEqUja9Zx
RfiHWZx8vmR4+H9QltLkbB1I3Omau8iSa8XHG7YPFVxHMM4FVwo7TC2QxoAOoZ/b
9k8IZkVaHjcOK4biMEyfrkYvNwp7gklwkSPyAMCMM4lXtgyDxt/jUt9RhvBZpeSX
XrqQP8FSTUFju2mVwWo/R5NSTv7FZY7ZsRVe2URQHwZH91H5hjCK7gzlJiZincBZ
Oec3Z2I9Rm4/+B/V9k9xPvuId5FVJwulVNdToiVgPrIWKjJHftFWQUQzx/HQVswS
7B5kjU/u42ZcSUM7vznIfy4nKrzou4fUbRzQgEjQoHjim36D6BghBSWeqJTjP4FZ
GaTjepzhj1jBMzmbahFU6WG/uHeOiuiZHkOU9ZelCg1B5OrESJuW/Bia0Jj00Xe5
8JbSTGSnkXDTh5eze4KwMbjKLPPnF6REtp5ZQvTVBewrBYgYlvPNIMCiaGWveYKI
8Twxb9fgGnMIRO2hHitojf+roK91BLiW6+vGzi8iAoj1XiMnjQasGfTTIEHP5yFE
NxRVgRiaeEAkMqaKUy2nPH8e4piHKDxDwIbSUs0fiClqlitd+1EOTEPhU0x/yxTa
BQrMzd2U6phz0NWKxHVPT+8xWuk/HK+qGJn28arwbbmf7ttNExcku/oMVskPLEv6
s3Xk/wL0XIHsXI1HcKrC2z13SjqfwZQdKYY5SwbfqMgyMMCdLrJdQtOHoG8m0l9I
5jaacAZerUtsz1nLFXr/tn3DCg+9SFovzmm1i5ZH2vMKrmMFQz0m/ppp55zBKwgz
OUTQGrV3JYNlLOS7jvvr4wTuyl/lxJ3pG0NMlJrFdpq0LbR8ZWOf1cdacKeK2XQ/
r5VOSI6L5XUzYGEHWvn0qedGs1NyQPuplQLu9uuDlAw3NAIGohhCBG/x86nPTPHf
gftYCRVep7O2LLjcFeG7mz5Qq1Y53L8dcKMWSsPdJuF+524E67hOGRuUClJJpQcD
X/NIIEowiamLMD3zA+L1LBbowfMd89oYPyLZadrIRDYKN/Ph0i93z7C3kKjnp8p7
wGhSk5eraOWZNsm7ahlB/7fUMwp0q25iLEeHXnsT4WeCw5I7I9QS5yBOixOFRJYx
lvjAS0v0tLwYXUdxdnpbvY+q3h+ZuMEHJKUdV1YJxkTAo5SFxOfXoEf2XIDbtccH
5R4Jr+souoeRhc4PkB/eEBsZCW4lUS4lOejCYAr3ztUo0mHm86t7P87YgKN837Ox
80b/Wz6iei2mXvFGvcsBZwM99tofQ8dayLph5KaRin/nE+VmH/vfv/BNKkzN4NoF
1yC4hhf0UxKLLxDLvNaE1lknwpP04cjW2X05cCsRdzRi1AkUwomnE2EY4k6bexnk
Zu1AmNSzvmCyDMGwyrMc5FsOSlSrJhX6HWQonaQp/GN3Z/48sASpM5Cp+9Ejt2Ar
9tyv2Q2zC/xiI2wPg71EDSm3uANm9H+rC2teYpC4DHwTnHeX8jx4Hkmj78gfgGb4
R+SSrhJzmI53/D620VHzJ69mJitcPrJa2wx7pp48/sMf5S0DakqvTxZsUscZmt0Z
GrUPwDOTpByb1oBLDeo7WAdpc7tKjpZtZxKLADj33sn7c3b0IO1UN+R/Kf1a58Ii
1qOV4cn8RI+/rFsyqRf0PpmPwRQt7R8IYwq7j27FO2kQjqcg6qCKXH7xL+62WJ9G
X4IDxDZsCi56NtuNIAFjp5CvVUTP6z/Wc/pyE7wEovIaTl0YwT4luDnFmnrMSxxh
Mk522EYSOJUYKLJPTkIdnOuXwHosGddrqDNT+ZV1X2fHyxq8Vi9AuSU7T6WEfQLq
ORrapG8NtwVAkPcmZyMbob+VBZ7wKGCnv0Gi+5ayFyeg3NhuEs6mBWUWEFqG5W/b
YdC0CaV2Md0bGRhZd3NxAkv+nWBP+58GsEnKiAHUwwXWGo0gJyV6m6MWEWsq/sGm
74cQ/WsJCqp/EgdDrEsp3FFgsMrKFbXgTfNtHNO0HNpdM7nUWrcY2AbTUq623uBO
yQbPSuCBdmhhCw1UTetUPhg5EaNNpbPWl8cZugaj9EIFwvJTGXQ5NgOt+1n33SSb
/g5P4dG4LCgXP6nHT2E67vD05ADKugD8vdRz610pRT2VGXvq6ULyplygojgipghU
dVX1MeoiTTcF9TeNsH1ZwvE6VQixUHpVPWFc9u4f8yDZPW4sBqd7RiEOuaZU1YXU
6aoX8c6AVpwF2MnCYBfqty4pWb2ZgiYpPjm+LH9C0MJVU5gwX3G6srMerMxWA0wW
O87bbDgij3pugoW9Y/F3N1gHI6TrkvBmxKZssfMj/DH8Nw7ugsrhn/Czy3Rtivsy
QASMorToRBUfSdwPwu6rK6EziRAlRuTJTupm7WoquQJis4CnRO917Rc7x0DJeiPe
tlJsZFgPGqKxFraAWv+L1LXgjCs9Hw2bi2hqa/Zbf7KnwbyE9MKgJuKkuQhNFneU
XaXQnAz038cuWApyU+r+A+vXnrSl4hN/HIjzdwokXYNm7RonCq2cVN5AYQCtW2Ut
sCMXBoClmf1ifdbJ8wIWlobfj0Lr/Q5RqTTPYhuTCZmBGE1LmUTfbyADxD4ZrhpD
LoBBZrRDaOdcZkxHQJEQnHhtrnVFdbmJ1an/0JHQOgTKrjBdVOn/C4EeC+bMyy4q
7yLc5X255FDe0oyFsWEYMAQRUOdggKX+eHisXzKxM+pKJU8SO795aNQOuMtcYnG9
m/jGjga6+C/Cy1Aw9J1G5UNtjYpf+ZvY4p/8xvh65mz1QZyU0ESkGQm2DN+JbrhB
8VUntOuzW0erriq4y9i2Tvoz+AgiIagKLbjKHorUFWNAIQ780UwVZB7kpEEjXSt1
9wFFB45CzJWAeEgD6pPIpE4XwocXuvYINU/1P1BUVRYO4nQXLXYU1aeQ+24UiSSx
BJaDepuNvUR8Osa1FrJqVaXRx4zBMHnc+4G1yeCz0NV4mSVDBgbIWIlB8iy4geTy
sfhIAGHp2UbhWqqkWBOnF5TOTjnVxrdHPaZaGsM83Xqg66llJ37egAwuO2YDHpnv
MvqxuyOmZNJO5o+0fG4QRAv49keKxe7caEfnPuJqA/Nv4xycrnRKDe8lzG6V581k
iRJ4BCRihwSccrGv6aw1O6KFfett4G+qRahy4vqq8Qz8xjKfwpcMzgdnFkj5Qe3+
WscntiLOQJSj/jPRI/hLrxeB2AAUo/5VuDgKsHBKVlmgxgjS6dG++CuO6IxRI6Pg
F13bOBdxfKKXkR+9sLr7b4ON0KfRv2cQcyc0Rt1l0GiElocz7/y+uxI5jOalFMIU
eU72F9lsCr72bKjrFCH2oDlVvVBOaSUh7/likxfVFZn6y+bbWqVMIgf6gIsuDxJj
LtfcCpPLe68EtBrI6g8XgEmlVVrUkN0S8qbS9FVkO4jxI6MZR5sP/ph4BDLnArg1
4Xf/m+oXl4BkZBZzuIjLDOJI8LmqOplrXGcI1Zixv0vPsdGtIRg0g48DdhxPBzKe
1dNT9bxCnvx61YUt5A79g2RcAJhsuTmFklzh2wJy1SDVHhuOEtUdeYhGW3lYXpWL
V+PQGvbRQDYKRS7O7IVE8PkNdtC5Y/isM3K1vqjH06cBSGL0Km53ApkMKIJBZ65n
H08xX5AeuJW3TUMJDSySm1lGdpIwf4wZln4hCHLw7elLE3yAEW8/7eszAEZpcV3m
kwCl9d61UGGm9OFAyj8JZ4w6xNxeThzgo8NdL1CgDNPH8kjBwQh6NJlWGLBkE05b
5YauFbp7vu6Z620GGRHtb8hkF/4yI4sohxUAVfV3f0djTSQ/JJzrm0PuaOBeOErC
NrsQyKGH/Ke0rCv4eduYiaeMat7lqsiBxMYK9T0MSanb4pimdHVdYQNsAomf8+7J
Z2hwkr/QfYDvWzaBlusDKP6nza8TRRZbBtsJe5QoipGx4Fn4XRLs3aG7ZA4iqs06
6/RCB1oDi1SvRUD9pXlb2EWhg/3sHzIKbPNx0ES3EXulQh6U61ZLGEB3KN8rDw43
ivy1rpt0x6dp3MauuOhiMNASwa66ZQV3/cMT/UuWmftwgA2UGmSQrBTVXJJQj3g2
GvtT7gSaG+7+hOOoEsqPyg643EfP5+fJzFoPr2EynyK8hVZvC80lWeOJR9VbbedN
DF5fAwlK8J+GBwc0oMSFnRBu6JHj74tOO3iSt+f5hDcY+izjRDcn7EKqGMbKNUne
S/OzpA0zqHC+tPtM9vg0pHkLS0IlU7XJKxoctg4Cm1Or2lAI41cP+3v6O5UP+Uuj
NuQC7CG6ZILiVrPDJlvVy+kf7k0+rII/9UIKh+HZRt4DI5ITBMEj1anz8WjJ5eSk
lfWz3aSKAYj//+PJaEK6rPBM5EVc1fcbFcy6X0nFPvmRKS5TMlDGTXyTV6kOhwjb
tsA26XJMaJe5fLlXQRnq1q8Th8rWqA9Z3JJT6CIAngCP0+7JyG0pTEQ6svbfNwfx
lQmXcMuIUerJzMRm2OxTrHfHm8qPMGLvkUHrbXefa86mPO8Whh2tBWbnnhjm27Zj
CcYFs11TcIDkwET7/4X5pQcbxKCY90o90D/ZZ04MlPx33BGJPJNU4dExiGAUmwB7
IfAl0yvyuuIi66BP6/WIuvHncrjv+YnNE4atl5SfoLwFQi/IqMfrbZGHIyxpAO69
7yLaC6heZi7i474DfDz64cxWyx1yV/O1JnnXZ0DDkRtwSoI862Gihn+DDRkBQbFY
SHM9gj+/PNMNo6bSdvWdhSyxLYt3lgp97Q6aTUQ/A0ijaOaFu8ChORZZe/K51qMX
4biM3B0dHI9wKZKSbjve64hshfYccgRq56t6N4foNWyyAy1VdGgJxDZX9pcfHXyh
Ehh3ISYayq8UafjWv9bPc3QOJnBtKa+7CzuC8wGnlOLzqRxl4rxsW8F7S3X6YO8l
WTN/0y9xDTF+tBDVy04NrGO0gOFYrjdUzx7CoGvJRtgOfyZvY57kDOc7vx1rIfDM
2cUF5CmLTYXvfGavYK/Qd7oK8f9D+9FDeYMcveaZboYOz7W9vQQMlEnroAyxRyEj
0YiGKPJ53/xH/DXyi5RHHmKkSp1pHonmGMsk1SMaI51Y40hUrIY+86Hz62uCcjvA
yLcIHnfQ8WEJ2n2KkwlOmdzqw4fopeS0kXlc4cXU27bU0OXxGwG7WnJP4ucMJoT7
BIJNEHc8cBYkFBuC1MI751vTIsjR1Vv+eiA9bGTxCDw2MQ78FlWh6nu61SaNVutX
Gm07sHoCUfYlRK6Qc3aJeJJSnVz8pTrCU3UraD+wQb7S2VokUx48nV70of6Ui21k
3jcMdzPxBzmY1pHDh9rP9AK7E75smBHZOl72ixNYfF2CEwxipKxOtXkqQAw/vSLz
0xUvjOP+bGwILPM8SRp1lof8W7CFGg0BfoAhCPCnlLiveiJ1UT2byz6S1Cpo9JJp
4AOIwiuVuiAFOd0xuCMxA5rOq+GZnbO7SWnjr9P8KqE2PtpMwy4PhnqWXc2AUYY3
TV8NJMaPSCgsVo8BkHxdhANLBct46Qloo7DT3lmrEfYIliNRVCVL4wLNga1Udkj2
oTnplCQIesbEcYCudNyZeBsWJsoBiORWxUVR2EBEePutlk32609GEZrLy5SjPyKb
mkSiv+G20jGrw2tA3vRmcOX0OAZRZhJ0vG99iMa+c7sk4VSpssWf3gZDdp8CccvO
+QJKERHJJ3JJQQ9pGmowWeH6GYA4AkpGkW0kATG/kYr1UzxZpq29FMb8NkDCp4no
TVSE/voMbtLhgd6Yyro2Xio79HgrrB8ugSwtgR8jFhf3zA/KduBKqkPK/Rf7OA5y
RdWhX1Efv5TV2pJS1kzs4omxFK6JKr9XlRBmhBFnDAFIs5Pg0A8GDYwLyE4cj9hG
CRewJ5B4yZ3YCwDR305UKZN9rEMHH5uCqZ8YeUHYyEzQRrQoEfKZm2DnLrxg2Z+x
SrKQzLGRmkyKFJois2MeYW7R4M9H7w/naBh6Mc6CYSlikyyeNm8CudoR3jUkontk
B8DUrnsTvLX/tvsL6nH7lGZIAQOn6J7YH5My0UHMm6pQwXmXGOZtnDMoUiNHI8Z9
vIumwC56bgo4eW9IjHZcUJfMwzNXw3rkrXu6Ucc8qw9+MXGk0ab6vCWvRdBteXWV
Yb3xTT9g4By92wvrVpf+w5X5jR9ty7exa7/h5VJSWw/qpY3JB7yQBCegA5FKVag0
WgZFHGHiLOHgyQHQKY5SiMyfPDxAGrielD836jTlJgBSYQ/xKxzbiHBatELr5HyP
OJLS8EDIMdmSf3xZlQSV/uzshJW+sjM41iBt5eRw6nysABw4FwYQyVM8tfxsA8J+
dnJcN2ElT5U+B+JYCGlsQqVxwfPsDZWXgecNVKrmxWudubYLJJBuMChTjfpmKADg
LuJUYEkPc85P1ZT5RruaohlSmDEFh9/f3PcrIHSib0GLtpQim0IMkO4A9y/lnz9F
GU/tXxU0dv45N3XciQ/sqh5BzKw1KdvQQzdLGXh5q4kyY6/vMmT8FtGSEThvEpAy
ZrzSj3+uOoviSphdKTrlgT9Y29wRYotccsO41WgKjeHsKhXogDhStpTwrJqixMDi
lpA8RRfHo2voT25NFKkfRf7kQcbwdDUMK65pRdEFNO4Isua7Q2Gq8hjV315cOpMW
uoge51nJTPMQrSocP3wjcf2qc3YCF355IeHY62iildG7VRoSyadNVXbtgOqXR76T
kkxodWiv+lqqLtHH8veuuEtukI+MTF5JEj0aFE9V1loU2T46y9BU7BiAp1DLcFHb
+mn+djwKPROjYAxg3Ph+CpU1blNJkEQttapzq68W+NHY/WBsPTer6LMP2vcyUFDa
X9XQc8WisEkdmaKYLq4cvX1KlKrcylkMXv9gljUqzZ2/oNnoKgmRn+FTL+myAtcQ
/YSUfpECjykk2sruvSoTYdx75Rhs1iugDVws1wqRI9sir1+RKjXvu+eSvVnn8p6Z
cX96E8NxlDIjnH6ZosaKmmVED4sxu3z23YUU7E7tRnZBj9UQaZLb/+f6Vyv0YB8W
zWP6N2XJMMfIGUA3unQsrahaCIXjcq7zc4eu2/XI6UK+3ofElEV6MDW48yvlyPGx
wity2e0Viyh+C4YSJx148b352MObwU+zf7RHy9qFqtQDCX4pZIJuX1cO8UQYvjQN
L/oB7KrduxsXNO9GYDkiHeX5V+Cx8TwwnDG97o6CI+HYOCYn9A0A3ZvU3wBnQvey
Zw+gkZLA4Olr10UzGzBibwPoIsA/5pWf51gfDEfugBkGX5wbz4gdjPe6hv7O70jf
8stqqurKZ+E9BqfWwwFtgZjggghr4aH+YpJKBW75jl3crP7i+btBL8CjrJUhNyTP
LK70E8VcPm/LO+WcKklXlpSNYjZK/lyyocdI1kuJT7c8RYjQrgf5XBRJVly5Q7P7
GhQ7t+TWkmw01g4nMlBcNbzPkErG+IzwEFXoRcslkISP0C4caUyvddZHHTjzfMG+
Sc2e+tVICTfdOHW2u5hzD2kCCsRJ29sC+gDi7C+Fq53wG2lc86+4y6QbbCwJycpH
UN8JxBi1zh/ZvpCDIcCGuEezarDLxYy3zMBhZOPQV3a1OQmYdiO2Zj0W22nG1XK8
t87mdYkLL/EyJ8efq1jd04LguElOXxC7SEYRYHvjlyaMiLDek7gBTcNIHxmFNGTo
atyhtdMq5S6UZLeJRPD72nL+/ELAZzl1PuQ7HaiRkYqqJsETz4po3qLyb8VFhUYc
sZxRu6GzwlM7IIrz1izsKF2neP7ddI4TcC0pkUsJJzU=
`protect end_protected