`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzbxWtePNA4xLKWL+TYXD9ygPEOOZ+QBcvHmkPVktGsmO
A5xYYUG0v99uaufGYHTowYmSOfVEoABY1HUbQWs3QWohanyz3IkIlu3ZPA/Bu4gR
JBkVJJoYXSWmIN2ouiriyJKMTpbwzIk4ZSOId43/BcGwXkvxLYRgO+/wIxHXURKr
fBI9gWwHWzta8sceneOOUHTD6ASfLlg3OgtkrXlhU+ZnHaDHRqK3qKJLua2DjmKJ
VOj6zB6xuAoO8WIKSV8G5B4GIVkWuUgPfMbmkyyFZxZgF4o9Vgtwu7/Ln8JFmiex
K45s7a4k6JKqBqsl1zXdfwevP5BXPdXeH8EQUxkhMMwvrIsn/WxOyQg9bmxKzpaW
u4urrCrLaEc3c1KZlLiHRFExmA7tOwXOExy0cKErWuDqMYwGLGWFX+ps4L0C43TH
aRhieewra3KGHnjQYTNDlOLTtFJWPHTzTMGYwtT13y3Yi9bKHWqqf2rwpV4yJo61
rFkgwmV+0mMIYnaFREzQ1zYwbFV0LasSeysDZeD11cLfPCj7vtYiBFl0bLNVvuNE
MJ8jIudfA3e8BtgkT+aQAMmEVpTlixNdpuDVDXBg2Rb7kLBOSLyaDtjoh/J+AFlG
zyeACrnKiJz+60d3FGMdYMgO/FP71nieM1KXqSHcYDOW3faYmvQsGcyX6kCkaQlN
Z6KeQLc8WPzRTcO2IaddWYxUwLEm+TmJcklkY9rRasUMXKIcegK4oHMr0S3f2kts
/QE8gB9M/C9fWYHfryO6m2u/vPf80h2sOKjpBRez0nqLRripHJb6ln+IK9KaUvhx
mzBDRfiJOOn3axKTiqWYCq96hQX5LkVf/OVXlUyM2DJtzmjD5uLUg7WI5zH6i082
L0kFWGA2LrOQy9Netw/o8mwSMkqjQPYfG0Wehyv5iZoMI/hrsIF/bLHQiZcjyNCA
a51RSW2kUMclxLbdT/Y1YNKSaUVLP3AF21RSrPlO/gkdfgD+qiNhPkIpE0fouRfc
e0mYOZCq4Ftfc7/X7K08Z9c1G4D/huVJTju4jIwWhg8pI6PC7Fks8KLWwti8vnvU
mAgkjSqY0vpPeKBPtryNVJz6s/DY1Htk3Ei0vXuC9bU2IJr/+Sq4GPckvi35epiv
cS7c+M4s3jI/d9HZDRcrO5k1qoQP9MIULlDzPDCQtQfhzEomkgD+Rcr3R/WfB123
DPD7k+6s0T5DHSoqjD1H5WRiH+C3Lj2VILUWTmj61B7PJT6m8X2fmmoL4AImF380
AqfYKjdfMSDbjwsEX1eL1ZREWpGfYQwgLPm9/l8Tz2cEPUOWje/yzYRNtUIucUpw
8fZBTSM0aZFgVyNdt1NZXWKuxMzCr3ORiMjFecncRZsjSBilMgBOVJBoLE7+1sE9
W27fY6HmA4bisH4ZqVxp5ww+uJG0Dm9RCY6sTh7exhURXi2BKGByTghSzpkMDvo4
4oLl392pJbn+37jG+CDdQFDYczCmOdnvF9JBiTOqBmsjEqweSxKFMNeiyTg1Os32
cmH4/F0fFOVlEjjNV+SdUHLUzw08XVlBor0ooMjpmr6fIurh/J4FfiTT6FbTTFyf
XsCyreMXAaawW2UdK86K4xGmE8JIZJWHjAJZEoBQWAwaa07qUITcoECcJp21vU7n
WFrbFHKKXhqp9ymnV009jG77iiasY1bLddHXd9G3tWKij1zh/fc/u5aNUZEK19oK
9H7OOHSz3M9vWR5bm+dqdS56atIiZ86Mg8AJlau7FGaHDVOK7JjpHcFs3fIm6ySr
s9QcJrEZ2fKTZDsIWwlAcdRr2snFcuw+c5anCK9DkKe29mu/9Wue9aSxrBcczIsp
7at4axfLXZHRyhVLR3e4WfiFAngk6HnirfXlKsE4j0I+G2XmaFaHGw4fYZXf9lw9
OniJ63GVL7MWQ3RrnxZamk3nGj8OjgrqzJQ59gFUZhmtvWyi/jECFyeg5JE2GotZ
OcxxRIxu6vyCzrt8Z4nAzHfJnFKRtoBd+kkngV7HboRKP1JN0+Jhd8hKZbKKuivZ
54bpkf7uWj6i5o+hty3e1niDNSyRc48E4rUA6ZswwVjxD+P6GYci5/A5uP8rnCqV
uAgY8Qz5BGLfBeZGS79UGl2clysPPPu372sLVitNcOir95PXzsN5MggKOYZhhjRV
+IFhUZSLu1SoO6hLJ33ZS2/fLIkA9xTMo0LnY51zmwDVr0X6sEFHXTCiiCDjUvCA
G/vLgOT7yPGPhn0dcviQfCRpYz12+03TlHUyVzr1MD7/R2O7upvz9EyKCUX3Y8kh
4IZ5cb1hQwPcOCADUNkJ5I7vmB6eINzDzW8iY7yq24Srb8oGxhO0BqA5Bmtxnruv
erl5ypN4eRQGEL8V3PL4MHvLaYl2EP0BkjF96lWPtHy+rXeUbdr2/Ol9y+KGbwAo
Vzs5T3+9e5nOa+7iVavHeKHX187Um4+vKNbGD/uxbPmV/sFLQBYKXPjCjexg2YSu
D2IMOlibuVTFGCF2+mdeg1JKIoqIw5G4GhtPyH1Ev1c4aC7Vp/dzBNpl8e1d7Wry
JRCbXFutpfatYevyEJ7Ru7v0RwmFW6oFDgmnKYj80VW2Uln0FwNh3oyT7mxlpXKW
36PY8gi2D9SCRrPanqdMUt9FiE6+2QLuu2VXAUE0KVuT4njMxUCUIzuwTlRR+k3c
kpZa14VdN07HzUBw3qk6KVs2XBjV1Eexb3+G1T2KadzQwQI6mHcoW3pg8GjJalit
8m1kHI/n2lC1k0RO0bQQqEmYxQ67SU8kVIjQQdleN6AyacBVRVxD+nZvhwX2TiF/
HU/kvvV6TSNsDl7eeaTOZhcJOpsUSH2Y5DSS1jXJHLXYlsowkuaRfY3K+udurEdG
VrrsnuVWy0eRPQXBgRWcyBrrQp6aZwwpH3XRhGexWuJNgeciaIYjLm8xi/u1Ia/f
v6vNBsTY1tDwdClJozhxq5YnfkzzA/WWCq/Xx/51/XBZmsP8N3q4pI3ThPtDSCDQ
MFE3JV6I2SMDsPajkI+WcYexz+oKHVUKvbA8AhTIlojNEfwq5O+av71fjveypWuz
yAO0+qsVSoOrsooVMhY+/npdVOcAEdgUrUuTpunQFQqSfEB7DxIuoEOqDqF21VMw
b/S9xVV5zXljIaxlzyzQSdzODe6WO8DZCCJN3hIgEQcxScBUVZpkjtLn9gsWiLtb
bxUP6MZzQGMV7UpLP1DMZyjLeM2OUMwl/jwtq3bymxpo480k7siciyAJoPfCursS
RkzVSFZJGWOts985PlDGiR0XVAWWRbshUCEEyP1EA2xRa1N1efvoHHDV0lzy4H1i
76yhp0ITIxhJ69YEaMGrIdMuXOwp4Eck42O4zIG6imfLq6nZuD7L5Hb9KRfQG8pM
QX8Ofug4+eHGYX68je9HyENaPSW+Klq0MXf70MQDkMYNsF9QY6u1uq9TNo3X3A1W
1eJv1y5Y3i8b16Fhzt176upEJpYFIgvZFunQnyOt3loUmdorrmQ0Ezl4zm+/UkZT
smY5ERo1NmbgWBDtW9weA13sMMr3CtBf/zdP23ysLmsoF7Sd8u1omOj3JLgobSNw
+ikL67faTWLduGXYE7upVRdAycTf+BS7H0TDWehuMKGikmkVHk/0z+keozLbU+Jq
gyVroUhX+Ol+MtEZhQPH3/8gIG+rubnXgzuyfI/1VxmpKFG/MNlJ/IPxG7PYTS2u
FnCi+c35Y3J5jy7zPPCuXGMBllAKUNL2yTokwrsuHqnY838O1IrUQoJNaRuKQ6d0
SUs7AU5FhaJ2FKBwZXCKKJdrnI65D83ogHc/enai/DL69V0Kas5QGni50cphNYAA
IGDyhitjvn0XiizY9/G92WQ2OSXQBwvhuzk/3GEK4PoH5JIv18yHIaIYzlCKlN4a
c0FVLNUXTbWPvxu0sabBgxm5iARADuA4zqfOlzJRGI2lL16oQVGEpeIItlC3RPnN
f3YKvHvaX//556+VjT9R52XxLGpUCkeSa7uYMWrTJLK13Z8UVovPXJ9mxBFbULHS
FRddCgZ8BffaqBnY+SFWcQw1AxCrtkY5PmG+jkis4Lg4JG1Uov2vWDPckz1q4Lei
P8q/bDRYAYqRVtqV6z4Iql1CfnSxA0tVdWGyNkpGmrXHdcYDAHuBdkd7tL+SNIyJ
vDVcPEhp2T9NTcA4Aqre3/T43/DrUfS8PoYRT9ghlYOhAf1dQsRNnUD4jq5bGSBW
drvTfyr14+Rz7RuvlBGotxREDnTLiQMSns0aOtnqfPBNnBOd/TJrcP3OjF5u2Gd6
EDegfIkzZxLSSVKbGpHEZybVnz1Uz5uCcgq9KqWoEPwYdzufD+o9nNafDM/hf5mg
fgL4dIVbZD2dey5BtnDH418veFi0VY11o/B0o4EJnUapukerDm6Gc7NQt2M9SM0E
b0hjn3JtovE+XAeLzx0c9wLhtL53R9eCmvSzMYD6WGqFWsonazqfEDc5d9Js3GBS
j7W6tP1o7ugC0texfd3zeF4h3IV1mc73zaiwvnVqeYMDt1XX/X4Cp+gt2WPtvjeR
2mAKuJjHRmYiiCdCCNudSNmUyfHOrptQIE1Ge1hsToGfikX7WBOoTZ8n8HgqGo1F
QocHOKRENsbKGpFMoN3tfcWFVCYpE/Yqbcm5p2gAWNg5y+7zL6qgJS+tPxCeR83L
ACslO6IwOKmEd2PizOO29Sj4XKPfjzccWUP/TT47ldBs6m2fMVAkLIACOAT1Bi1K
VMThAf9uyHnWW7TsEKRwFRzUSPc0Io4+7CLjWpopAGjZKvypAcgyhpva5x6FU5SD
G0pGdD7ejuknV75RODlrGBMfG7meHRHKQkvgKGpncUUTBQRSi+/9SBEybfmvMIoZ
q7E1TJnddRzMa0YdVyTCrrC+UdPOj/h8x3hVLE4hZbdzDN7FeFGmZvEyCnmSApmG
pj5ihuZFAMKfkN90LK9NQtw7Zsfef9iJ8pxSHx3crCk/JV0wAM8MGlFpI2p4PBDC
ZFsk7vqVDS7hweoLOYLNWri8GcAKMWUMX40UavP2ofnk8B06TRbXMxcWF3w6G5NR
d2FqQqJGwAB4qbCbn4fxwpo6EZw3903HKmSZuVqe3wuTnLk2J87glzqQZ8nhjruc
MpjWk5SbMGUjvaiY57j2kmNN/I7IWYdBj1V8FApEd56rZEMC0lh4GAgWblH8bBOi
7ugrBEepq59xsHshojYMoqTp6ZP1C08h3hxPAV0Hlq0FfKabxie2jcoiJdT6H0KG
+PQXhjVzKPuNbUpDGXqGjtzGB8TCEYXPjAlSo0zvphSK8qTJT1f2naBVOEY9W/l7
o2YnXAhSGJ1EM/TSiiurl6nlY+tIj4J93zqCzwLNjgLgRpXP7c3tJpEGqoT7xf0G
m+LR1m2A2B5oscu/Ia3n8yH9a5edBS9tEZzZ0EyB/daDSYNb7zqDK5nlscjur/Jo
qLDpHcG/EUnvugU47QDGdStvg5HG0H3mfceHV/8WJbuZOG7sZWKyBwDT7n3XeCi6
xrkS3gaTeW7cV/ofKSP01XeIksFkIYElRR7KormIjhwwVxvW6kD/9YJZFL0qmvWF
L284GHZBspHI7x94GEqw1QOVfabK2HyHILqR0MGO5hXyQ7NGhF6ynTrNx65I/xCE
3kDYl9+ES4KmGaNbJtZkCWeGJHXG1Au2HF3odhrAe2QPSipQm6CzI0mK456pWxMT
t0wqM9VZp5xkaEeYJivJkqnqmCRD9/91teFC/0Crpl3hxOWEod9pDPjsjCleq2Rt
uWlrboRCYFbwKtaTHi6n76C0Kzu6+mT+MXS3FZ2TOVfzt8EVEGgnLxt53ala/oNs
sr6aZdkf3az4DN8PHd1yUGqbr7DuWo0hWEP7exPrqlrCPVMlgho9ug4cAHI0n6Vi
xnQPdoxJjjKVgHK2ELVm9bdTM7jxeZtdVmOnMkMwOVvlPECisTT8B9PaFPLFmb/c
MDV4S5AXTUY6Y8ghBheX/C+rYuTFIuR+8brN+CCPm1GVgeTX526sbU9JqpMXy1q7
2RqQeRbM4bAImoacE+irpLw+tud9Dyy1N24AO3VTO7hrxBPsKOYS1MUdjhvDYdhY
RJrE0Dt1NsGpkIl3Ome1EWdBgD056QXhfVxBPe6sTMhp3cujolKl+Dm/Lkrduo4L
vYLnIE9ChuksclT2jluCxJf0GPfDmw8w63yhZlcK4wICJxl1kjalss8Pyil5uMQu
xdjjXauAPS/JVUe+2wsconLN2T72/+HIFSNmxosXe24r9fcY7vK8++s8U3njhIBj
b+IrOY/aQatwXRBFRWTXO2nI1/VqsE9nLs5oqVy2uxYo1x8dJaZG4yb2jXynOoF8
6jxn+Hdwp8sdus+ob9r7nac9kjz1BWZkby2mWN3Pg37FN7E2kGE/oIjezCc/nPF3
M4LY0sH8e5+uZ27TPj5JICP1OWZZhnIN5QXqSSVkcDZ9j60DwLiWRehB2XS4triu
A0l/R+zN3xh6yqb1HXhSwwtJciCc0Sfj8l4hRjHvzKgEj/mybCXlHOnTMfCvMy/f
Qqyj+BYQPrNDh2yux+1g1icnqMGuOTAaBvkqF+IdvHJCQsWzXb+R+om2H2MMGffH
nkoaCVfI+PtqDKL9wsqLc8Zt0cmStLkrHOTqHRJCP1Z7ZZoHW9MlEN/IBrr0Jxg9
u56t2RHjFSwi4+1gNKXOmv3T0mlIydHLGitlVwOzsBIssppqge3F3jNxAQ6ufo+x
lcuStPMYwgq7jP2Vx6rlUJZWkdGaaBVvcDPhyz36/DJpiiLLjTyiT3PIfhcd7cRX
2z/4eFVopiIiLs9f8i1FTmMr2yCl05TxtiFel2Qs5jaKO/qTSjQYOwKaNT6frLIF
8Sh2+MTWf0RgxTe2ctVymVZhrQg2nDOBFI8lMmGTIyrXH3ROYJI7BBSRDUv8inoT
BpZ0S/eAcyPFq9JcV5XYkjr+F98IAmPsobFnhMfi/axz9YdQA7Dxl5fj3z2NgBT4
JnLX12docrXkMFRMSDsYNfhjAwF0E1J5X9KAUK2qZqN7Jd/d2yb3RLInPdnp45kq
TI6WNB78YSJw40WXilU1fhS47+qCdsBYNDxWnyjI/mE5M35ts75C448qYdNbkAH2
l88TE+0pNQqWEZGGCPDhtkF5Q10Xa0l0jsI/sGFFrmsnY6bTn3Tp+0Fjpm+mUDIZ
3Cz9gu636kb+bgtMMQW0HncPXNBzP5niBaeDAbAyi6JD3GK8FPUIvWHN/G+FnhvC
i7ACtIznLB4jOWzhHOkejBoWrLKU8ch0kQt8AJOdlBi4nfORY8No/o7XNsjzNIXO
G3dU6ONX42dZQ+/KzRmRf03NKx7nV5vDts+ko/5aoc5FnC6b83WXUZFaknc2u/An
nIigqh8SgqYc8CqNIf8HAqiZwDA5km1H2euOZx6+UEXwOM34t2RqKGOXUeIecFqH
jYyxprP34ZSWFjTK//+N9rmwfRhTrIaNdyR/t6brPQa0Suf08CokF2rTaLE+FHgM
bHH7UC50B6Vodkc125CAV8Q5sWUpxAKQm3F1bS8g1VLEoglXPL8dp5GOej72/4tJ
pYPLfQPmB0Lv0navAgcwE53bqve35ZrnQpaTaAGgy99fmJ9JTYWD4cyFcCPvx0ty
FkV4rLVdGPTyXPv+rjN8O8if27KrpWLzPBn6Dw7Op1gAGJKVV2zkIdVAhUotTujS
AcaYV5oyeQZOhVteXAUwLZc4NqxhKrV0d6enIF414RxDuGO/fNbQtHdf6ZfRkV6d
OwNJ2Fwk9L8NCYPFaIWNJdC0TMUCTmU5zEU8+P71uMaooF1o6K5EXM6Pw0smxIDB
JlbNrIqiySkydPOBIWyQ6G0OPDuCtVT1yquz7munwbmlyDp8xG8PX3L+m57WtwQM
KwrT06QTfSAvbFXLfRReqodHwyIbhd8jfoA9ZIVOViOF2UNd/czINUQ7sprzeou9
423QIr2292RjuYEeX2zVbhossJFKk+No0hdWJU+wwOF6KNTO9c49vDZKOwKsW32i
naflFOgOVzmQpztoPFQoNvEGui4PVgSYM5xZusADX7+uSff52VMGQ88FAagYbXi1
9TWfARj/nNQItiHJdHHTQCSIIbLPizmFQ+0G7uzadvoFa427OfPapySVZm0WoKZ8
377+n2ehVdeGrAgHh0m2EY3fpn435IUtMmfPBOHQGFPHw9HCMK4vp+8QWaAZe1aN
o0VKbFyOkAr5B+L9TUgzN2bY9dkKcZnCj5kY7fG9hMbpQz9k02T7Iu4tGJrvEIcO
Yvk9C0SGssHwiq6moiyew+FpC8jkbydZTikJjxxY2GV9mImL1HpD1yz8Ggyvqob2
ogc53SECM6ly8XficMV2EOQ21ZvhiNsPxQnDDVABYg/Zv4MYzv5EwZg0y3rGRSw9
0z7DOCyD/4U2UX05DHfAu2G+f58wakS84dgR3ypsbokFKkPnTYZcCUuyZKOm+209
Cj10rBV53avzvqUeCBjpbL7gSnWEz5qPjRdz+YqIuGT/t94C1YxZGmQZIrq7d5/+
Dq9tM96q1tRaQGWwNUdhd3tbUgCHMR+qXIgTTKvZA7qPTdZyPsOOR5Q5cPnQkLkA
6KMjDMX+gmy0F1RyS6bmF/YS9/cmicKtfIYHX3WYrtfqm2N8CnhNGipgllZsuHPF
UpO8J1hJjU7JLsNdDMpvukYq9kx3dHW8F1S2JWHE6l70G4sKQGC7lfWpAczdQheh
qyxGotrAiOUQjZdzAMF5pfW5Mlh4jKYF2RNxFhark7qyHI2CgG5dlQwg1cBnYndW
2P7YLCC3rrpZYKOf30o3od3Twbm9/B5tC+Yu6cxHOoUopMJjn5fzQhgrJe7YR2O0
9w6fELzf9N2WvLb5nmiNfInwsLGPQogEpDVvXjiwqWZmxPKjFkV3Lxq54Gj39LrQ
xA0E6kYdNSlMaFU3/bAF9QH2zh0We+L7D4Yo978WDjLqcXp4r+MBoxm65fVgFa8q
GncaThulwj8alHrNOn/lWlxIjUfkpajG8X8QFl7VQWeIqpya3tGlGOCrrhrghZRl
BhbdI7i/ayv4Zbo+DQkDzSIFbWWAtW4j8ge2GfecnwLq4ha3FM02kas2QMt49NB+
srDPDC7Muw0kqTGGHIGQMDWGBwgXTPzyehsWe4fOxfJKaJvZAzdqtkQeCkz3TfZz
j05PZ7zjVkZWtQFqzzWv7uTBetW014uyORnX+3YTW00eDTkWJWOH/ooyv96VmMbZ
MjlkgvKb2UOgsofFo0LVY9mnhIoSPgFdi9tN5q66bLONKO9qWz0E2EvK0/Gj0Mm+
pSwXnTV9arMNuMrF7YliwHvLz/IHXfGzgOUoy9no1GFga1XAaVn9rHyIW5VAlS2K
3uav2uvLzkqCilY5kr+lV844JVdlX4CPlraZHTVotglwlioZwMmyyIxh0Va6Axic
fBUovdHrzhqAd66EcXohoYP8TlyFNNO4tSWJfmw4RORNbzwFSLJaRXYS9x/OZQ+7
pe2PDIaQHNpSVR+2r/NIzSKMWqC/Rd/j//kZRRtuXVezJn6A1eflrUHDoZ/yBfS1
PeAVCJjBM36Q1483iJnarU5vZ12KGglzOmZd5c8BH0QsSA3NF+Yn8Ej7eQjfrDP+
WT2x3w9Ja7gYKsoXXZqee17DKpGLIsD+J11/8Do4McDafejfJRhrAKjMfO7O8yph
XavxvSjLk0UrIzdTIU1ZwIKr5MxecEfHpm83iKYonkgLiPN7DsrD/Q7ki0adRvCB
NFZ0WG4UIQlOg7cm9b9+KA5vFkm9R9ea0V5QNkSDJjTmcMPlB0wBIDVZtczVsU0u
YHkN9vxgv1cMgl6e1v3VbfodzMmPAQtXuojQNCfJYWIvdiooQ3Dc0RTJ3/WCyjC0
7SoTENAHRRMCYqfVjc5SdQ6T1BLW1JV3y4aOgRol4gonbIGRjDzBzAao+1KMQJig
Bsd6XLN3CjRx2B/36QU1lWE7NaFJ2HW0J8J7ZY8vAMf676HfGaGQNapKEELvEb1J
GBJHjV9it06orc6L9QjwBDVDHaUzxQRE7Cy+R5Fnn11tpTF8ZB+M9ujvIJRL27ES
1EJZZaPzgkmTLXozrCUQFbvoVN6x/OLeiFLgUH1KgQQA6ICneMehTeFRaWKAi+OF
yOAIE+qMzHkB9ZTnZJQloKtq9vdHDzJr/4Sd2WOZUXZo8NYncO+3QUrqv6bA7p3X
LSfHEziYwk4Gz3C/7RCpi7Uicq0aNZN8QPguWJZ/ZrCuGX4cs66+HMx+2GKWkwnb
I+I9/0z6pdlykVjNPhOHvg9iRTkHofQEXjV0uyB8sxrO/DMqc265kxhNRc5oUh6Z
m8NoWwaFmaw03Aq0GlE+u3qWZjptevWsROD1CAAgI3qZ9J3UhPcjEHQt+7B1Ld4Q
Xfdt7+L1I9fvPCLsfYwBQIk8MiEUW/ybZ5+QMOILpJd5r4jYwUW0RzHax9KiIoQE
tsxLyZqamL9I8SKPUtQ2NRFNTEUFz/XHEcsISb/0+/rtzvqNdC1XZvX51sV1r9Uw
SXw0lvgjdTih4RT2tWRHQhJ3Buw66s/mYd3e6WA3qGtWvCiqnVRp9HOeLh9/t8W0
uMT2gJMEfv6pvftbXKc5KThbVSOPwsvUFzaL6Eh+/00SD/UWek0wI20Du7/lT71f
e1hE03x6h/kcxHnt/Ox8FODR50+Ds1PbCuoqzVPo/Uz8U4bQwwBX+YoHw5reUt++
+Ru0vTYU9MHMVKzkJA/2YaijuOrAwoDQe7HUUpjB9vyXFMTq6XmiUWZXn2kydkiA
w7Mku8gtDFjy1aXQZ4myUrSDsSGzTaRsvMzgwGJLA7e9w5FdQCVyYWMEjUC7qc5W
X6hNlR40AprJVbhjHH8k+RZhCga4X5p1ql5NWfOe4vPtgaVAHQvYKZ/tckYg3mxp
HLGx3aAcy2n9yZNBfu3k1miybwCkq9Nd/i9q0ZcvBUc724TEdftHAOPZSbAcfXBv
EOez6CgrB5lYguiXcwLvKHcZ+pnpviTmPph8SXanXVBK5fGPW1sPrNlMabl1mIR/
YG8unklvWgcrFjBcVbFDPfrg6VgqiK3Ke8ro+Ez4/RJufJ1XIGsRE8YBpGjdXQln
sp1hL4fl11UYGnISiZ1Zinb6OHvaQJwfbbYk8id+Eiht66by1N37BamxaZAz7bOG
95zyb6c9UyVZlRBKsY4Q41uFjB4m5kvtnldAR8z41GhRwkfgTkLl9XvR34DA5/eU
qMFAP5KlmTrFVrOawh3CcveWKUbmXS/LBAT/A4xEe0NswKRICNUPgC2je8EvdYP8
6ya0CmTpbEzY3m6GslftLz9YQpbAFv5a0c/lT8AzMMGNkhBfkOgwkRjsYk+djxmo
aAyxSxfwdvtu2TNt6jjqJsmPCwDbPJYUTuyOrKLK/aSwwUliuB+6QVr4a3a8Q3dU
8iGHeTOwXV/ytEmeBp9M1BHJ9blkRfh22pGv0fEvgYYwZ5kTTSXaAywiUuGzLa7N
mk015ktMoA+Yk/PqefQuhan5rJr/BWm+QxrMr80+0J4SGobzv+zc2BG2FhJfDk7D
i49itURxUkytqO0IGWr3Y0/8vVebbi6K1nbYnuUCRqtQLtjSpjX3lh4/kPQKxkCP
a0GUXZSp7x4qx9W6cqPgNR+PW2lFGjABHUPlP94m5C7zKRtoCnBArr+E1d7dSo4e
HGE04cxUqAqJMLqAXXcnIlayGx72AWc9Im9pfWINO5DAbkWJqIWrrtaY9LP+D+lZ
YG1EP9wIKKk8wHPpUimXqdV35wQtoe+HOwVyfPC7NyUsZOYH/3kXz3LlIv5Yesaz
6pFd/6NNnrK/wLJk9JbTP+oDDcOTC46hpDxnHm89mwooSR8aMpjDt/k6DO9HFISt
FbXS9770sOBV7cEWldMrK30PRLW9uRCUU6StikGmvf7MQXAU5dNRI64yKT2UXHQs
V5GPjvHwbGgBqlNij4cTGVy3nSLUrQ8z/7b+rI5nMJRBavmMeOivld87Cz8WeP7s
emrHPZJc3uXbYu5wVUsw9Rfp8EYck+gj+o0q82mEljabTI+HZCkj0K/qKWaLUTPo
NLIBoDEvSxvzIgrxvNZ9x1G8YKJOO/WHtGpvb7IuSxHbsqwuA6JkRoLef8Uaee2H
PZ4yq8Z3BKICMjJ72ex5e1xW716ps/Kzjpr56CvLfilYsQ+QuRxbp4FEC8z/7eM7
Uw5OuIHNJdqQ2r8p+NdxUaWLoDBHGSubXmWDP0rXAWvgNevwi0aL1ImLTAfvwD5y
VTCWCC5zRTLaVIfFVX/DQVg8TfKamusdxCBw85vgUUvaWVoNk0Y/XVjO2LzBuxw1
1tVRSE3T91UU8ZCRRLZT2A9iX+p8XRww5vrKPUWKOMQYtRNQCfXVgmK5PwPUGYMq
Z+VTt+hKVPoTauH2RcgBRLi7I+pswZXHMuFUcFsnVTkp5ben9K0CQA8dmGQTJef1
6ettapCGeghEuZbYRXBf6LVg5sAPRoNOvS9h/uTjV6QEQvOh3+9nB7EsYI5V8meC
8+ZeehpT2sYI9sN+M18gPu/q+AD1tdhHsWuc65DyVtHzzeAyZ2djoQ3Ra03VfEz3
y1JlfcFzvwVmQ3iZRem113bT6nGstaJ8GJrHhmNmzk6qGM2wkBDU8iBpVvR0VZo+
lPdYla/TOPWpiw3Pr9KIDjLSGmiQ/tjV+rBtUuiOzEIGgPy2hN1BLX/cjfDjmHZE
eDufqrSSjy7WuyBkfwvSyGEVyJ8qwPBvSQ/UnwQH0aVyzRUHWkwd20v2lzSM5Hg5
NDw81lq3aZTX/xtoq+KpsDQVc5NiDDgPt02XkmBy54cd+zEzS4ABMAfvO6gobFgN
auMM2FTStH3f35Fikuny1Tj2096Ooeh0xPZL3gO6tJXLCrxEZ/BdXUj3VHzGowAu
Lap4BUnAB1s85fDXSx8/BTWqYzmeKJX5whN2rLAThIiB6vqbeXSoifZ6tEb8c19w
u0IKKaP1IUlAdbm0eoeNcECd+o9GmEzxRFqOt+Ok9nNr5JV88Z0iOaiurRXkVcbI
hZzBzbCo6UKHpX4TH3O5eXWYoOAOkmTTB3NTWqnRxU2TSP2c66xoKfwyMVVzsEZI
ZdHsO1SILulHD9utemJwOw6s4EwWOWxLS200D96DxQ5eAo3gcg640J5tIPCdUuRl
B40Ti/vHDA4FXwPECYpiRsphqhFDZgWwyhgEXBPJmw2LgYYHpWpB4BYmy1LSCZIZ
nTeSKXRjkDgHLQj0DIbrQnhoJKtD8RKVwqAclTedI2kVA936akcyHJd6/khLrkB6
80AI4bD4lr2XjAjpiBwA+UVngRvo/gDyYl+h3NEihCyJIMRdKOMT6s94ZfhoEE9X
7yhS6ICRNnAYfy+mckzAs2sMD50BUj2gLXG23GigMBIg+4mZ2hzr1JNPLTH6iuX7
0UcH+VpOmyjP/VIGz26guFRONMrPNLOvqynQnu077Q8rE2EfXE2c4eeHd7ssnSm6
qctNb7+UPbBH9QxcywaQK3Z9HZriAg+s5s5qnmpcCG4DyX6Ro+Hrp5LwpLScnUaR
tI5L9SHYbPu8m+IQMp6VgkuDtii9T6ZAkxQhloNki/h/2cLSID04UTCgowDQj+Wi
PiPzwXhCwiWA15MgwHfANlN+4DCiH2JzUruM3JYsSgrZvZDRnXhrtkFgzFLwp2dQ
a1hHkH8TrX5jlK41q22IiBTu56lK300hXj+jp7jPAJEnFtT6rL1YvabdqDBZXPG0
CpeU5cGwf98CEOxZLlgsskX0S8o4gPeHVnC6uWJbD6T0lBEQJVT2EXoFNNWG6ayL
vMSjHx9BX2sOoCMGgQEeDpI+LN6qBDfTf/o+jgigI0BeLhTAk7foB2Fwcw2IbVpn
G5p0dfVmH0WvIMOEtUWUX8DMvjJspywtsZeRL0PfUsm8iDnj07MyErLIE0vOmfnA
gm3KFXuj++9NocmfD6eEuqjV6HdqDy61tXr7GRr3BdIgswcCqOjS5U9gZs5grntS
in8nc0/F3vnVAgYCvtkYxek4PbSmZ8noz6mqJ6idZEzYtaoVXGy86ux8BcrwhzHG
Ix/369i1ObiQNlZgi4Eeg43s/OveftGE1It9cf9NQINvb6hvAaWtl6FkULhthG/K
V0vWnqsanBLjffw7jwd/5xNoigEZ3UZQjEzEPXXOEeoB17+A4iWOAhdeLe9nnrMp
+nk09iaJSRPOFX5AnzLZv4nd54ohtzQZImE5STTw+lciVgR6vdUSxmhO/oVf9Pw7
qcOIiWFe1maxv8HxHnFUITPDCIeHRnjD5CydlURsoq1kSKVG88ApJr7kVtsnrG5W
OyEr0O/nAhnRh3LKsJJ1fge0eicXz1UjtVMqs8F+VxOFoVMRhQVWSMT1gNzwQ0dV
mGKlkm2hRT4oollbaEIhp13iQDT0ikg+t58lAPHi+Hbsw8sfVHHvo0///71T6WIi
cMFaovmf0DSECmFI5+iPr+0H0GIdPTg43Vw7EY7JX4YelnjenTEpq6tg41VvhJcr
pH4iPVYiq06T3iduainFfci44jM3hmmRbhwqRWbM1POjF+TBl7o5gvEOpP/uVHO0
pHg8uy8T4pvXRV2wDe2OtRbYPzwUKk9uh31d3SAg34Cs6fU3gNSkPppEp807emYE
3rvNp3AhoezSjdv+ZiCTHMW2G6TVHUuw35mpy6JL97YApi4OxzZeNwn51e+X1Ul+
vIDZh7Dmj4U9PFOhJRbuaDt6Iqe3LlgSRk2cm3yDVU/xGxK1gFBmCFiu65AOAf/e
hVI8b3Vhu43JrjfhFr8eimm9v6Oj6q3QUiO7pEZr68GDMpsoI+1PJnT8PSpEX4QF
BKk7R3nhtMZARXC52PiYz1wiNRHiUCRgtc4IESu9YUDMojZ4tFo/GwCDUkdvY9s9
ck2CAdfIzTZoqPAfNlMozpRPwo7cNagJCIiMIeAYpOgeno+VOvD9IT7eL4mKOiJA
fjriKOiKt9UOvgCc1xEA7MEQaUxSrANijC9CyfAF6xnuFGUO/lzDmKpbO/M+/ujI
BRMdxR5A2DiqRY29SEpSVMbTmuFFRxNogNBnvl/6if/5ECaRSxRnKD5QQln4UX5P
4/72x7zREf2V3yJfZDclBDhquUjVYj6BUHMoBcT+tDYbd2j5QiUDyjxzA9Q4n9M/
RU3SqbebJXISrJrqAN1FlHWQIFwxcV06zdcKJIZ1z1sGJo3sezYC6I7+7bdI5FOQ
DA2pIwaT4bsYAtvwFNGgHNM5O8Hfx75/uWASuFtv71BsjRdblrHklfOjjh/2EOM+
cKByAVEWj3wdU3PZHF7JSetrZE89ZDQpZDDnU3MvQQQIlCsY86lNEMMQPJYN1ZbQ
pPNRzeYfjw+GXaKnH4ie36OcUobH8WrK6DLMT9bLz3ZOn0XvA3Ta4kHm4CXa/d7S
3vefCQoh95LN5EHAUBBIRaHDR7v/Uu9X3gk7F8PtrBEJkAXkNHPDVcFKjjsTcmS/
WSKuDCqpIZP4YJ/ApCWLgqA9mtmx1tT+HUxnYhvg6B+cnIH+7008XMYJaB6jXLjP
6eiCvTTok4j2payumsuegDayUC9kjlUx2gYhPKIBGvhTQqmdscdcJY5x3iZJ9xPk
u16j0HCKYDpY0dk0SLBRIwgcwwVD5HlxhFxfuOpyXodZnXLc1xHW1HWS3xmnKwY7
HWRKXWm/L1BB5zv3HYukXU5Deoj27h6LqOn6hcRF3EsKppzvKkE3f213AHWrahYo
0E0buk18kEqYdhlmNiquSA2l9H/1tTJpsPmfeBcihBA/UrDZAMYD1oNzIh+Xwnx8
XwB0Vu6KTQzZq4IFb4654XPb6XXxA5OiVSsrUS+YmUMUzr7MEAI6BWjStcgPzRJQ
/xiiRmL/79l12RbkBCR2EEfNnEhSP+z56YNOOqO0fDf39gaPaDds2FcSZb5nV8Vw
p/YeQTJkXwyOSqnYyslPL1t128xtbYr2o/bfxReTLNDrcySv4oGX0AT+hRwze+sc
xZ6fT5uU/X4RYJcBkeYgw7oLVgv7yuDup57GsStGeUtyVFib+WYsMAhWqw9Kf83M
EFSo0/BsikIiouidvx5iuh8hpg05k60e51cNdykiqbNTIRrp0heoUxBpANVcmNak
3cqAjpQWBBA6/vwoAYsNpw==
`protect end_protected