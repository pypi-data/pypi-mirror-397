`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzbxWtePNA4xLKWL+TYXD9yiHYeY2y44D+0FuU5Mr33bO
VJb5o3IQY/D5IiWxASuLi/tF75tFglfGFc/0KkXHqaWbLJqiraATQn0NcxqjNOol
rrTY9WkPof0YBDe4efapVa972flG/ldoX+U3xIoK3/uknU95vYMFGi5tJB/QxFQC
BRxY71rWkceHKhkSNojvccSYrVIhjlInNRmWa1CFrknPf69fk3WdZ/a7m9x6yyh0
1RyHTtGX0zekMagi8JYiw3NLxWzzTtmW/jLAfgngNTlEue/LRfYGJ+snuiE+sSyf
M0dBORHZ/qhOI3WWeeh5gAsZOLxhVy8jo7wVwkjyg9sHpzyrYvtnKhLkgCTBBQTi
82qehMB8qtwjwnvUQ71nztzdZUOk1+NfebPUCvCI+yWYtYklgOvflj1Y+9p9PgH7
h157osTR55HSsYwmP4o0TXiMSFw78C2LYbnAqSj61NkuxdWL5Dj911qN1iv4QIPO
zUh/ac6MJicmErBq5qX45mY6PReRlQJXDSnDWxjX5OakLgR5LpGx40mGUe1ShbBZ
dk50NNll1+9CkjS9/VCJjVFyEIAAqWgDcXNq2O+80SdByB7La63Cus/igY6kwftI
0SQF/9rYZPS3c/eYrjvebMqd9BPz0cNHAmlr08XP+mHtQSPSC3OL5qo/ospf0L8f
S+gYiDyjSKpPnx9EhTpfbHPSvg7tX5R8Z7E7JLzKujWV1hQYuIywn/DFWbCKVlYq
KhbZp61G/fquOqz9Ip16XO2Um6BDvYDBlNio5URojpt/q8TgK2npC3PDDCPbcpP0
TWzevJO6Do/U+E43Nay4UtXWoHq5H9sZBobH1aKhIi2Pz9aPP4WQFmz0Wd6Gza3e
FTyJdld1ryQXACZWpSR38kinXIjeRXEsRxO29o9UQoNqRpjNB6luRTY8RKZE28Q4
ygpbe4hSXLONr9l+n2k8dQVWObEBq9z63awVuwohn/mL2AkGQEjxeaOWOwEjwoht
jMScLY3jN0Msi0Poxu7LkfUu9V64+GDaft6e8g5/hVxUvqkLG9iEKx8m82u1yLM2
1RkpLXdlAFEppA0DVhEe3zmp6Vyz8OZvt8YZxud1PhQLoE4BIl6xZy/AwiTDrPRB
YzF2RWQpAWWseKaHm2yDt09Bgyse2gqWEWn1l7H56F0pUfUQA/+j07FspCtFhBkT
4VXBiDMqlpko4JdfX+eS6q77Az7ImgZdizfEtSINQP+gHz4L7lXwHmQMylLe2vlZ
yEU8RldBUYXuD1+qnPURJgcHDl8IITswweuroB9lMeuhEhzhz0WtKy7uq7XBFJXo
bipoIDmlui/DnArzlGV2KMDQC5NROGqNjQrrQU03W7ZG/daOLHq3bTjtiz7/r0yR
d9aS4iBcxweME6SQRLIIBtfwP3QIHPETLPMz8O/eQcZnqVFkj6Xe5n4a4CvwYIjj
O/RA6mLPXODnqFb9D4N5AuFLxVEBgdbY04DvPAvXru8kw+4mOtRAD34eZL1T37hV
bp/ZSflss3ZmygkpkoFn9kALM/NAsvFRYqJPqWR2rGI62bm772i9M0ri9gV9qOhw
xevP2OkDKjMlak/Y4ffVCB6G+o/oviYZEelYxQnyx6E4ZYZ8xWj5bTRyWOmBH/xC
Z6I00yovckz+dSRYRd9Qm4wDOG/zM0HhW03Bcpw7fsH7XWqqgFtyeErCgswSC3lV
78nWPHtfjtuO80QwSnB7VsqQ8mDUiRFDQhWdb4gOG/pZUuln9aLmjZc0B0KoF2ba
65hCzMuGw/4ebp+ldCYUkGONhYe3Ju0Tn66GQPxsHKt+irwDzEQwoo/ixRRni44A
+llTo/ah5psjElqiPLgwQY9vmsyXm8VU/xxVvpStsMrE5MQl0zucCWF8Nan24pxg
howV+xUmsHWkfsr5ZmxgjZJWB8WfSle6+CzZUhLwrXMTiPidP4SdRZoBVPGX+avH
W4Ppy7z6bwIly0hxgly42sZ2xMUeO2ByIIy4SMyC+KAsVKK5pisRDOMZIC8Pxy8S
2HCzJt65hz/I+dPXb1gfeZ/Y60zgBOFp2ZjtGH+Y6hkziPUfGdNUPE955LLZ0say
3naQg0PpRm6VbUKi2jAlawBmdyaYFWw3iN/LDHvhpVKKWuAUyYXZOwbMERZJdMIt
OzSj77XL4/KJP/K78Gq1fUU1jflziKQNfzfRo29VHR5E+O9E+cYKfz63Ek7hJYk3
xgNiQvtlBa0THW3X7TkGF0GcLA2DxYzWrxgegAPZxvym+hOlnz0fEk5QsM6xKDFh
dTfoSRakId0VaNEQmdZJqe1Dvh6QGqE5G+h6OnJyWUpC+axSdSSdkHujnLsLg4Tt
/rL5eWypFrgQNIDKZ0zqzwd0m8w9AGXG/i33hPpIL4/FUHKE1GEdb3wjwp61aa+S
MltiQxHzQVONVersJRScn8mTSIo/k/c2iuk1ClpQw+g8fcuz/BYty9VkITkG1uPt
vkbhovksSlV1ar6bx4IJpxBuLhRtzztbmXE2HRpN8Zn9f0zDk9LWFE5ETmF9JN+I
KdiWac+8d0eopdMXFYYOj/Nn5tKzNiiL4byLvxH2QurWeakcAV7I/inLWF4hkHNb
RCnV0fllS63u+PfsDvkCGPzmxwgkcdt7AhMH9OCyyN9xiZ0rXnb0N3x7KVcEZkDD
RHs/wpJqUOE91YJDAR/fhmY5Z2NvOfAUzh6MMeVT4mMhnFiKe59tkgMS8qeGHRxr
gBK1BDYlais1gMspWeDscYxPTRnQKHGe0uoExR6O/iyiM4/ZHOxNmPhwRd9+hT+o
uu2r/4vJPdeRrKFhrh9LOIxtqCyshkagNNFpPa5HqnfpNvCKJ3k2qRLlcPp7CIzF
ATKbA+3+pUoJTko0N/Yj0wdlp8356rXq+k0lQ64eH2noYPnhU2cfjZVCCJaAotlV
3wG3O08yjg4m2oxoFj+ZtZ1cA73hltoL99upDV4252inWrwA6+cszheNABfW4IRH
U3fa4f7vKt/c2Ey3HySST4/nZgpT1jwfo1Lq4hNEWcih/DwFpuYPVPM9xkkB8D0/
ImZpkaOrBiVbXqiv1/6wl2ipdjvbjmT8n9Jp+80+tW9kmxUfySot86eu0bdmlljR
e1bcUEENFf+3FNDq+ympNyY0Lyph6QupV07OoQULhPbZCsGPJbWWv/k+wE4q2QDf
aum5Ic0yJc7j9RESRk1eF3TytlSFcjXL0b+Z/0iduTAYvNf/RYUvWLlR1Gmbe8i2
XXyxwddwhRnzgpUajkom9JbVLsIEpC7jvygQoKH75rp1fPjwivPVbw8kWqqhKbp1
3K76l1xz+ssTKBtYGN0WiL/EHNhmLCcJqaN4VbcGXeMZkLJMsdqaAbSYqVW7e6ZW
S5tn7tAZS9oLNsE17w8jYAXB5AzqXQc/UAUCHb4AaTGNw5j78t0zKUY6AZerKqks
3/EkDfa4s1mEdKp4MdAogG4tJf+w7Mn/HHV1MAu+14zV8SnixPVxYZJWpGtdyhSp
f3jC8g4OZpDVX2x2Elm+mIq4EjcIKMvwfRtzk9YuBTiR21dvjubavVsXfUBHhfz1
bpmRcgHqEYabd96h4ELwDpZbr9Pf0pjKCLeANiXg5Nl4XnEzGA1c8BkAXN8w4Hy8
eZQlzKIR7X7UJsScjO3LYeVqgPteMWII38FJAG3sejT3YIr90VLAfxVTYhuqJVs4
ABlpchL2C7ITPnb1Y9ubGv7HL/6N1tWqDNrbU/lQkqPF5WmuvldnPMRI81X1JNAg
qiPmCIZStp8I4q4pLPsGdZeuLtbGCTK2GRvsAKvKgqXmuBPK5ZzCKQ9qgGqjmm1x
gDwGcFsMSqiZbjpSh2RZ/NRV5jj7dL6LdgPK89C1WcB5+I9Wu8yTNEzFvN5zrH4O
PdHr8JFsEzlJ2zVnwyYdpJQQVX0QDI2iRoo4h9PKV8BcQ4yggnTzGU9D3D9zNc4t
2+J2mKTpz1/NfTEpYqQkGHlv0+Mf3yFVf8qges8Cox/vk5NR3qviBiACs5eQbwSd
foRAYTSAY8oY4L5VpvOW+mknmhMcpkaqi8GJ15K3quU5UUBrTtD76S+61nuaM/6K
HKJBdKcY98BV76ucX9Y+zKXXEbwSES72D553cBU8kTWqNIraPM5DoK4XwHgQc/3n
AP2jW6vptx9GIrACO+Kb3OHBLpBKbPI7Cj5b2mb/w284L9FYWr1IyN42CqthVBHQ
jDqiRQs+nh5MaZKy9Ya2dnfxe7mCFVyI5xlFZmvZfSBgZUMYzBGvELvxpErCQ09O
AvRFQnkzChYGvdefkIQq8udfDFoI9+fAZu+4dQW0LJ2Vp/W6bSu1YQ/m0bpurGST
uE8Wh7eKQ17vjfpq9Xo4PtxIQvk6H4IHVI08oTJeWV0wZ6ZJGlmEjtTiyWFKrS+3
pLIZtP4CDNqNPREGoXaZNokaJzrWFalD5PGkgcjYCiX0vVw4Dhyg2Rk39vNHas+8
CqXz3iiNNLJeIDoc35Z7ohdGLVOOooS1Va0xmDWSf4k3uRZOUxXswe3J6FhhGA5I
g+vSnq9b88lVb61Vm+5dQmKSpmG301psT8Vj41EyPntKjOZr+5nlgxOvJFAUzCRv
uN4DX+9nkMYzHAv34m0WYG3ovbkV80yOQZeZGB0rSZyug7TvGmyu3avdrvr6R3mF
e7OyJ1TloMEffpSpdiykLXZs4rWt05qwC2kTC0oFfLclSzv8qdGaOWxHltfZfvZ3
QcBZROubuw0jGlNm5LC3Jehh74cOl1FhUpkxbMrLgbCkf4cjIO4wcym9lt4qOkux
Rhf2xEMCDk86MUI5uKVnqSN7xj5KvsWYrs9WRafBPHPQBM4NgkDlj6XsT4SwMuDT
y44KR7cee6lVUDekle3tqFGlvKyhv53YvkcRYQcS6Iy/GY91fHT8jMwGqQV+do63
sPbbuUWjifO7bxDmS8yvpvnYWYxZ7NF3Nof+dnYSHMr776F0RecYo+ddKdKTgm+w
Sz0WOw2bPmbIzcq3mR5qZUsLfBcTM4qv9Q7/TjvsTYa3HRnmSvp2iePDjOEEwp9f
oe8q5XzEYxwkm9A4uh5VPE9+i2AqTPRqRZHlCO9jy1JRuY4Ckbda7O0656oSJxbi
qORryChCOoIVuYeTq6p6rK3rS5dZYZf+oY59u41AVma40X08QjUv1fAgSoiVPo2Q
g4ntqG/QVDGsgev/mmWQXnc2iDAfPXGB+h0Y5hVPwh7N6EKySrkXiBGdxXwHxUag
cqJRJmdDaTIJaKrrvjfKnzWS8jqPX6jNJ5126q/1uy1pCn1J9inI921O6wV/VLxh
xZm1WexioIt0TtS1k3r/C5PrPiRD7Lx2ZF/zHNrS5cY/V1n3VcCDB8KE0wIuhQpp
v1E7JWGLPDS0Ij0Se0RzAq+W2t6K3E6P2m8stnY5Af50pb9UWJ2eWKZuQFWba81n
BYEWq+X/tEBkzjVhSxBpRqyj41JkEiWceeVy3ZggD7bWZZ+AIoIHNpCNQ8ZxFxM/
mQT4DJ4FM44SJM524x/G2lRPgUqCrLbUAB1fWxzcoDZ6QvjZf3z4Kh8127qg7wTv
mKC8+CdSK/qahyybLYqubZ1JlA4d8JNiTiDVmK1dcr8Wl8I5B9gnvxKuCiGlHOxi
3N1cZ/mbiCL7qMPueVOajijPztrkDnZbE8Ysr23+G5I5GiG+PZ/zyOzGZSgw1VWx
RdF3fOOaI0VfkPgcrBpVtFtV9p34Wx4vsNfVb/bSJ+XeBON/EWUTIN0sqzWQgG4y
tBfrCc95wiGmaTLLh9M3ZLZh0WQ+RugQpVNFojpVUvw3c9A7LBdWYsLLKskI6d3i
ZCoTbbTLhN9P0OqoCg5qgaf5ye8tzmPyjICXGrBKeD4LgNIavzK3RcqHnaB/Efcc
fEzm79KSE039p2cAdhakLuoCOP0/8OG9JQIjmLcJVxWk7fNjv/KZTTH1qbBSt3TX
7vGv3uxFvXw6T9t7mXKHyUfZpkb+L9aPiA3Wj/teQLaNSj6+bDwP0ovNpmX7LrD0
QSLexVqyEwqIrRk8nPUznGasfJoo0d7+4zegyVKthbOzKioR/u+WfbcxEbRwk9lW
TxqX6pdCA56YfMVXP3TwelLQLza3DXk93qIcfnlAZU92dPzi0bdsxUCYrFGpyXjq
2S+KMInZxWLQBHDiRBsECvGrD8RQS01REnZbLj4iLuihlKhIyJPbXrQrRPQK8dC2
i/evRhsI4T/gm4mxQkfkmKrb5fcd6joQYKcYqwoaHblOidUlktkEC8Z+lKgFXl3G
jAEK2Dya4Dx4bwqwFDxtcewEtNPFvoGuADz7eCqaepAPwQC0rI1W3oLqrUIZv/2e
rxukD1o37Ali4gpSurZDq4xGTVXe3Al5x1V/Fpz19YDUaAfbHqofXkGMPuk+w4o9
jmYfjSnfds7G+U3GpOfXqMFNiQt3NNVP/Pz1MBiwHOcbF97V/8CiO7Eg6k9tQj86
E9IR84fl/n2LppL5lI0HXf2lifZCorzGx0EyiNGa4ITmJhridBz0UxkQKsxZ5OFd
03DhBDz75mPjZGSa/4rczq36PKM77BPI3/tS+KKBFGMKlNH4CCFHrpUGmFW5xvLz
GW1ISAz+k70ofleAfjM2Ntqr6NcjZy3oL5kyAhhebi4PLPUHFaRmLeTLWzaSMcXz
DrxBIPyp0Lk2jzxFrfHFfT1o8PplJhO6/aiANbEhbtva7gzE3AMSU26dFOFJK4OL
SgDR6Djqy9FlB6evtk26oQR+sHfKSiYZ4qP7v+exQx2oNSseECqVEU7ggn3O13Y6
6NtQ5Xq20S75XsiF0rwKxnidirtjRJ8yc4qkZ9JGjH+F4GbRmlyDMGOSeLHCXsXR
mfco34b9eUxFxOYx8+Lgfr3wJrVBbk8uTYoYQk74Cb/WnYmr1GRyY+B5E7LI+/s1
SFADN3wKXeB+5BByjPgpkG+8XFGyicSOkOSBbm4UFphIVrDnJJLQ8ohaIUpO3Ewn
5c9JgpGVIfQ6ODDz9tqSbk5s5xXiEoEkGAGZNHKaAd06Vub5VV9qm8P9+7J/1lvy
u+z7bm+WU/xvEHDMDk56tRtwIOEUrLHb56N+R7xodAGeDlZYnIBZIPv7+zcwYzs/
xYPiyKlgXF3+yA1kFA1UwESApsKBl/XgWIllXA0qI9CvHMs9S5oNZGcexh6EhqWS
4f9szK8pqL4znwkt6rLpxnJ4B4K5ZyZksfQ58hulCGhQwwr+URPD9lg5+vEPuNs7
tzyHYGEQx3CHYyQ6ZvA0fLJDAOZ1cicllGWS1dEaecUKldWNElRcgUI7n566ASAT
cfx0iyiSqI0kEsFKI1hwNjbPsCgpNUUpIniKiX7SHWLf4ZcOPe41NpAtCfOVf4Vb
loOiQHgnw/veZGVA2rU9U7dJyCCVC8TvNydPDrCytvnee8QOPZoOUc0YAkqkCa+K
/b8tzvPN5we8UMzipOzbW/deDvW6CPNWGfKJ7H2AYjvM/JoJIP8sPMa+HHPHc1Xy
KwWshFL3/wH9TgowK531YOToqGaloMjD2iM1xOjh5v5VClQX3U1gu2cJObocH6Gi
v8M7JRVnss+FDOh8jbtHnneSmugxL8ISwzMZfIcqaPLpOgAkKrWDrlNVfU8KC7+Q
X3WAwDq2L+oRTZjbS0lVt3+hRU4t4CFIN9ZQw2Qnqp4Ma4iBOoxHJrHzZ66iAomD
Ns/aXGE9w0+a1EN+G6GiVWJaUZmNzgTKwEqcB+5TTXHx+1JiTmI761U+ZM6l0nvC
qFe0imHgsEgrM/cZ08CzuDIYmEL2Kb1wyqi+vhWqW8uvLWRFCt0xh1rbTBrdSN4G
YtwYDVY+/U1dNOoe21ydkbgxcjV5ldO++n63EioX1NSfnLRg8l9kWdfPqdCJMmpg
aC54K8Q3SqiXa5QZNAM7n0Ilw7p1ISnFLUUQiJuwTGmLind/9hQOHJUYNiziOPEU
CPedHltkL1tVCPsllXSYYAS9LE+jrrgwA7NJi/+86PsSFJkoUxkAvEikObEtCmqB
oruJfaNtizL5nzGZufJ9IjkI1mkLmJtJJqGDio/Pe9AlVpqp4xvG/hVzDbYp2oHo
POvlZT14+2KD24YNzj1qwLCH7iscEK+5cPC1r6UtccdTIEHYDtI4T7ZTxj9Andpq
H7LDyaywULvIr6/W2FTWELlMY3HGx54tpLu682Rl5pmUXbs1MPXqdFejs5DyYe8B
UFk96xeySXhOBua8XYK8w4qMXHo1YGaeob1zO+gscNza5c7ny/GvktfPNWRitC2a
3bgIe3X5415aBJcH0TeNNKjM/ZH1gBlYTDP7e9qg2EbbdL+Qj5W++bH0QCFEqH1h
W0HDISbqDuiKM9wam2XKyHn8B/iYtB982h9uvYFEyUM06A8omIPHlKRQpQoEbvIH
MyNIcYocHrl8mqLu6Mc7Bw+teX1llb5B0qipEojW/VoUmpIzdm/TSUlz9mu1/Luy
SFeRQLcFaGdw1bgzxL7WYMcOEuO7gHW8Ie9w24E66qpVLzppgbTbbjZ3Z2K2s2Yw
9Y3FZ5V2tdRZdwOJOi009cDtjIA+O424jd06z0qYnOa3NwmzCp2awXdk8uViyNUo
QdgTFe75ZVt358JSRUpq46PqSN9zJdiX6XZAUHfFSSXYUAuOIqGCmD264VBfjlFB
5yO7NPZiu7d74M2U5hwz7aTBuc+KrWBeotC6jIt+nYVHSSUX08SIdzt6giqfszS0
gHV1mmmL7F1j2sQ3+B4n52RYb7AmbN5yK+ukVRqQXzwDH93daqnsFmS0EqkjQZvg
BEFFKdgJec9uHbUj9aj62nOT/+jVGt/Ct+Vj0h0KtW6PDH1gRVMmYAJWwX9tiDze
C8OM47xwRPvGHayAj/9GUwzc1S9YK+OW3OK0xCV62I8QfmX5ZyZMOASocX1OwzEP
wYF/TATC6QaYTm+iLPRmNf3Wky+sgyBD9POq1gYWBXU4V8fsvgUKXfFA6A6Bgqyx
O6r9ceKr5MX5m17c/QhVNheYqAky03Y0ixODIexPtqKgQDPi+kMiSi4RNkDPY1Ik
IEydZE4Ao9or+Rp5PvVPWNOJfSVWhxqcVd5QXQekSBcP9FC0hJEyU/j3PXmynTyC
FUNTxzBR4aBHexUhKQBIQlYXn46FODB6TvX1A1rmz7Y85QtF4mIwWxO3bAV7YRqZ
R9XcrdLs86/oRwadFtLLVf8MOUVLsRTW6Hey0m8BjLM1owtx+utZKlG50fe1SB2G
OA3unLz2a8Y33ukkgiBbolgW8B+Q+bjZINNgEIjA9j1RqitxAdURsYcgF3gW5gPV
Bk7jUAe6n82+0YGjq4+VrHD7UNu/XTbIz0ceDGAtzA9sgj3I8KzuWtTKhbSBas5M
f3OUFJS7ClYTJ0a7b2oDR8HvAVoJu7JMX/6WVoMFznmx21FYIjTm2mLrpnjCGjOf
AeWrH5joKwUWsq8o10Nem2KNiaaUostZJDxS/cXT8X8VnJshN4p0kng+d8+WiUir
rn0t2glYJi6pRf4UT/P5/HjxuM0H1FctXXE6c9itPotfNgoAzlHZBF9tMtjOstqs
kAcQQeakl2+QB1/ldaqZTctymSPL4FSRilSKkN8FiwwmL9e3zp22GyRlgV27Ff2z
eWSYbutOYv/vnXZW4/hWBGRB550B18uLk39VbzcB4mGDhs/WKZMiHgvpP3dhXfO/
CFcDFoOFNQWmCDS/kqwXsIWtDAt96pa1Wp4ltfwAswy+AMgkPok4AxrqwjZiBg1J
c7IddQqvoshnXqBYEJ12NNEwX7bWPCjfN7Pc2HtysnsbMEGV+35jdMzu3toMiUCk
KqqZntjCUxZ2/kH8Ww0LmFr5/v4fN00ueNLx0qYYi0E2ux1i8ndADYst1ZSVgZZv
lboKiN8SbGbHcGxAqZtaKwQK7F+IvSGzEmy9EHp4UPTPvuGZSx/jCmIFj/UWxuy2
UdalpODQMqqNg573ANbzMacHdOWRUP0jCl8rG7ZxsTecrCbbaS4E3B3iFCflC1Pv
tucDagnb7VzQj2uDIP6D3lw9Jg4MI9kN8ecXuMNS8ZmvNaHt+bxd2REipldzkkkm
xMTnDKLeFrntiMK2cH4C2z+2gNOsuyCwKZ/0IFN0GMqePY0NSaE/5HzVhgMSw6iX
joDTtAGEFvmq+LB6Wk3cWkls8pfDG8k5+onQ42FQz+uFVyG3B8rSYA3ostpeC5fK
00A/hvZUcv/3lnfVgqjXbOqahCPaRReczpZciGLk7RSXViLlMea9Tq1nf72Pt5US
P3im3KTqMDknOSM6p3pvNy8WjLsi1wriaEDOUxNUrXO0KrWywLnQyyzS/4ZxaIuh
j5MpdQELR8FsEfluuQEeyDMkbbr+h6zXNAiDJA9an5WgFUbSsjl4oev4XW5Ko7E0
1putUw9czW2qL6V+wvhEs+M3TpYXITkMoAB5H7Wq+/2uVSjH1aNOheQ0iNGI4I0C
ld4+R9NbT/LVuxrvuhwHQIvSJOlmnoei6Y3mMVvKKvKwVEDe8yt3VJHlP0n+9nNm
sR15ixh/8SRjpdFjQ6exAmsmbHsudhfeQWwJc7/cydYDtr8coTnA8dYY6uywovTB
NJf0JHTtUOtIOBpkpo8OR3x7ywsawUjCNrSacdnILDgygeFEwbO3VhHWwL+jTy4A
lKG/hjw3vaf4tur2/0/ySDWzj2ik1adG0bs9pPpnQmbmH2+3QatUBN7wwEbHkc4W
NKOTOxQHslkgzPHd5LOIFCV4hzGy6IQ7tqjbqssL+fpYQVFjluGu3LQFeKibc+W6
EsnVOAGM3n9V8ShEMl2iTI+mpMlRZu8v0t7I8e0axZiK1v9g8Xv5MTduLoGbOnGQ
+IpBGiJT07F94wNzaDVD45BW5jIrv3iUFObG02yquIVq9VfDEIVg9pdjc0Hk0XzR
se5Xhme/6el+YqMgbJ+dVyqf9sS07OE6tqdiakSbRwxQ9UTC3I7sAW2UpAy7sIw+
HuUVSQ5k8pr2pLHuZQLY7nlmk5JIZiliLAN7I6uxlW7uNRmwgowmmKui11LRbVsf
Kq2eF+tMHWN505Z87y7Km8C9cMohwC5YdjM20f2c5tkscSYxtsZnnzqrY5vkcZBg
sTj2w1NkbTZGaKREnDDvohdjVhB/+qv8BFnFro7MuXqkLTzg+41EcPGeRrZKA8BN
j55o+16HiHS93Ux5g9h32qdCX6eVVp2ujD8ulSoNOtFnElsorZl3RjNEA8mxqQtC
KGC6FbhoTIIPeE82UuoLjVtt58P+nB+doYhF2VMr8wSe2p2f+yfsfXwtlQbV8Uis
kSkun9zVez3TWDz0DwFGeF9cQ2TtAFehY1jc9/5RepPbvaICQyHpCs8iTZhh8xYk
1zJjxKe8AO2oM+I230RFXoIfqr8SWz3d9r19go9b+uJqgrHYtu1qlRRkVUXWaMzB
E7DeLQUvQLxbIBCi8/pMrNn354eoLBtlL0ZUMDuJklVzrkqXht0MzkkVulyqJ6mF
lgeZXXw5nE7rgLjHk6mNQcznrXpUENFmnQ8vLL0X+G+Q4Kr5jt9F5Jemrr0aO7zv
Dc/nNQz+e8WUGpBiFYcLvtl/tie3ZAHlOLtwwxLM/3Kj3caZcw3qVNSZLgmBXPTi
pVdu4kwkwCO1JhDmaPO26lnLmtCCDhpGgfCfjAWROasSntx3bler3chKhRDiGdQB
zKaWgV9LVn0OZXOr8eCNDrVN+Fj52/qQAFIR1W+RvLcugteRWTk+n1VCBAPDMbyr
6VSW8dDlV++DVAW0S/FaKEuW+HkTyjyl3YfsuUii/cKtAJ2EVjIF2u3LgeDMqCHc
o92MXwVKgYXHfHHt265DnQ3u4/pvnX47b1HtwU8q4PK4aymokwrc5/PoJiZUt3am
5Q39MZd1vkc9AFixCUvzNHPL9numW3cwA61vwqIvlEhu87A92HsvCL/O3LzTzctL
PbMlORA8ov9GnUUABUbyUkjqr+gOJBN2Qmxh6EBYzyp8o+8N1DpQ+YpuP++9EqNx
y3XsjOT6cZSqKbXa74u1cj0qBUJl4hHX009zjzUu56Mk9v+ytOYLCQs79aAys0Qf
rEZX9FkR2T+kZT0D/FqQsEbSj5zEeE6yFCuGYSCRNg3p8R2zbcZnVU23FxZeaUGX
9GIIUMzscUi141idLKnKAZqwkvqdwbNghH19GMqRj+U4SN4HtU8TwY9twZwzcyPB
LXteZvQLgstc3RH2MqZvE0swQqrHZx+EgQVYAlwzF7cFPx9gN4AsAQq+vnSM8U4o
sEMt8xP6rRirz0fbuTw2tdDFAxlF31wfWAMIjOtan2MTo4n/qJb8iKuwCH4tdxD0
ynTAFvPT95gp4Hwv2CEusXybPOEsdAcQfPAhwQ+uDcwwIi7/z2I6cea0YtqId2sg
h+HWPmjrP+YInWq0WhYE6cRKf668e8/EE3zwEqc/RePmxdj0H+uO7U3Inag3t0EB
FzXCN1ofZOgAQRhCFyCa2SOIwZaKgUBDjvhKcZ3pUWzw7aOEX8Hd02cJNVHox64U
KU8oFKiKlpiqfqYJPZDJTLPpGDPTt68VpCjfWs0tPsRadQ85txjxeRJTWp58uh2W
uoN4kLrXd5vkUTbHRDx9M3p+AACACoaUyNobb7eZ6QRuiQ94u9wq9Vo/ZcORqT90
Gifu4W2OIgFW9YTQeZJMy8yk86UzTsZNA0ub7AHFDwxcGbDlj0MvNkv6bqI3tAzh
UMpnYAANOrXdCzCUKxAHCqia+F39Rhl1kXDiwgE+rDgSESz8+HnpF89O+jcVQb0l
BeVXvZNNfSq6EsO3/TGgtweLKHRE9nPNxCzhRWR6pt5TWkCWTVtpvtm7Pz+Rk0Jg
isPssInaCzawDsiYhJvayxAh1dU/28qpWfdc5R6MkgiiuPa0UrsIP+CJc3rMZ6Gn
iqB6MISPiDY+Va0WnF3A4Lx8GipRsRPeXiVkalMCXtiJgVxyoezGX5e5AC2DpRA4
w1efUOz7/cC9BZX05c0lf7qM4kZ3UvkOZ/vSRS3E4KdU1jn4yo8f3Uyk9ZbTNijJ
GI99MXrkAzFlI1Pv8rb0s/HV8wDZkdXj9G8x9errJS/ff37ZQeb6Lw4hqmGfW1Xn
0BeUmCE6rwGYCd7IHSPmcVayRUmYJNGY9qG1PiMe7obcb93Kj05wwpHDnxENTEVY
zwZCiiRUMASkwzjLImd49RvbAoOHSt3qLiZGgOzltR5X0uEScLJ65vZ2kuCFPrWV
rr3MwDEExQRTHEZznVtWlKwMp7L+fs7BT35KxXBtJ3Itf3PRVF6qNgwh5qNBkONK
cFh7Q5BZq+p+eKF34rtTcxYmzutqoicFxLIt30dUNSnpb9zfe+ZNaCPXFMRhlYHM
QgTb0PCjNLLLAOxD5tzGM8Pz3jlXPr5y8/cN3yEGb0BHSSMPLkDSf11oI3W+i7ub
gXffpBeJXlS2tSJx9UT23/OF4AnLJzbSkNPUklpzyv7iH3KaEXjxkfuZJlXuNT2g
JJx9NxH5xbGlZCJbI1cuNTduh8s6dAp/fn5Z+FSECKT04SgtnocC8mnpNzs5jsUq
Jo2dmQbusH4+X5unQxhep81NGladlR3LI3+ztrdWhKh93eleu2npOt/FEpRpmMwY
UDOBhrP9JXnfWbgvOEOAi5Lm7dCRiwKkmpY8/0sN1thaBIVHo8hK6gY0PtHWSXtv
PpB7K1xu/KsYjnnmxF14kxBOCORjMzwY8gf8uLONjnwS4HetdbO+bD+4pdUEx1QJ
qx3VgMSaJt/XWAiZf+9EPpYYx8AJP+la6DeFP2E1GkAwsak6fPm/FQn4ZyOdfMhB
L78+r1waGBaTa+xFtFzuXqBRyRvQpc7d+u7RkVulqVL+JbH9SG50HLnvZ7fDRRCi
oWt/lKMJ3x0BsYdX7tVmkE7zrlnB5M1WnhGWXGEW/LK48Oi9GySJtLkFrDa5sbq5
sdGRrWIEHjP1oYVB0/3hW6JbRsR9j/JiP5C9bg39pDqJmdfa9YZMVm5vM5luCa4O
DpDRreqg8n4rzIBmHmEgfDsyLdY4nfzTZXKbL2gywkufw6dLa3PQqF2djpenk1MV
THC1iaXB6B/y2su7dIUqIO2fk2UEkdY1WC9sW4YVcuY9e+xgoj2TAs8nVWE8oVqY
7JsmEk/SBErOVmLe+ohXfJdCJQ1AzpEoDlXA1f1+/NfFhi5t8aM9GK8e9BB/Obhm
8+cHtqluv/RGspm+kZWwGTsPc9HsFIpUUlHvH5kv2B4Gv91p1n4KpP/cv5TaKwsD
pKx59f0wJ8qMlCmOKWNe3HkNWRvQTUFhYE/tny04/BOn8YDR9lAWr6j+YnAAcfTe
UvisANtCo9Dk/uKiWZ0pt0FyBnZ/GcvjacuScnbxewGQqk2q2lpdyW0QCJ7ZK+P0
CGSg7Q7m1M6XcQ1h55OvESHBJJVxKTH9FX3Py37HDiPkfsbp6+kUi6jdvwKv4W5P
GqWj12I24v8pANnAXRT9ZhlX8PE+p2OLkkjXWuZ+MdD1Mzwk8DYvq6X6IHpfZMfg
ZSppUoVGolY4Y5bt6c4B+Qhj7koqPwh3XOsWulpmy8Tr0/CwKPGnLCRcjkDRy2gN
3IcjGvxahsECsD3tohBS6qlq1Qx3dPDhrt/D6nqogMqhP828eXHJ2QTfX5bffFyP
ueO179RTnW3eT2+9jPrEUE7t9atVzdUeVWE9mZCLBZ7WItWxtLVuLNAGAZAp3Izk
r1UE6doIpXThqH+/K5t4uY06w2ZgSUhuptR5Qt3hZZ9gWnJZs8qoxDSptlYmlo71
OIzjj+GD1CHEtv5pQIBy4/DYhB04OAwGBH6y2Zyk+qal2iNbsf/l8F8Gc3NBtmUQ
/igK/+DjhL6/La3q7FgVNHHsRdnoz0yo7CryXUWDOnbGAxaVMZZY1+ss0702GPGx
TrxMFb2QP2orNTYG1aNRNP4U2vhodMpd+cFcjAQThnh4iS/9S3y8NBdp7tYpMB5v
bElNkBtFAh9vgS4kTxwA9tMe6HvuR52N6LW6EFuiptWNhlYCfJKwEEnhD/lLsYWl
B5KuMPkHc+3jp0y6aVJq/MQB/Q0jjHDRR8i+wpfMtkzGUwK3MUF8UjPISebIjLA4
+tg9WY/DMzTdqJaF9Kf+A9yiZ3jtkQPem5WXdLhy5HLtcnKOH159K5FnI5kw7+Z1
dugHNowJcFsigpQmlFZFCziSlxbpGFXgqw+3F9lpYz8RDzb80C/g2KjrT1p4C3eL
KRT3YSSmdLcXAxCdsEzmhlgOax7qczZUM/8ja/ObuE8LRVDfNM9Z3P9p2TfQmEWU
IXdGO/Xd/l9tFoXKR4c9Mp94VgbUA4hy0URwVqs+J6YtfU/h5Sp0izfe93d9dDEh
eVx736rl3XQ+RifJkOdaT8GLUAq9KEmmlF055iUJUeGjrP2vTynMkZccSvsJ1I7W
T+2Wb9tyGDlaoXwuzYT5yCQPj5ajEhbQDAa1pRhU60SMaAuhaqaLWbdyfLf8S3iX
BKullh6xMLFhFCurw7sqnQtFPoPlAGZPZ7iiIRoQkH2SWdY8LJ1tC5Il0NuEmj19
juCUP5xbCCaZ/Zzc844eHLX/azeCjgLKFkoo9iwuaydiEAclngyefvax2vpS0sp+
j/8t8bwvrYhVVvHeYJRHK6I6wHdqvF1YCxKf6gh2GKDYLQMRkoNYA8feVO5ivvp1
Ma/3uygx/CksN1+vGqsZugZMavmatJNoba1L0EbuLQmDsHj1oi1QVb48lmt5fKA9
5FlRaWyMrNDvmcYXHT7ZQF3HXCNrb2go128vfOS/UowV2+YcTokoEaS3zzb9r0wk
hHzNVurzgm2YtgtvoiFcoMvMzSFMEMPLY+XVLm4nHcyTiBnYeImY2MbKwGxdxMFk
h1ux8RSStU40R2InFMpmR360CYr0vXYx5jOSUNbJSfPYpYu9swOj99SHWuSGjmQv
ATYoxWByajinHuswv21rbgUgk4tpDssaW8k+K94AJD99YpH5xf8rkNsg/JwWZmRd
+TrwkL2QZ+hg+UjmG8dMBJ1HZU2zCO5X6e5fdxVRHwcufefo/fyhc1vFj3dUKceb
OH9/CzhjXAw/TeRUvy7R/yafs3+trMi3z905GzASrZNW925VVU4H0ywyStHNRot+
eNiLpXfmEWXGG6nkGTiidLv5Jb1YI5N/KJYIgqbMQ1wln7FMMbjKUuvudjostJir
mjzKVLxYuv17u7N9z14+stTODcKCuJ6BZruSC7KM/9KKD83X7Ms9cr/mYoFBzjcY
MVYY49mBxeOJGlr5nTDZNrbAzq5tsT/VCBz0tdKgKBjcmdVsrIL3ust786X9Hygp
ECOtIHeOKwSiUhAuYyQSq0Wnb1EU4bMEeOkmvjeVW+81UebmG/u0o5UEICnSGhuH
JphoNsL0j+pUwb3LjnEVERMoFc6BHx0lIjBejL75Bg6P4wa9GJOfo5oMqYU45zNh
HAuve6wqyMmsMC/+N7Aywb5RJfMQ1r+lq40EL89E6TdwB8CavNMJ1jnvZADcDhov
V2ZACbzm5edv3gVrenyZJk1lwUbu182jXmbnxmnwUV5IWFr1vlpMnuhEn0RrDQ9m
RF7O0XUgGIhlY+DjqVZPywIGWA2Snpm5QrQe9axomSSgw9G8Tz6Q3QmvSFwabjik
i3PDYZbXM3CN2XXP/DsbDNDgJ4BuIzZ+u5jvGJOTkKZD6cllAuBVjHfP8VSl1rxM
Odn1l667jbbW9f6sqzec3Z0My4fwB/gHLVLSclX6AIhhHjSfHa9aakqKfkKNJgnG
AiB1/wiQn79aXHX4Abr4kHKpQulxfgB4vh8GrRvXsl/a6kid7aFbBkYF5o4pEooY
fdy6psvmJ9M2TDo2ST/EL7ri0MkuVfsLGsVAO9OG9SUJJQYLqMEVlwE1gDa30TXC
I6e9ktyWrGaelRnvzu4e20Aj1UzCkknjUFiVogw0gT0I42ewedcCwoOfZgfz0HIF
JPVhQG3BtmtUyPYBSpw4X8KzQfyi22OjR0N2kTy7gVdw7KvWq+2xFF+Y3reHQgXY
sMh4yjrDpkiuC00AgXjfvxLSBLekGkxILFWMUkocVd+kX1vE8N3+gkroNl1H+VU/
7j2xnnUOx5wEjSCibTD9uSVI9/F5i1QFZVmtmenWqpM/TjutL+6nQ8jkkmX7g0on
+LvrG7jzMYm36qDXfVDpCV67UdkD6ovDX9vOUQtCcinYQWeVuAjexUUecg20REVv
P6fusMe3N9mgDnARCQ2D+7LJLTHesepwpmYE/PI8CYXIQMhhCUWlUeAOiyklgfsi
5adXI0mfqGm5LDhqrpj1YcmhlNxiWQKww/UV+1X/PrsTYQOgRwGT5yMS7E1C2Ewh
RdhZItM8bq44OAGeqZHQ8dYKdMjJRsPoRzx10L2OHpYVDuF7JvjWZYG+gR8ufujl
sk/gnlQnZkbNr9YlhsifYvW/y18I7/GFMlcKKbnnDZuf65MVlv1rjej7isoG3k3N
Aaw9rhp4v48KEAMImiHsTH1QLKX2jqYKYYVMywq4Blk6JNh3Q9HGmwGkJ3mMoQch
TwGV3cicKpGHKvXpyQpEA6Oe/nJwo9ZKCYAZ+zkXzP/M9OQsC6QdMGwfiC6Xrpzm
Ym5QYgWjcNzQ9KgvaplXO4aPzUq4gJr463dxn2WFxsdomBS1zpFSNtdSa30fL9cD
+rPxnAT8a/wMWLySuWLhMuTpoADezAx1Qbvqy0R7FDwNNqomCce6TBSm1v/KvUtL
/5dqi22/qLCjKVuSrFtrVOf8Fjd2zCuEGiBplfKhXArSQUha6GPkeFf5GGiRBysf
iXRbHTBZ1kwoAfqlwgxpENcCN1ps5aP3pcwptTV4WCgMpp7w5INiwaJ6oVN5ArD6
TiFKB0jHLNl0c4O8BNVOWViE2grwQsuJ07xCfi95y42QvXKXvCQ/hHBTe0W4MCuQ
jA4VLrvB5gwlv+Jia9SEbsCKUcZ0+Eg/yDNq8FEVQNm8t18t+aKR+EhXcnNWka5B
63J5VTnY39p6jInZZWiZ41PGhmVFeE4CfvU6B5Z9Px1NC77VJtdJg9CvjR1lQ1Wr
eqkbv4dO5P/+yEOhNpzFubN3KMtZhwFuAiezQts7jPyCwCmRtr7ardp5H0vlxApk
nO2qFxOXphvfy3S+/9jGoZql8bggEB3J6ydR7WPFq2yKwVh8KHoWwvFmXZI3A5CH
+vTIJyxsYTNL0tcQ1IXvOkuwJR6D7BNZa6d2H/SAnc5dmyjQwm4xvxp5znIozeV0
sFT0K9FO9AgTyjWWmSl+IY8RQFX0nikpRUBXUhipS4UC6UWVimpIy0CUE38p1KJ8
wRHeSgOBPGPJ3kXrjYSQ9gXmJla3F82UOeBKDztmeTjsMyoA8JfxmLERIzxh5ofE
RYMjfsqbezgU/8saPvYk/4HauQ62bH33Q/+NGZgL6Edxp/wgKQfClb3eTWiWh83h
ms/5Q4xmUJWz/UxQGqwJ+RsKRzR03R1TN5Xo/gcfOtJlPF2I07EUthNTCzzSueca
tH9r7FRHBwFrgLH0O3AmFKJO8KJQtkUk5qJRDmArT0r302rzRhIcEerj76ckPr+c
sNipJlxfFbNyExhFsZtR58gBJUaLDSiLjLzp/z7HZAzd6M0azpPFVu6lBwboK9+2
t9ZyjobYKg80Q5HIDQ1Cqkv3x3mhiBzQcRxf+0eOezUZ1km3+tpJlA/Rzrq8e5AT
WeuIH9TCOLCgXNpWEyrmkXzv0XR3II5C9GzT4SfycDrqCIeuOoYnLGfXEDj9bNFh
5IUKQg15eYLh9ibmIriL4nSsH7wsvUGmkXor6nNX6nUoAXYitncOl0MjqGMLyjnA
8QSM6XvD+AQPcozUdf7LG3LZpNQr5jlpQgI6A2TzvQZw3srlOYpp7k8+cbTy5y5E
jYie4pwkb8RdgPET/YPm8zQ1i1bQ4ZaxTmfwVCk2ENy8eFHlCNoWdI1US8B1bLWs
gVrx8Q+Ec54c3ySULZwC3IpoAxR74dt4lry/21ODDnLCfCB5nDcyc0vYNRlwmz8I
mLDXoCMx+lY7mWYjGuJQGvR6YkOn+nwaDQ/yNcAW+btjJiCoggjYswJRNThh26Ri
ivKYZU2z2S4u5m0COHAZ+lfRhY7u2OnA6jOWTmNZxzeIdDAxpYjil82xRqjwVAAE
OgQNtffJ5fl0bgqojR0vNBb+cwD0Ft01VRN77gcAm4YHW6ieGA495aHM+DEcUj7/
+PXIbWEjvqh0tlVQhuK3ekfTSN1+CBeDrkEPqYxPq3eTLn/IuTYKDP3IazoY7AQ4
1h+ut13IPWqtnxld6wKBB19cw0Q7aqZomVhsz3s5HoS1Q2GrT+e6+CdT/EqzxQhb
4lkJOA2xtR4JqpRhFy+sAAG64rbrwYQK2EshsYMHjNuwOAubSogccVgE3HEBc2Kf
4QSL9y5ZGjJB4ZZlhJsXTvs/YaTkK0kQF4sVFeHfY43DxIdYI0GVSSt6MwaQDElt
E9g3ij9HXsPdFHW/0WZFOK1p4weSLu9XhINMpw9WVzdf2zBrVqjZV2YlQg812THf
mJVN8qx0pY+qT0FoYpH70N0QMfC5otB0YhF7Pn/OsJyTUoG52QUnpu6VGCxGpnYX
4HJ8VURBsKZV1HiNd8JcjbNTVn3uCgSoMHi4Ujh7jORd5D44JYw/YrO1QY7G8Fp8
Xdr0Y+RK811aBit4erCrb/LWhxmxVEEkxgRkjZ84sTaBOi3cqbqxbPxlEnRVX8T3
g8tfG7Rw+OOSQQGANk+LE4zXEmEQSzViWtKACZhZKjuSI8kSuMqrU2DdhVnOENt0
bDTsbRJKqSHa6txIMdgvG9NroTZUkmFOUVwZJSuNLJbtsFfrgWpgVX7LR3dGpJEq
ayzCxuN87ysgN/Gz6fB+QSvOh//oIen3jvRdU93qwdENFWLBN0kymbOzTz7KcBF5
kF4yLzYs2WCg/A8FuBQQ/JOTEd3nLvuT1V85y+QcsdfPPLUUHzj5np7a7gpGrcYT
IipQ+BIg4YcQSBRonnGt/X20fRt0/hhb4s5qEnAHGaV82jfUY9Jzx9sgNlKeyypk
BZ91uPNhy5pLo0NY6H6z9No5aOTGMULrQMbN0AOnW7OXUbfg11g6fqXAi2fGLJVE
A5JJ9Q0TNKxRrZHye8iH8D/7CNkH7SIPge90JsC8Uhwb1f/6YEpYhsWAwbsrkPBz
m6Gyty8nrlKSKY6vi2Vh1CGmJ0Y7baP7SQ/VQ6rCURpphHE54X2mdmu9e8jzCZ4L
UngUmep7BQvuvbM5mMFmT/Zs8VFjYXcqP85MMsnHSbptCxxaXx+aWfO2pzCMmaN2
m2ncrcDEs7YxCTra80T+4GRbkEm2a/eQgQG/ZY9rD2Ht4SkNq3X4n1w9QIfI6Ty4
0sEDC3wZyDRm2KsqU9B36uuIHFvfuG2rMiOI25fZebcKVUKULmb1EsPoWK3Z4o2Q
UACl+yDB4SJMiDOnQZggiwksZl2YOxh4zGKTcxbes1Q5c1WoJmCZa+88Xh//Dc29
CqWs4rk/waKnh5p5hiVqQuAhE4pHIoH5DZIn071COBjY+Lf9Uz/5aOcQvUwF7K+1
lGv37+sW7afIPwp4VhCOSoVcOQLSrgyTQUDHn9UfE8mplNzQ57JmuCCV+emn/c0o
n255pjg2syr06oQds2UgGQzNCEH4TvHjnxOKIXjC1c3nowvDkXHQkUwzpj4Mpvmh
HzIV+1P4i3MIPSfRecpoh80WIIFIIOnfs/4qLK8MFQAHwtRpA65MNGE1ECl98Y6n
TCEJzSEUlLNZOfU4lVksCgVrEVDvPUL1y3gQGrNVr2Op2fVdzc4uud0FxmFGJgwK
eZA0v0w5Qh6I5vjwwgcC4BLPlxf4x6qQfQi9WNLvlhBLlxMPCPRPZdYCZ/Sv8xCi
nV+5wA8tnjt8ODRxV48muile9hTM+6ttxlDxhnHVxAI71lSnSKZKPiN5s+jMbMqB
AZn2QZzsLTAnS+jJ0TT85ChCIjOZBaXh7yGLPj/bVZlNrJ07n4cOJxHR5mDt+fQ+
SnN1d+g6yXGqTFhql4qzFurTRkj6uTMy5ykNhWW87jXX8iCySyxyqhVe/O4zXyoM
RPMtPj7uZUoYQ+fVZ0oT5PIQYOEx+rKaTWzCvFN1is6JgwpF3jxCIo0KLtKhNHv1
C+oqCvn/9wJw1UC8/9jHSVs6QJwwXcQ05wzvH0E7O/yEjzn+49Bsu6B186jN9NPS
xeL2ZakGC9bhwhWsm1Nv0+yHo3McRPXEzBC3qVwuHD10u3ohlMnSCmiUEGhtN0n6
A6iLbhLA3GXPX12A0R3pwye0LQNVcklbhlh/YhGCM4La3RLa9RgVVazhphwTG7dp
brGn+fMd+V0Qjd06lsFvklhz0+GT/KFHR24gLE1jvLKlufotlue7tMu5d7wuXkFX
8gswQOebgTvDtA5kL5VsPqp9er7fZ/vO4szxicB+N94pFmH5OHVnVHjLcJwBFAe/
nEu258hi0iheZ9Yp40/N9x0+tFBOA5cJFuv1ea7bX3WOKtplb9bjlRMfaK3x4un0
pMuzzQIYox25qVP52rPw5l6pGnIaRflxyCZcUNow10PC3Ecgo4BARM81H4Lf8I0r
Fx5MkPNG5S9xkIOZh9UTiaWlkU6jcryeod6LnEO9fp006/uI8j9cowbSs0i8GsHk
DA9K+zu7yO7wNz9gT/Zt+e/71ZMLypH+4ashBkfBQqiYONHzndeT2pEOsAY33xRD
aA1QzH69Fh+GNzGFwM2YqFmRvhLhYOAfgWdfwm3ewSL1YzVfszcpZMnrjcnZ8q4x
Rwe6k/j/qxgINeIHOHkXDz1zRvUmmNKfBfrR3mgBXRzaZY0ufS0z5W5I83q1sp2L
ryzXy4OnZB4fA8suTpLCFodTrHe33Xe3uoq3gEUsRNhhrSxXMv6ih2hbkYTZyHDK
w7PFIO36cdqKdB6s8w6T1KnhKJHa6ZmAAt6sjV1fEIYzFvrFUIaPowLClCSdhWfs
4yLY4t/gYLuIy97Wy/Mga5uTNafoDi27NLMdE7FUPIjQYnPOffoVkkEC92njcdS7
`protect end_protected