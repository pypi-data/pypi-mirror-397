`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzYWDXkSHoHPtaz3SD2bnYC7oo+LoxXHnIXwrqJYUwMnC
JdMoyVlRdRLVEqoznNy0mQlrfDY6Arbizvu1hY0Q/LRMxvQX678ahZtwvV+1+Se4
WQqsNfRprEypzhmECSr7fnbtsbNpYLNWP4QYIkLKnzekeNX1lMsLUtuXWJWx1jUJ
GBaDoQURR/Td+mNBUihk182Zj9/RmUAwLUe1eWiDjGK7gkiktdujfOCgx4YW1IGf
iOM1UCPxbFBU08/uO2xP/RPHQn4XwqFKOofNMSUTcB1RAm4aDZfxK4ldd05UiSHs
6UkRvwCn0XrSOVCCd+fNximwL7JogrcfZtWCKpKbGdmOT5HM8dnxKeuED9hJswut
dGrREx52iRVpCAsGxe09fywiOxQR93/+pX7eLrQdgz4OSQWjaVRYPjgvDQ+3NOsn
0As7be95DKwbLk7WwcN2J/R5Dn0KEKzjFUrGZuvuLXDvzS7I/1jirLQtQZtw9iQo
Ex/mPRaOv3DTacWgpQa14OMznXPz2QdpIdCKVxMqHRkkBT+GD8fCHRt81QP6IbkB
tzCtpuXyR0xCP9NcLxcEp2YLFt7u83h9rHbsIO2pZndZibOXeBK0t4ymdwTW4Sj5
V3hTdCgGEyQ+eHD5+uatcq27F0389hftiWSP7FTu0Z2lUFM3Dmpwfw8jeiZKIoDv
+YTOUEjp96xB7PK0aGSA+QhHUkOQe6t+VYmxNTER9Tuqc6xPVuNd4lzRyAcsX+QL
6KbsV4o3uZXFEyKikOYzs20jtk6h9Z4m3PZDDX/HLOPNx2qlWnFPHRAJmCl1UR4K
RmB8iMdvZF0hRk/dvRSnjRivf1z/ZuEnMRcSnmyhcQXj/pEoUb1U2hhCK0ZhYLkR
a+onnx7XoJtCNJzBhb09WBUQ7bcKNW/F9I3Q+d2ETtAIuVVI72APreiIMqiwRFTx
BwAVo+a6EHDl6abYFEVjXLON3g+WCPP46IVIKmN+r1Fof9owqV7Xz9F+mLPJYpDM
U2HlmS8EPvEyzuNgGE+b1KyepQETRrRfciKMHbS3f90BRAZOyMGF0Wxe1Sbf45ys
L9ld5GmITdFP22hkaPX82m0MkdLI5s2WqcNM2TeRsFMwEJFUktXxQpyNiLB5Z3j7
laCu2lm31SUrNFl6oSQZSfneZKVci1Ay2IB35QhdKgm/KicclMmi1EJfh2sT7ZyF
/+U/x6kuhLFnU6Kd9j1yOorYDKb1OFlc9XbRFNWM/pWLpAlnqbnpLiuE2nE3UeYN
7pMUkTVbl8Nrglz7Nq6zlBs/VgLVY3OeDi+m9Q1CzSDHOrEQ3lNxr2iRdFv69IRp
QyVAFwTaVcc0Qigzug3HQEaS2ivd1n0tLu9tbRdrFyvwe6rNrP4EP+xcs2WVWI28
Z3SAondTWDyZjo+X5wN7B3ByLqdgKuF2SlhR0rqAyRc2hBQQneDHF0LzUmnb7DIJ
gw+a4WvNmp1BGO81ialE/wzSgJGpPkZg4l5lSxdge5CzSWL46/KpR1kn87b+CbCt
lA4YOP3S8oTPGfIcnfhzD9RPm/uMvcqY22IlAhYvDI0swO7euyLnLlM3NPgAeKKE
kiXRuAp3fOd3+3MgKhztQelELZHeqmTtsxzZ7UkNzwV4ngrQfuQJJIDmbQ/ImGaG
SkcJC2scSY62VGvuv1PheG8/NQOGyhRR2tmShFQmPIHVUSVSSkdX8Q4RsjPScl9D
nu6sUIrIjJaW4NssbmFZ6Vfb1zEq1Ln5HZS+O1CToucoSHB9f5P5l5pTSpNbhnfh
HxVXzIavUJjNsq+ALvO4WI6LgczVHjJnJHZ4qkj3dHsYEdLlHJqpa7fNKyAFIDMX
EUdEqgxYNrVO4dCMkxosqCcNVaIp7eVBrWsJrXciARmE79gMeCwRd+uU7opgioPO
alVwSX8Fb6e+uo5qFsd0bCilEDNmJYDPKGvdCjWBUMhX67naVwVfBVeeFDEPux4Q
gx8x4Lc9zc5nD/Fqy6sCpcMF4STAslPPP3pinqkJHowwtVjRpW9+h/EZZ6GmzEXT
T5euBo2wgCI7HE6nSna22wV/zr+SOTBX8c9/naDmE5gMdvQ1iJiZAv2PvOH5lKoI
QsB9OmiXZSvKmtZ4u3Br2AQA4qB9pLaYMCKLT9ON6dn8iY1BgHQxImDClTycifbG
bTmu4RUpUcjMdL7wRAGrFHVKp+M2GipPoAlCridWvfbXWqT0HKq08I6QYDEdTPq5
MAxXvWn58irl+RMAlls8T5eWLnNWRgepO3c5y5e9W3+IGOklTwgCcGa/H10fi29H
OVBwrmhbMmXNB5oT+yFPJE/MohPZk/lJwDrwj9RwHbswbMQwtfXAQqfDCxI9eKCN
74gQkhi3K86LkQ+GofRt3gyPHpR0t79fvlIO5aNYPadcCC+tsOxReKP4iB2b5gQn
qHsCSQ1Bsa1JIgpm908lPCthDNVvfUv/FoLCnenwfWDKJlJnGN6hDRjtsVjhFB5k
xZKsAn7KSd9jngVvzUShY85nfHWk9SaJGjVZr/fagzezJrCeURNOh8wU96mIR/Y3
B5z9YkUbXqe81J80uXqBbG840/86EvDha+GdawQjT33TB7y7uyPALNW3HeP8NVxp
xo733wbXWaRSV8Nyh8kSL3JwPEMWtb9g43hcu0ihdkLoQZ8ik7/LI1y/SWlQfqnX
drwdJxRLXsh5LfZ4ZTPGr3enFZQIxCawWGWIIuYtja3QPyXuEbdJQ71Q8SoTXrPB
Kc2xues14deAU9EjtSWhQNgxet6KArwgLCAPToGzoQLwGqBajWctpgizrHaMUsXr
UBTj9Hxy+f5U/LHyFEM3i6bCaIzrUM9NQR1cKytW11bBv7s2rrn+k3ac9tXRAJny
yOSzR1SSKmx8hGaCitRS5rKZTSpydwMah8xDWIyBMDPSUobi0yd76159bjW9iZXc
4IFRTefnNQl2uqGbYXNaGkNERroX4RUMaLCgL+rEr/OCsYHPMQa4LkpfmG3QtCGX
jLqTnIbY3190/LIV91Pgvt5M6TJl25V2BW2i7WRnYs6Wmvtcrnx77vreTlbfC+G5
tdlJzAMH9vwYxoEwzhVq/zKFwCabWqHA4qcsVqcS6/+DPFWqo6RGfFi7lmfOchqQ
RYB7lFg0m6J8ly6ca9VpfaCy9tRaePqSGc+K9Enuh94ZkxQeS6swSq/RIOHyERVT
8FZeh3zRP09xa44IYSMBRUYic34K/ozdGzia4hQmWoCPPk5J5c5CSjYunBnVMHvB
3Yp50mEIibAfD6u10EkOHvpqyHCMzL1J1QW7bKABTuqmZZWrL4mmtz8t45KZiBpZ
UzlSuRwvf8Soy2w3fa/DbBmvZU92xPORjzgWap2BA+2Kv2flXok9h7QmgRU7EnE2
wAm7aYkKVJ2KrsFeqMyEfxEoUZke49iVOzJozyoL/H6qs6OW1wSjRSmuwjrY2PuG
rcTH2SoFuTVyfYzEjTbCbVipGZlQ9oKsQRF1vqLYH1+T2i8aCiVmaEbXq0SR+ZxY
GpTf7MM3CKSomSQsOWdsgGDFuP0QDa0B/CO1VVir4wlBrCMdY4dPFtK4FzYiFhIo
S+9Wkvhn5+uR+fmDcCuT0yaecDtYnwv3d/ODCQSJU5mKccdNIsZ7gn7t/3WYXCYy
B2Uik7LU9rc330l6Xh34Y2X4idxrMwnCkXeBwQ0+6ZzpUZJ3XSz1PFiPgXclg2mo
4GLxMng9iDlltaCdDRtTZXUMJgzUG8NPuMll4/CZ8N/Y0Eb4uwNEpMoqQiYTTGhS
3VAUDlpCEo1MjdHYR6N23ZwwOYRls10n+h/MxUIa6Azsk2HCILQvEJwYdkvvKQSa
vRanL0ZeySx/Z9lnTeQMk1Un0oAUSY6cY6UMqaqWXBHEfivLDmzv9XnTnDr9m7ND
c8lTCn3T0QXB9wBr+9IEx4whFL0FdaJLry3s0HLEUXQ672f+wEgW3Cbi8Cp95lPq
6nBHR11jRbmVa2krWefHtGs6Jo4iJOwoV7pgP/FPIAiKA8ZOZIpewVjW0TjgeFYM
aDtNhWFEqLOZQGHx6GQmPPEXobWi8REsFrjgXvYsehMMtrPMUrn2oU3+IW7U3Bzh
1vSaeQq7mWEgM9Goqsxs/XTlNx7UKsoYHnmmnFkL3JXHHRosWN/V/AWCBTUfGFdH
snn9PdGnOcozq0SZFc2lOOXLDLgqw1y/Q4qwSTatZ8OIxi1HFLMKKLKi7KA7Desc
zes5fuYKJa6iNh4ie1FZ8GfAAvSSmzcnxjOanVDkcYgl9jw3hUWZy8ykkzzU0jlo
7FIfTB62Ofb5+YtzBL+z9RwqvaC4iiPMY5/0stS3tBRB/dj7HemcgvhJ18uEXVbI
G5fFP360rCwIZreMp8s1QC1NmOoW8b1zEgGMqG4Iyt3KUFqZLvCn8S55+WnDkpYy
iIVeIXDHIGhLdKkTzkxU6cT28EjH0tKr8JMIiL770dDEZO+lKziJ/cxa6Z+7k83/
Dh2wt3gwL4bHPq0n66CtdEYuR3cZj59RjxKn88/bbJ80JiRva+qzXGr9SofpAw/T
e9N2iiYz1K2/KX/5BU0lZuj/dHswfl7novD/qa/2oeLS8+KWgsd6A18jq5TQqWw/
v4qb7QFVaQweAAkWWd9s2WOpvxpK4N5N4ZwuLeS/NLo/yBRjRdYGUmcEvxHeVH93
Yslsji/tPD9fglNAjTehQ3QRGTEPT03XruIS9LzOn4KujBXC/RGFQLKLTNN3VbdK
ERkxrQipOde+/2Aew0PGhnjmHWeWuAj+9voDwCPsUCZXlvcrWAW9fAomgjwzG9bX
dPAdoASRai5qyrvaB4JVftCtmSjqASDfd9EFN8oCh63Br7mhi2azfcUuCqXkhysd
5UueKU/3DhhKaD0F9GoEkyeVsBYVcPba4wmVEJuzZ3aER3bzUYPKuuWjw8gBSPwl
zJY80RWYaBIU2Fi6/cgorP3pa1wlnWHxgRhhwpVAgXMtH7cLxzOHuju26WBzELjE
Vbx1KrAv1Iip1vKP2uHE3wwlPtRyFE5yEL1PP01wAX/W68ydLDWT/oZ2RZCzMIs/
aMSpy7SrhZwfwEqMNsHZqh7EXH0f4vemE21psfKyg+CY5VGGuhWM8BlkQCzgnaTh
fbUtVugAhXXs1TpGG7e8MwNHptL34w4ItwnmX30bKOckpFNwOGDtbhmMdmqWD2Id
D1bRpcWdvK3N43CaA/BP7X/3FiHISJ0A78CdzVdPa23Yg5XEc2eo+/mGfxHjHYhe
zmE4WFsNBZFckDj3n90ClQmNUiWoS5OS1xKqBehrHzFUZT9YJgA/gj/yAAYR5eDO
sSzqsGZiqDlFgAkXL54XVyhwr8Gapkm7JZWR70vbM33U8XxycqdusTWgLCb8kVV9
8/q6BagPVGcNn0wr/e8r7nbr2zARy4ngT9QsNS/ycl2GLZWXE0oq/zzT/YNR17jE
kHnVpj15GxymUNoz12Sn13hL/DFAQrcjzBVB4esDeuBOxx9B7TplzyVajN6rtXOA
rQmEHOjuh1qR//uKh/lhYEyRQuHWQ++5A32z3+rQmtO+VaKyB3u9EClehm94BkzY
35I6QZY2iHfREjJl7pY5GDW5qB3ElxVtOKjtcyMZLQoq0pUzdtdAvut/EQ8Ze5ll
0HzEPTOgdLlQZ73n2mqzKJU97s/imQrkC1zgB84SSWCT2xfpnWm8lHbsRKyZbJbz
ROL/gbS7YbRS2U9SxORaN2S2aGLseSo1pmgnNhZuhZKAcCSl3QZ0hlWq7DDGdMm2
7B1gbC+gdxqJf12NLN5IOVi7Lntviw80uf+QCGXIekSNGogA8O/CP9//0AYGEDPY
RvFep5M8Hy4dwRCDqFZR1fD4bJcAh9VPjtfr09F7xpN5EQiSgV01Ys8oFntalO0U
evJeZJVMRgJcPUvJ8OFLSCgdnGnfRXu2UW+BKLRekjMlg0kzlCBolWo2AkouS/SA
4/m3b20rGDv/5RqJ5vQ71Llxp7PlMaw6UrdZILb1KzvVfAD9c8Kz2jDMYj/CRkbb
F/HljeCY7A/LkYlVGr4rjDcC6Xf9Bt3qUfTpcLegua+aQ2K3dNcjR11ia/Ja2AaK
qpPaNYXWx7u3/Ca4ggTOSqd+F6TbkHbbqjKdYrfeVL6mS5S8jvR9LUAGQJeQP2XB
9De1LbSK9y9XOlw9CMdNEyuuvXsAMMiIuo16jJiBlbQ3iaPr9Rm7EZ1n5rt0dTE5
9TCxpcDL4dN+aTlFc+uxemzKhln3nNWnaCMuGWjRgT5hYVqvR9PXEO2JSzqwGFUl
cOxTeFxHRpyv0lHrp/gUBLG6aqOdjNzIhnopGWffL5LPW3ZAxjiSWf3Kvr48Qhha
J1l6znxDFnvIw6rXR+15jXA4iPBVpxFUYDbWzoLubfr1NT250sD4AMW2zxZBtOcb
yHP252Cj7qz6O0puMR9fIDtO2KdoZIrApDrT+iwEuHaTNnoYoQ8aUnXY0+QlAxD/
s61jyN5L8hjq4g/JuPOzbsbnXixGNhth2TFmu0PPDqE9AIGeeKRZIOK2MshC9yW6
7kuYZFjzWoNDzgngSH7tBHWx6UOS3U5jgtd7kfF+m1dme4OVwX3rcQLOhtnuk5CD
jJf2ubCJyW2Sff0gzrrgq4mSt7l8brbIE7uV+YTS7BmSki6toqwqQJIMe4ae/JKZ
uaBQtxx5/47VORF1m+3k5OrgbBwtB8RzeF5eCMt5iInNAXPMGSCTQ1i8Fmbo0Ttz
yqOqNsK8OAkWsXQ9Kr1OD1lpYUB3eQ4kQkCdnGZW+DY4cyudc9CaqvmmLXuYsAC4
4UbdQkZy8Gj6PPmJ7RL3vwqJXJ6qCMW3dsV8F9i3ZtslnQuy0BZ5q5MmJzxyrVp5
G+/rXCfrUos80fn2CCsiLqw1cI/DiyaKbm8GoA9n3x1U5eX6poDlVov9UQM+MTJi
vb/x/ia0EgwsWWe6L7NchQoBKCPI5L5ZSYjF2cynzRmcjUNHxPFOHJ4vHEGs7ajl
vULhNYDZWgUDdHRbZ4ZmC+73TWh+daM20bTm9ieZD2K0SHYJ8LfbyPkkJti+QAGC
RjLW0k60+xWeiNUNHc+yZXOfl8AaMBNI3UVR6V/whKTamwAvE8CZFkcuQRrdZHPL
/ZZmrvn4TQ+RvIiK2cLE5RUtj5djXL8kUHxIaCjuEZJoidTsZ0g5nbElX/GeBr5u
i9GP9Yaw1+m7cvlqFsuXiiQMlxIYUzyCbzDbtPA5s4yEKw0t3prczlHvuO/Vfeq6
yaDaU9g2SqbxJ9EBJWinMh4EsGwOsstUCIrhiBKMCTUlvPEnfp0tlmwIP3EVuBAZ
CvQfIpjhad6oV0j6lI9sMNd5extKB0ZmjvkM+yP/HUYcVelSENuwIf+Zsk32y4hJ
KSDtvCZaW9D7TwNLhhJv3hYrrYDbMkfnPod9tLeMYEa84m9vsd83mBZJE19m2FeP
08g+2M3W5emEO5qAwJ5CV4mSgivS6OlnwwhJqirevb13WoTMRoeBwhZi10NE8IYx
xwQaoasFURHz2T0LxS1qhMyAApYVwkK6GQh7tmsf5P/xNK0dcSBsE0rsL4Fr6RqK
43e7pECM9GMrVk7PPxzCsNgRg9wdIttZUxn6YV6UwkPKpxaimv37KcaeTusEaOtq
riNxVr02C6Jz1q6R+XLWx6oGeo2WJyhH9apePp2R7TYaN9yCpl433uBDYSUwUhWU
UPpOtR8+iTwALP146xUxAz3QJJpMN2+ie5VHg1fYpyd18f1Q0GQ81vvLjXCdo3e3
cXODJwZSs5LAjC0epoO42oRXJJawgam+vJtUoLTVGyUpa6oSS8gbDshqGzkT9bo7
AcIPNBaEyzjT0xsvitIXlze9BEWRBrbOAlzBtfrnJ+p/kXTyB9OsZuwLyZ2PbHey
5RvhMPTFjS/3seb35tK04rkzIa/03l96fNP6+rYyCVrNuUR9Wc+fgKH988YNCojH
8pgc5ZhNzdirfaonCVQ41OnFRQ/DDxeDBJKRP6pgiPEDIC4lbHR1/VJHifYkLFPZ
Z4Cd3/QtYa+OIUdEXfEyz3SBdkdtqfM6pNEqi+RoeKRZ/0kKs6VtM+suwY1vIVgN
3D9j+MO1gFCUhPw8wTbF3kOwkR46qR071xayhPVE5f5ouYuNp18pumzLW5+oT0i2
qoTNO1hpZdiHivf+zZZWuk3utMEVPz+/3lH/Vd++/nxdRh6UwxtnCCGRa6Kmb2Ip
7be7Vd9qicHB5bBFfY8KgioONEIl80m9YIj0F8YQFhqQ6KDFdedN79HEvLaaG/Tu
Ux09KX9BuPs2Xu8fyFyfPd2YGckUpGeLaYZS7QVyO9LokHnOrvNEm9pj4+LZbiwm
J6+rLwTNxvuYBazpFIhHROTE2JwPIo/EtVWJc+Ufpl8sMVc1g23HtK0gNYYuIwmK
aMk0sqqY+FM1DoIrsBJz85iLhHiLZdbS3jVdfcjCZP/4SfqkucVfCoZvWcnR94wQ
ksoHIGx4ihQe2VEzuN+8oE/c7I9c2imLs/idDAQWs1pDXR1BJAVSlGiCD3/0LC/s
jxvpZnyPGOhs3FHzOw1+W6WZzuFFqvQBuT4ctKQIVytzDgQvNPCen/SppKnb8JXF
Ds8NnX7ua/j9O6hXkj2jF2PTX/ljqQkwvRmPMPIYOJ2NCpn5yZVxqV+lg8XoOe51
JpiMjmEwYHn6D3q8h780N5GQAeowmSgQg6JjmDfxLJKkNVVsnjxJ2o20w9XzR5+T
33y3duf88KVA1P7FrQu/DIEJQiTV2gTvc56TPDNfRDox5h3Nt0guh279phy7MY3O
rW1YxCsDUISW3O6wNWIAetoX1hBIlCZWMDUGy39EFz+MpWOQHkUiGAh2lpCBj8aL
fj4Gyk0EdUwL+Zfl8x71fvPRZDv9+EePmMzcrp0mRg4DsOmbPYyaqD3924M/t2GW
j0ZE3R6PxHUg9xXW/NWeF+qhjKrMP81i+9kUua79oms7kvCkS5OQW5f/YD7222GD
XSXbKbeI5rB+PJMxtsuIRRTFVweUFdNhqfvBRBwNGdv3dXEKqSxHtKLVce2NAF84
M3uBTCRha0FIfZeDyUHgNUcfdrfujXKMc3nSy9ZKB1XDOPbC2aJ9I55pHmoMbJaw
JxSGPXSZHfalmVJNCgVY+/XSBVrLFvcu6/roAmwCjF1GRHe+iHuR22BDiuhlTP1e
CD6HL8Il2QYyyfi7iMwV5O8CueYbu9QREVviekk55iSuWloVevHPzCPI4hGmN7zD
85as5pR43VscRYnwT7bcPWduydlnaNEd3A0FbsSEZUAo8vDVQDt/5fS3ZyqOoYlt
8/0vt8FMamv3PXjd/VyWVSisThaJgMzh+Wd6udKHHUgW9GIj6ZkxCC/ws9amLuG6
5oi9eA45J2kzVOZIcjZ8mNUDDTwbDODuDtYXnyEwGEJK2aXbB1vx8h5ZlsUmXHG2
EcdwT5i2DcTna8HAiFd85X4HXQ1vSNjvb8NYe8KjEmFCKjGMH5CJsjBFmVILhezb
AJt9amou/aB9azOHCrK5TmmpCJfY+ZtzdLzMg6wif7tH7bigoZFNSD9lIoS+37Iu
40qa/cU13zSvndrcDw/IfORdCK3XEn9RFeeEnWEo4QzpeQIaaGNTDZ1PIsyTNByz
MFbCmJYHTV/I7qKTKYyHHQCsG9ZUUJ3HyuwKMxFL4O58LFLEF5uMqqVsa7WQbIkT
YDG9uNrTLVsjKuZFG9mIGbbsepAvRIcARwIOD2Un0myP6tiz+i0aAPP8vwb4D1N/
TYA7KjnYld/7+QmxvzBpKY7GlwpDcBLGh5WaM/rpiAkFJmdGISC0uKAT3lcdieEQ
oq1Fv7+IIloHfQ5IFBLrAZ5orMnNFzieeddyHcGCo2kAxzpJ6SyHu6zB43KvAZkO
yK8aKCpMDb/9ebE4/E4ms5bK3evWSNrTHh93QKe4vBXyHijWNTaXBeMv0ed9SdKK
9vkpMXpDaedPqhbaagRS7pvodTSagg+v+DfyBwv7xkZcGaCu3SVgCByKrCE8gh5Q
0N9aItXGzRHqf/PQdk+LiPEStbu84yz6/BmYOTcd/p4lYeSLNpd30j60bKRozWGz
aG+5/o251DZEFwClFRjWKU6OPhmEqmsqP186AEvrMoxILS+NHMQXnIMiaThlf8o5
zPAs0Z8xtjG9UMKvKkj5smS28vCdQNFmmkwFptkC/DqlI71LN9cSKvas3yuc1yms
B2ss29UpwckklquqNPH4Ci6Y7chcB9uW8bqNzgNNrXvDzbJCTzF1l/+u/oTOJmBp
GeYVahIx/vohp40L56ZPoQ1YogorxM/Ftn+DGRPdJbnTM0goTypvMzG0NHDb8Pbp
16DbspcvCV6alyyex7+jCoFLIqJIdFxXMFdYeqPXboyx7fN291QB3OEmpmqh7pvD
GD6VREJqVjKwTVDR1BK6xO/jIISIb/AL9aILI7fZugo1xqxdwkNjLZUGNBXSdjFl
9XxgQRxEjG1nXJDg8+o29Av5DifVb2DkWCfOf0KdGAPDJChdsOobMejo0+XSKjNf
Xw1+PwK2PkdrQXV5OsJBwoDoGNrkLb1zK5kjFrzG8ZcEsSwBq14xnJf43pcaF8S1
6F1cOryyzCm491P7qUgHluYalTU5LWVv4qVMsmtP4Y45yrSDJyvBXJZ4esF8197e
VhcdeRFJDKhee2/8K+a+ENlOlX0eIUSs+nro7FBt5m3Fq6lEKpQxRwNLoYk8EwFR
kwlLQ2Pn3WWuqiPZ1t+ytFLuNKEwwT2AaCfCJ4nMFeq2Yy1fAZnXhXYu9VCKxFPZ
g8uuvu3njQUc14ADH8KliETBloNk3e2cmmwKh/95LmXjhJbC33CebukpjiL4YdXp
6fNONFMdJPYbT30+eVJ0igZ17SefmUxBX/iant94vbRUeSSwF/C8XIbsoGCFY18l
LD9aWdus+gGSU0nJUtO2l3j/+ZW0Fk1NuLR7YXv8fwL+kcWK6nHJqBpHIxTzyJz8
E8oMBpnF555OH6wku2V9UMoiNH1uaPjU0ujyZzIA/TFFJY/mNnw0y5ITPNLUG8o6
1UIAObISfZcHNccgIbw8kMFaomuiVzlkiZdVUVb5+N9lz/aNLr22Yex1N1u6spho
uzLh1wyvjvykdZVi/0aaZr4RU7/nOjyaIrcOdcqg3nRolsokKOWAlAMP8JED5LyJ
YOSHXFSLPuNvHK7OT4D/9/g4Zl6inXFsczwJ2OQTamTTRZIz+HoKS9Q2rRlTe9yd
ins/SU2ggnkEWi8L/kNjlMH6MxRkg7t56SbqB/VhrqMM6jn7+bJhS89jaV5iHIUe
iE/W0fqC6qcLdIeWiwKnNkpVXJc6YBuroHxGwSAqc3LmGHz+bKXMrBBpkXjAhk1h
UMwZ6mlZ+XKaTj/E+eqnDVgcnGQTdjyMZxqWl3Q2izMcsGKXNYnLQ2E5RELUUU89
rzmFt7Ea9qQyL2ha4rTBn4ytSqsdZ2Mkf5yJehTygEK/bfujmLKQ/sEAX/OGLzxU
x517FzRwp3GPzHJGheAVNHnNnq/vDoWr28pbQcz+zxO+UskjJ7MwBlxkHp76kaho
Dw4LH3sd9zbh7uJIdQlhnksv3hglzhj6ozyw46u09hPhHLdx0csYUWmnxNIdksWV
K0fdGn7UxijrKjhVfsQ8BoS6tnFKv20cMFp9QscPSqU0d/AsxUJlCkhISGMo5eFS
YC2aZRWC+/vvUjFDnmwnVvdggqrl/YauYihMIgCAL2PN2gTZyNrUUB9NeU/zyTIY
5dpWnr89VZVD3K1klWH+65KvcLgHOhvfMQX/9OPEtFfgPHg9YUcDnHDKHuGHXBFu
IcBHuAfxjzzFKP10O8220EYgScXsGWGk8oaQMuxjxs/ezQeCZh7N7eu1CjAiUGiK
URbSUifzLOeFjer+ek7RwCgf+CDwKzs8KOFk5KKLkmBQwzYM16grBFRiRvED2y0T
45bAtH0Hf/yxXq8nhTKX0GzBM5x3aMovcjZPIHnKu6yG1JfUwrIoAh5gzc1m6Msa
opOr0o2a5z4EHFwA0O79LClUMh4JB7g9EsXoRHJcebMXqgtoPHBND9IiJfmllsrH
jFno0mE+qqNr8By72YS1OhSq0XPVCMXwDi5QqTCVn1c+ZH9lXU1rdRWq1NocSWp7
+bgiKFWHIx4rFt8+71WydclLL3V9F/hUlZ0uZABj8CeCTIdLQLLKT+uMZNMybBtl
Fv4sd+KqSKtaZb1UJhHmYXGPCcRXkqrjAmY+xSYcreMN6R+X1AhZmg4xwvATCIGj
L7Q32gqY06EbgoHZkWbBOh2aUqth8xjb1THEntRFGVBsiDucR3AQq3CqadVCmwYT
o0lQaT3cUo/f5yfN3KZ0fvQrjh6ZNIOE3x0YobdqlBhijgaYeZGDIk9Ebo9Xn8Gv
dEwms3JUzSctyZcWYAYy2ixkexUIpcxdefyAL9l1Ipi5doetPEqFjVaRO5PUWKVf
sCrhFKLYr4N+TyzYjM5Q24XaF7UZAuwdR8i7qV+wdiYsHYIh/ImP27M6QuD/NQyr
mWSyvPtnxUD6DnPgDK8ViarogQkbFKcGBMSNIwR9fJrqPLoOMbum+Z3jVOEzDN8o
jNDHcg3oKCw8k2GDbut9UO5ZVGuDAqEAFkYpeknccDo/E0/x5ER0hxQICBWWmC+Y
VdqnT6F6e4UgU2Pk0wBGjOy/vr6E2e58g2F2rttvc2ETh4lvEq7V/fCuWWTvUsV3
pJBtB7WKSwRn19T0VjNnTpHDNBEfIvCkb30vlb5+Sfot7wR6FevMjL54fuu2Zxr3
a2PuIGeUZVVSiEYEN/IbacHzLb/hOVB/hP0SC3E9m+lvoc2mP+hrt+c9P3H+hDx0
YWAF2WgtS22Wwk2TIgKOQCTAn+Lgh41D1Km4VikOA016AL2We1qO8tFmVZHWl6SH
P8zmTdE7f0WnS6PuVJRjCyVXXH+XmOciJhjeK9/2uoYTg3yF/+3R88cLvu8B7kqw
Qp9CDw5g1f3/QviSouyJLuhsLl1fzvE2fuaAQtkERo/kn3lmylCWbIS/ik7C7YIp
W8ooM7hnahaVohXtUWxHpOffUintWCA9iukQT7S8FIe8uFRfum8BGWE1c5XnGipd
MjdM9Wx1DkivxKgixSyYOw74IXQFf3i+z7ny7frZJuTzivVwvOhjV6er/NKZBv0U
lTgBjkuRhoDHwcmV3ZvYfGY/gAfBme1XxHZD39543yFSTM8uCqe9M0oiICJvc5sS
CCbgSrYJqo2rOHJaZMmWNMzm8geieHlnzusqkU9UpAUpVhcXxPNyXQJGD4VUyFrI
spOMHnYOUt+Cc6nUndqWnJd3AT11BgpBgXilHR1RaMMwKNZQ4mp3Jcx/YtNpvMGO
wqRjSgE0+hplpnYCm8SfPwVrvsfSoUFfajvHZfcziB7EKLnYiZNdzcqPGWIVaKhl
RHzMeyvfjhYYsKTnJqCCGZ2rTTLsGLPSkwYCv35TTP53HuN65DncsDtT1dZEKzRs
HA2OJgDdJJRGDPRDUx9Dp6y5hxdyt/sASvKqf/o7yJJH/D0TTiuKeeYlFed99/Vv
e8qgiZSdakx/4U0TeVluLpeAVEYSyLx2KZAxTMrTrJJey2uBbcNdOvf6h8Ax+2QZ
+IFgq3N+ClvfVxPZAkeUkTmieO1FrrQqf2oET2VCoCUoR3fJfNUaN1g8MthLrzJd
jDRiUTki0E8oxjyR54ZsO5r7jyZqswf5gVC1REBY1ztSmZjdYUacJBy8uC0uHkEN
qxuv124Oq33dS7DQjF9bWR/+UqfZ+cIjAIcK/80xl9//0qOaQt7BwPvxU1BTGezE
MwYxbpDmysCTzA5P0cqsM9EbTtjrhuRgKNLgsNj/YBST1evL2/XhynIAyBYYE9/D
4aHunCXWcy140KiX2VwsFr1OlbZKzj8Ie3S6D/J8Ios0yTGFze83VAzePiW8w4vD
XKhzun1BcZLlHXIonmmR5AWW5ORIORkSvb135is9bu4n2gC3TJZa8T4lTGIqSr/6
HTNlU96qdfTXxC3AtZv8Ca4aNbJFj11asUieOO1wJlfZfBd4hihZRucTRACIw97C
gfwuKFnifLTvI96wQ0xpqtbDRFiszNnhbVjrIzzwwO7hr4pZklBFeKUL8EsnSv94
WUxgeD4QRbm/c17mN9ZDCggG5T8xxyq//CukjsGv5qAygEomhbXUaHkG9+zak4zz
moaRtArgnSpt7dQkfr6WxVJutqQ26RDk/h1LFokMj6jz2i21RU+XbWWgEYyPCdr7
Zf21Ohoe82x6bcJONOVkZrKnU0GQ33nj5VoJanT+NOQFZzm0ixOypWZw4ENUDswo
8l3KUCSQ4iPQ3BQXTgtAcp6PmtZ730rcMijbDv6JUtIqQ9Sa2IK0Qd9Fw+PDtUGE
BqoVDzC6J5+0Cmo62/rpXCNi2AYXKiiOIyQzAwRX4xI+/3mpkWmGe6Y3NJKwLwHk
i2TWZPRAOp+/dBp6HHx2xVqkavDnXwxUmPr+3mmG7gswac+9aLH+bOheHrSlF4Em
6cHf5+8utrEmCYoXfe708Vv6mpgbE0qsUKgzSilXWakilBV2J9PosyDqKfxz17xi
ZpomzjffIjFHfLn5tQW+hI29S0qRcu6Qa+aqwttJaFwBSxm2Rr9PwE2Eq+j3jrQb
z99SvyETL9YwE/+x27csYq0F42Bdbn2D7OhMlaLXofPrMAgeZ8yTWd/ziTrk4JY3
MvZmZb/hwdyvDpm+EnT2sFJUPk/1KOPA+TPeUwHeKklPVRd8q2ROs8AiLalpDLZQ
e0QRDwq45YKsNKG4TUPl1eVbp21NioLIVLQ7cKd38/S/EGUdq6y2A7ew5aJEgCQI
v6ixYnO2Jd0x21zAfKpDFVXXaooEQ8bQWbcpqnybMd3UaHgHmcPDJ9N0QzRpfa1e
f6C3g4Q7Xg/r1yYbhb8ixd+sTZyNwrMDWkhL/UwAaQyFw9nFh6zgJQ+ehZUe/d7M
aovOnrFTz7Se1L+IM3X3g51dKpxE9a+Zniu+VKll/UG8IINGEEKYnpQ66k1wKRvq
gOCC25qDWQVTmnf8eAxOqa06U80mc/2dM8qqezINfthi7Q8Ll5rDoQq/u6EX03X9
s8YpBhyo/N41fB1hS9loxCCH8VcLuKLmsqHRDJJQsBIC2GlnqYXdV0SlPNsLFqpn
Ukshcr4jt48MrH7GovmDsy+PpxCWXZ8HVl1Qjh4wsyzoVelYe+Dvonf+ivygmCjw
sx9IIYl7lmNqXDv++klsFXSVngXezPZQseNNC3IYcWajD+wviytmzfPPG1x3mJTJ
PEBs99oSNtCAmnibunmLU9+IOSPtfoNrdSM3YEts2uA/g5z2/Ndndsk+/+oXedTm
yR7+meqvM7EDgDn55AfgLFbJJoAclUNLd9vUGiEtPl6pQSRVyutM4RGF9RYbO8Ar
wK8E8yYl8Q0uZRTC45UBUM9auFqnoFnL80FCoerca44n+uXoizEhbIDEVM2nbwn6
fGaanJ9qheSP+QFdmuHzlykEaaeoS72fbc+uu0S2/x0ch36ynwXaIV0J7EBLGyC4
MmUbwG3VRUDV3HyP5RVbkJlMGS2i2YLnw5WXiI1Kli3XLbW3gzyV+KaJM2MpT7ej
LieNbKLoQCRfh708hsEdpKaTL3gwDA9mZP0BJaF72R9epG4Fz+6wjrgVq3lhvjve
+70aKs28GYDURhLRIMHY5ufwhtNVzZJyY8XvmYqHaS/WLVhUaWxjhPsqXDJVRZ+U
0A7RlojgT4GFLwfWvUvbc2Ajf/TxqC85e8XERXWgKLxjBVGnWdzls1ia8P0Gj5Os
qyU90vK0SozXVbthxEy32LFn/szoc93csQpwLDyhEJHY9OoaiumFs/uCOHmRG4IE
nazmtgWxKUfnbiQs2SCyK8kYrPGT5xaqyOUyWEksn6L+hbfjlbudQv39fzAprh0x
aGJYzjOGkfm3mSrjNBdXhqm1TEjTIXbPq17KsgiMKcz5NLABGw4934GhQv0rxn+c
Um3lL0FdUsDqNnb9BOqOVXI1gVUeh8XlEAC/GF4Zzct5L7UtXusUkjN69hLuG32h
IOCiLgRcxS9X1Flx5XbtVGjTggQ7ZEJZFsdGlSmHnoshocMzOJO6M/d06gHLbejo
w+RyrytHYSLz7AT0Xx+NdMnKggkFrtwbO+024wU2KMKeUHIZwQZDorzdnpM9GaRZ
p8vclXtcwOhpUQ9juuSqR8ROhJbKk71GsQhLI5QWpb3qUREjYKNZn4jqQuR2G9w2
IHZRdYNVwSozSNVH8fRTfXOlXsrvF96+fV7mXnucCrA8njl6urllDKFk6z9GYbpG
p0G8BUXLRCO7Gb9QRgJlipHVOPVttvoKefZJxIFjv4c/3BbGWEJb5xh7sP8T3W7h
hRYNjJEEc8MRukL8muT4Lch9jPA6Z0yVxIBUAwrKQe7Ls9mpAw6g4KPzu5rI4VA7
Y9uyt+DE0Ag0OBy0Hr9upV3tQNh2PCvCkk33ZWknky7NcLZd5nEu22pmug2yRuSQ
wtpJZzE7pjfI9O7W8+v4p0Q4HkbYwm/LXdKIzOVfrL0feqarYpKgluMOFQDjrvig
wQQ79y5E6+XWvK/exAfUea4F3HNLJLYMZ6x0ZP6NNAlGRWT0t9iBoFkFFavUvAjD
/hTrxyEyJWeDTxd3DYNzl5piL5CP5EEZVSlKXhu7BqXMe6ozgwLj46ZUw1mOpXTd
y1O83mwyuf1TmlAERsXFLTx3hUrfIeS/sdrGB4Fk8iEhJddDb1UfENkuWvTPHoEK
6FxaSMuU67S1ntI9fjI2ZnKcY5X+I5ctPSJPZcVEROgWZK1AczLTsBt3VZ4H2knK
g8BRiFHyUve7mWKhj4oyfNRJZ1DT4lTrl4Fs3pWdrdig48oo5UfUCrVBQdEqxihB
mkYvZGmFaHWjTaVuygrlcwfBSQ8ZAOjP5WdanU3oGblyxWY/dRK6hlLw/bP3dBWV
v397yzxL2e8fhOXj67C8xJKWtB/LW57zHhOHdrCCGRdqFInrc4e8Kttz5qO4OWfM
KSi8RyFiUcFz/bsALHLp5+bUd8MWYrKSpKHrLra2PCAtnd3+aHy6aEv97UR8Jpp6
WSktrvxusxD6PQ2Gh1ZfZaOYrZa6x8ISlSAvOvAuEPqc7dql0ZibvukBwmF5VrWg
jWq3TleiWqjhcK4X5+kja/KQKKzI9DytHvZtsPW10ViQecX9MD0HqJe2jl1zZLy8
iafWAdvN6/DYFzTc6HIp7Ocsj9lDeTJ2K8PnLHNFAefdF1HwqPRzSQz6F2KKIs22
FZprdEyI4BYVxpTzHOcyaUx1FJthmTYp59KM890wbdo23Rm0urHhe4fdJ9F6sU4Q
y0K1YE8ym34OSaSZ8eA1CuVDK9CctRrV7epW/d3/ivSdBD8cPNaoPhIn2X9+IG48
ceKXnyrmXLV5YR2la3F7m5c/05Q66zwsv//PsQc46MhMeW72JWKLIF0yiRg/4gkN
X6Pw2l5ldEEB3MKt5zu3MFMFSADNEHcoWJJVDgBd5sABNM70pPWznXzodQ2A7CAL
OvETI74OcvsTPka3nLzE70TS4ypPKj3kzug1iL2Mg/xRf6mnEyP7t2HlknzEAS9K
6+VRkjr/DZlXVHXN2vkvDQTx1BpQFJ+I+KDN4pDRgRLxwpgHmmiq7cOeT5Q6wvtC
lLXQlPfTAc+wuhiRZEK8JOsWU72030Ek3NjZpiylFcVUAeFuv4eoXw8U7E/3MspA
rva3bSdR+WkJ/xgLB39pDWdq4eMyxUsTYjk/60I9ZZwbPrJzWyxOUsaOuuQ9ABOn
iooTM59c8UxCKGPfZTaAwr+Hw1wdjscEhRp5jgO62JdWZx6y0thzBz06XzixNLqx
niokEV0mn9v2ly/9emBGjS/vfLyE3tq6SoL7J5Hp/LWOZQRv6K/9hbKsO4eAecgB
99HusKOqqkWzsGFoZZLmFqUHkj6QtsRSxl0mAqeMhO7R6n4xDAVzeF5EKY5szU+K
7SgV1X7Tj3j8FZYG2Mbr+GRFp0FXU1uwryBa+rn2Ap9fH35f5dwoKiPD8iAX3i11
/pSQYvNWhOLUy22URb+bWKOBNf3YFIqI8+AkO+hq3EkpJtfQBhneKJ0Pff/0HG57
bckaHc5FQmqCgPkGeCKBtIyHp/88YKmjlnVrYVUEqktalK0xRtVd/jxyk4NUMa6+
lMYaVVI1Zm+RizZV2WW+3eh+5rplkEk2Lk5eH04GYca9S2rHxYo2x9IHgeLEVjD/
u8IAF5o7OunpCymv9EX8HswWFbf398Q+evWT+ERg6ZTlExwxDrYyvbpZleUvZ9ae
2et9FdYHS/Q+DpiL3VLUxPJicu7sjvHjEDpW2tRpwmB4+gg5AQ/7Mdp1gVTOI2Ff
KGpK+rd6EDIeUvfsbR1fkqNW2H7KeO6STQcs+XV1aNyHE6uoCyIRN4O3hTQQOIHN
Ws0Ns8Udox2UtZvdysUwOA08cbvV1+z+YQKrTY7W0L/3WeffPx09gjxRRIr1/+GJ
ZMBt/95jduySIJjVygpBWyxihkPQGpsppJ1L952McjYoDiBreYl1UvaW6A1DVSVu
3+azjf2k9i+cS2O5qkPh8heQIZd9+4cO1P/+pkHbrPRtFcAozpMWoeDlvu0vnhK4
dTVP9ZLFtqfPz7JEKLbTgirg2MWguk+NqHpnU5X+0Zvy+DIEyb0CWfoBULKZsJfg
OqHSAoVyUq977HzA9AM4sUDOvnX7MFY8CYDuTxMLHFgJ+0ncvkxXBVqpggJY323K
EaTzJRJsG51hK2lLZ3/QKGnOQ/JL0cBCLalt1PC7pzbicFlwXJhMuxdlJ7pX6yVt
M6UQiQN7raqeiLTZ+rVzvhy0v+S9StearGY2yvLKAvemrhnYRtYepk39fsG1oHGp
Jwa41xDWDNmNtdLyCrvZhmLGXH3RaLlTkeyL/GDS2/kL+Jb2lS7WwQ4qvJ3oc/+w
tic2C84poFKaMOdLYxDxixmjK7GY7UBvuQ5mn6RXbqllzMVE4xmpbx6XS7hbnUgH
LlGWN68/0U0x5+BiaHIaU5DP6vV6JYfWkGJoN5O8005h8Xc726nx6vSsKHb6IjYx
vFNasky1RwOD6kQZYVeclt9x7pNavEG5lZ+Ry3398Hhq5bMHYd0Bw1kqhTMJWyUW
XgYGfLdaDgl7F1kS2az/uUQ3KITZYKT58bBpvp7fgLGAZMh78HPTW/QViWKR+O6X
g3RpUwvsMudu5N89rlGXuU8QFysmnQCvIPc4UUUbJIuMt3FwFDcSYq2z+vRJIR/0
XMN4JMR1IZShvGEI/cyNHqi7Y7vBayUCMYV+ypkHWjDS0yTCRuibqW3xtq8hWJqg
K7X0rzMERrrNKZeHFlZuZr9j+eoUg/AoihZLzNfXicHtpjp6tUMn9o2hjHmFdyTX
kXkUqAjoXvyAElUXIim004h0DGOiTWsfWDAHH8aL6ZYWwxx/bKP5IuuP5rHqsLKP
rCGdynq+hpMWzLnvft/cPJB30v7AG4KRgxFK9M7074N3FeNBDBfbSU3piT5K+M0x
AvbKYXY5/aNUN5OgQ3cH9TM/xyiNrS1fPFnDi7Jdosftjd4777IpRXCWvsT0NJ/m
lZxncuGouOkSzLhfv2yxaG/8kG/QUINtpDC5m87xiUJwl/GiP8HlUKDNNRbNYwmW
j4PF3EEyidEPydXn9PykxafKgCeI5dmVxLtYjhl74XhgSHSZbEB81W4FGD5HDXZI
Fwq4mUHZHxEXugWmUqDOPI/yxnsgFEZJakhuITnLtxYQsj70bAVOXzXAyeKqe3eK
geu0IvbN3oEjkcICIeI1FlqbGw/MOzpUniCE7+NgZjby5D2qP4s8KaFKZolNAhII
5i4Oj/rx9A7Y4vA176ZHfO1TlGRFf9WnwahvXaXns9wEwtV6psyAdlGk7u543PaM
QDNBqtw/E9SLaEfHvTd9cCgPpR/rUfcFyMvPT0cTLfMZAAHJXxKVny9qEzcP47i8
9kXXNczqy0SvDcOMh071T356m4usazI9aOixWaXF/WZk81aWDaIy5CmkEIXgnNVN
J5zFTOGU/SepbvI7zJHYDN0hrFPSwVZ0JSRlbQv6uVIAVfjOuwokvm+oXaA/Q0Hp
vMzTnBL68iu+O5a2m660fY/DZqhk6prFMDdZbIYFWovqYoJtxD35erJNwGH+s9M7
FolD9ffK3zqn5ALHxIcr4XwI92LK6etVS7BtHXQ7MaYAqkxLB0dVeygB561BXaz8
A3Mru1/VXzgbqjyNgX3jlOm1iNw8GLpFZunYl2ggyntpqxAOqIKZ5UUpG3WiF8Tp
IxyWgCoNqzkwG80pHzIyLcmJlLp2ZQPjnfA1c5rDrOI3pglJzAhNbWCSaDs1QoJo
xfqap8glxkc4mJl/Q8pTnkPny0aVQVC8kLZ8SF9KmsLoucPw3ALvaD/La687xxyG
kr7Gq+ic9OcAf8OxLCjQRJt0PNN7hheDCmUa3YsCLDDlqTvu2K0Vk7FBCQ4I2NE4
4LegxHgLZuV7rgpPaaSih890fFtKcNQvBEnNHkfSgYQn0ZHnB35EwfPqWmq9S31k
Ju6Nx9HUC+rhIY56D19nSoOzB5By1zPcHD6JgZ3b1Uk0WpgqnILCL7XyksVpVz5r
CLLW665+59TC3Z1BuzuX4R+pbm49OkcKpaimwsfFRzDfkUTPLOEHIu4rTRz8w1PN
g/Fwk6xj0Tn0bPT11e9YiktWqv9tMOCPYUVpfM9BP9cre9oE8fyFy3REk7tZJVQe
0znUS/9UVFDfBlpBYc2RO0F/XeFDUsG6cXX1s37kW/EBpSG4muraDuGIV3aiaBZE
ZCJlHl0EXW9pY33tU0hrkA80Yr5OeHJ3BJaM8N97oF0TmGDEjiCadEtBhV9APcUU
NGkDE8oz99qo8M1jnGytyVEYMbxOdso4xP13zCmhKP3V/3vprflFrX4OuBp9cbeu
9Dx9IFUZvR1tMDTOGofynMIkFSjKOwbUJCrZUnLgmSZoTyK3zT75YCrWlFPidF1l
VBNW1vHI8HovnmZhxUiZ8OLopF3qSRSqSAspDVwAZlhbNntmFpnDhqBr4+9CEGVw
u2o3MtEB7exAyS7maUKbuOD0OAXyOavEqMkaeAZ/kcc548xkBs6YlFtWThXzLxXO
erwph5S9fzy8Ax8Jv6dF5mRbY6MaK4UgUgnnQOY7WBunWNGQ/XPYT8S+2qPNiLzo
XYXf9VQChOhjlHsYa84mU7OKKXGA7I4qhj20L8zx5lIYD1Tuauvj1RVRi66sNT7Y
5iO3nkfPLlvh0Jfn+EqhwaAg3rJ4ln8fw3YvFCQbSS+iyqRpxN5c1+pcLfxXfUDR
6nLHmUijXm8bUMHNWzPLFM5KQC7PXRgXtRduoUgRx+qlJ/h+t5FsmSCGNlTaDnvj
jzb8u3wYcXpykLg4SHqwKqGDfKLuOmg+rmyNs3VqeKH+HCWm1d7tQNXzGNsW0uMg
sGg/oq/ydAts/mwkBZ+KZudrdM/7Pco2He2vxYnVvalpVQqvZK2EbYRX/numj6dJ
mFQRzu97zz/i6WEfOOqmIKTTF0qZ7Fc7GD8P2u26os9mjPnzlqlu7xv4RaRF575D
mjbkf6KB7zRlUXj+moK5KH8gGW4Z12Z8QwT3X5X7Ts1g8MaY35wD0TVfEDun7JYV
Fs3sDsQJL5jDJYRJQOZ/mL1wogzeSmkRapYjG5udzvtqUzfQBFeURer9LyZsXNyI
8RyD8uR4sw6XJxT8lEDcu+W0VFZOpGKWKfjSG8swlvCtf+i9RsyrhC0dOLOzmr6l
MlO5LveTNzKyD7TTOJRgEQ8gLA4xWilsOvUNumUpscSPmddjpwTRm0HZp87W3ZYX
7ocZPQgScjiijblRvfqmJWWtAWm/bFWHU8U1GzE39b3DP45LZRM8P7qb+2y91e9g
kuerHFxu6ch9hdlrpfmka5LgKhzJVV8DRbujwJcgCWWpl4CB6xs1l+5qCnpkHrtx
ri9WIoMGdVBdc8Fr8mLMw+2uU4Oj+SZGrlWCbPQxWm+1hvxwIUxh1h2a/GurW8q5
n2oswTzyz2z+vkyZHA9XQFkgV/6f5h/AVslhisvYCTIELS3/TH2T5zCaUdGxp98e
90gjRlYUft9r7vyL7wl1REc7leRBfaVWpPt1I3qSDcPd16rD72zWOOKHBJV+Pstb
PfB+6gJl2tcEhRFi8bqiSbvYMbTHizzQ+tKNKlsSYJYIvdLkNF7ZqqrNlzaTonEC
1tbfItwZv0zjiPLSlOn9bRcNYoBLpkuWro/6v7NWH05mXJPXbeYvfF/l2JAkMCtY
2YnCVQYavFxGFtPYK/Rpug4ucX7E/gDEOEjFCPpfbkB4XLKK5inhauuOWedOuism
qtqr42No5OC6frJ5v7WLCHZ3ANJcQbKhuLOamqS/oEGJxpUW8N7UG1Aetsgf4Dah
XSs8SvqYS1dUwdWP/4P3ggkZXDlPkpDXRjb2EefnbdWMRos7WO6QpnxsHvJF9x2O
Z4RnBxtz3EA1vedrAhgymJSRiW010rDKMOgUCHYl8xBuUCOo1t54A9XcENv75yk3
VZSug0UAb2cAf2Y7u5g2lvi9t2pDqseI/FjdvGED9eP3Sv8vo6SZidG+iYtHV2Ll
MvILsVeWuNbmSUGKMm6TIHo8R0HJEHJ1qQ9ksUOfxO1srTotjZJErZw7AwWIfeVN
oM8jZ2OLMZ1orOj7szsbsfJZMeVxlhOgOTz57okLvg+1VPp79lc4HdTvjK0tvEod
fy4JvlN5Z6E4cb/W6rE/Qlp1TCm8ocKp+5BClKQoYKiGXwx73DntN+xwu87AI1tt
GuS2AfKaBCpkyYYTMXC53dPv/Ut2kRaX2WHbgZO0zquQ1hLCIvylHbucTVpb+1H7
5wB6cXxWfa8BkkTFaazUgxO3oduy+/olXjM4KdDm8vmjM6u75s/NMt7P6gT0800g
IpIDy5PdveJ91dmYaYUsNkcbSct+7vStbc1rtqVPB5vKfxK2UJgDst0zMk4UiInK
AyUunbB1zE4toza/UC+eSRxAYShUjRj90ST7tbuodx9z0GgkPx7sBY2R5bf4ZrKA
sTnWgt7xN4jgDrAD5QoXh3G2fCNkFgRtPvo7G9wn3AeFhUBoJyBpnDTrINbyBdyT
btnJBGYjuNkSvyvfyXAvRupe9odLNxNrTyybe+RgHfwqtUZxqjoQ6mS7PXVuIdJv
A1L8RUr6HvFtOjrdebib78oZquHban1rhFjkno7TkFvtU/bT1KWupv0aBvSl55HK
sUg4sKn8b6jZWGQxn7apCODO0mzuwVjAcMaIk051uhkYWn/mvXu4Oqv/YagL6pmk
6u6KOX8WjqMLWVPc8H5Yc82qX8CbOleozT1Fum3IBssjSiIrJP0LE3pZzCJEGO2w
4man2YDpA6GmwxcPHxqr/l35SjW7pygX0FchNLKBf4Sum5E2inLVGIIkirFjpkKX
XokXO/fe4FuOdKsUfl9ZxTLemr7ZY8IDTFsUM9UoQ2RjcMGQ6RIOa4amUdeA8mhz
Rpz9qghgPLo/NeYaXp07XaorOEMOHM5aDkPdIXuaB1b6th9YecaLy4qgbRqWkkD1
W6e9sqn49RrAlyLjwhubSisHK5ITROWIzyNn5BUNn6qrCHBXO2cbxA7yNQv4dH73
20dzdMUNupWrFl4GaMUnqJCitWLwJSLjvfqDHhjDBZH7uo1c8qWpTHssZCy+p0AC
Ek0SQDVMY4atwdlMNBa5W9cMx8WTPqiHkzMLIAb11FW10shiQSc85XI3UUOwFnbX
ZmnYQetFR9OgGbChirTzo/slKeUZQ8+uuQJo17U0WGkHhEDqG7qsd0PuV+6oqDi5
bMRqhlRgRtv45uX8bR1jPWo0zYDQ73g7f38vbfIN5BJtz1DFCiJRy+i0epfrzjtl
HN5QQ4JTfK4lQZVK/7K+0Z0Z4W7f4c+Rf6IbCcbYhYPEh2OQO/Bv6KIM3M2TCZh4
GbmZWF8kr0WlAsDoOVNPO89J1+xM4V0mJW65QWqikcbhbnSSZTpaA6BP6kMK4/BS
RkeZXarI1O81BYIPXzgdoDu+Q4iFTgFJ7aeywCFUALt1XZjywT3zNrtN5uXlVTHY
alIWNI1t1iTWLOslvGkzG77Fc+s6oBMjsJW4MfyRusmiTsvn0QeeHgG5UiUlrO1V
Dvj8gvCf7cYlWbGYGFc4NxLe1QS1VoWG1qI+AaFtJMq5mTELqZj2VlG7oLEsSI/0
Lp1sFeZHsq1ojOZOYa47fGCfD97t5KO0Dwv9Hs+xjkqgeXmhnk2COSybm2fak4i6
oK5WGGzIzn/HfA6CJDWUvtMXYBR2PcSUY6Z8mpg0H0g8Po0oku4WO9OtI/ZZjttG
GphW8YlT95e5vy2nravBw2nrblWQu0J3+9OmeIeY7+rbCJc/DVRM2kR5bD83MWnj
5vvEpbdDZhuvZdRsTzGDv1Ze7BUysDvsCAVH9XdpMoWcNoEEwaZ7TmfKLeti59Xs
57/u49stzt1G+uls7U8a75eyt4nUM5afqpqxJQKghHs9OdGQDGccJQDYa/9f2xDA
Nhfo6qYzuOHJNwYm+y6VKSg/yxv4Z+8T6Iy/SrOnNqnEzY1eEGVvy3BpzErSok1K
jtLSUD3B10ztmPb6tTzMmSI3MZWPc0UpGW6Nkp48P7m+UiIMYmoKiMWCrzqW8RkO
veNLzB/1FlZN3umtspkFgQn785KLnRs+HE0nTmoQ3+Z2vbE4aND6PxaVRZlCAKax
+6CTySgvuVgrZi8iVyL9iq9eMcMEtcyiM9Wox2dmPYkT+cwF3EnhISYhI7lzvRve
/py8bTE5h6l8XP2fJi2nWzjWB3ieIkRnjvOWee/dyPm77pODVZMVrmgkz4jchPX/
WYtGtoYmdmwwQ2RfzfakOOMzR8+LDg3nWlRDqhI057XR+pl8y3hYWQaqLzjBJvoA
n6RODkHdzzcAPrs5x1ExbB3E0mbOjEJdVYbOiSu+jxYtiSr12UYfaXQl2SWePyWN
vONbAs5jjx0C3XWz997A5k+CZR7eh4558KAr3pHGY/HssLaULJtWDmhW/5dm8AEX
s7kzd+LW3p9fpidV/oKyxT7oELhwoO877mNxP/ooV4nfWaUivyxUrMhrsh/JAM4L
T5XS9P5p4bb/nDrbryb5WPVUB2cgPDUOEit5Kvvfb27YgpnLTvLHbQaLQjLiXdhf
YlOMUPF9q0V9QyRYf1gMWE7K8iECzNiCfdzdcKkSFdchFQsCowIq4Gl4GwDu4Es2
xUp78Tjc/SbACwUt5NSEzgqVblktcmVWV/gpDmGP/xZ6Tsw40cf3XsfRIc0kI8hZ
VLv1ZflAL8kkG4yUWfKNP7tBAniP4JgCqF7ATsCQjVchoLPYM08GIvLwaBljhWzd
mUZ5IzsAsLZ6t91EaHqRtvrG8A8cf03ScwgrhjiuSRmyQ1jh935/mXRrhkknQvP6
9KEPmDS7khR/Wf74dzMTzi8V23qRElo/9RM/so119roW4qI4v4DiU5j7quJJM6GH
4sRra2RM1hYnbQfs4UAoTqpSpyVgK4Bto47v7De0mt9opqcHfmdY6drNnAGW7zGR
zjmzQcbZI9R5iromPQ4GOqWxWKww8ZAxAOteAwB8QRnMu3PewpS0jld2t3LXpOQz
YZxCyuyUEnKUJKPmSPIexv2PLLPGjoxaaPrViIri4Ovrn2RnKGnaYsSvD7wj5r7N
VfyHtT4QiW/3Y56QkOVOHq4uaHCw9Nu9Y4Ls82sG7J/jD2oyBEUvJ4nXxeAvB0Av
mA94Z2KxKfpiYlkq34u0FIMrcjD4LQuoAM/a9+/mFHXBnGn+uTRtcSzE0FE7OuXm
lEA3h3hTRzhLayqQE6tN4WUlDlz5PK+64mMAjL6jrpwOQYkFbvyGdLfiPMeK2TSP
xSF/0ulEQdNrN21HQvjUXPGs6ebs0zQdBkTXG/PcswsASvyxd1QU/rfM9OztSXyv
tCkP/J3SiNs69yvOT156MGHpNNC1/pgZikn2SEMqtpPHHYArVU9HAvXRJa+vfdQT
TBv7SRu4zDfAIu/mio5znxt3Su0bmQUrbOUgEBl7qIf/d1AkDmbmAxgWnaNW+CAs
CWhS+Nkztupxc3P4eXbUew6gcI9lrgHfRGaA2IC3pJcouVyevV1gOWhgdnNUFpCd
4pRnyN0ahWnDvwdMjZCmy+TrcvHPkHGgMy0TpIBE4BNt19V8XXbRNTVDhInIboxW
u06+V4783/jZlRVnAtYvzRCFXZzPYoOmWi2pe/He8ukpo5JtCa8U8N45MYKLF978
vkWrKw6OYz6PLEaSGcM3ARRa4zU7ZqpnJWFii+Bil+4I+/rXP/ise3YXwTxQtK3Q
2L4i5HQoZa+8Z0KFALYj3dwV/bmBDgx2FOZ/QtGit9Fbbu7xSJbJsZ4yk7HMTHRE
AxR5bONEZDpKHOmwQ3VXhFvwkxHKiJqrAyMpuGJ+uTwyDMdN4G/HOOXO7P8nOWMj
mRpmYJnVPxMzVCq9686p47uhvq6tHwV5+F0CI+PhXRZD2t1K7t4N4JMaUHDUDtPt
9Ek2r0Noa1QlCwZ6YIB/1/4uzZjknRQkDspkQ+k71uueNM7pFjlfIQb/GPkFPfNh
Z6dpXMhmjFRTCU9UyZrX4w75lkL0/ZXLUmPfvJQ5X333PKem2kIh994MHsVrpmoV
y57m6FgKJDkzxKPVtfa1DfBxGq21x2xMoUEZr7QJ8aTbQZiHD9tiFXQsjRGq9Kiq
UVX1olIqgZYq6suJPHL2BCjrg8k//p3qjkd5UHy80FNHjX2VfCz3naF6iwixxsy1
Qnm873eS2PTQa4saOiHxK3I/kEiEsz3HhiQSqrzeq3g1PEs1SRgqoQVh3Sn+cEEy
hfp/vtOlg4mfwxKpUJVlCVCzg1t+mKkxQNNPexLKJ6ttqWZJighBwb6mTuCJiC0i
ajyLCsO04fQ9uBObeBJg+FDiCveq/UqXlDyU3oe4es50Y0A8j/EOveCbAmwZAdSB
9Qna7iGtKYdyWIqcKjNKRmhMqnPZQ2Y1bEuqsyDMh9ytlTo+pLGN+tLchdWk09h2
nBHkQ+DKcsUYSXlhT9fyZwbdIuOfNOIQh+dFhsrNRhf5TSjLn8/q05K8lRGytcqR
b9pGIiutOaK7/icQT1x76ArND2lgMQg9YcYM/dw64AvRU5mYnHPbPrHMh3zBxftC
pu9/Z/a/k9ieu9QVpoUZd2+/iWe+tXCBOUTsz4eLan2l2WStjK7HpWhiTGwSOKnn
3SIde56zrKSVVInmHz1q/6UaHV3cRowGsdMCnayid8z+QmzGASU4BIJD31I5uYga
8Xm6CjZczxpyIFlAwalvQqrojRQZZpgAppkzPJCphwzA4WTALf3AZLFC2tCsKdFZ
hBymX/EgiIBzZNmR3R8BCapnajYsiTQcfzKDEZJFgOrYBespNU4djTB6d3WUUSOE
a8IS41niY56l19Q4fQIe+mWlV79oqvH3hJ6WKwlp7izlBY6tT0p3u4jMjxtSy7Vr
CVa88U1qnVS0AP1cN0fXq9KW/IaTxVxsVXWHIQ2ED8094AXB9JBVVOx1oQghmXmg
zNu2cAonJtL2twMz7AK4whspNxuhwkK6WO4B2AfvcBpXYYFhzvY0LR5TzlDoacQP
5SB/wxogUPFpSpdpGMVHCP/71SrEvizJ1R6yzdFB1wsICbeZxgU1scOSrYMCZNyf
aqtCnWE0QLEVLGRqWLQHhlwx2INvi/63IeDGvaCEE15vkYXNis4CLNazcZZPuatx
1P1KvtRE2sUyKj9BDKPomrhgdsGxWxW6VkqYyklh71MICtpmCVOZ/NHA3r1xuKSX
5JZH+22OWk+0uVR1Wo3v7CDWcwPEb0vfPPG3faoNBqU3orI65kDmqdqKHImATCMr
/M0G1tS2751OUguAbpso5+6yfcBVvPb0KYfs3F3o0vN5aFR2QBIy37rCsGmVUhGx
OFM5Tefud04OLI/PR6YcZYk+psd/dQIJlSF2j19RxXyBiH+1TbDTB+xc+/MnYukr
GY1GYXSkxSIda1KsU1HYhF1x2fnygj2tkT3G/pPAnBlliT/cWkDCQRnu7FeW2LDu
JpVH6FCvdpdj8PXNYFfwNvJ2dTeH5xsPd9luie/RAhdrJ9Wi/ha5jY2LK0GJ1wQo
aj20qCwpHhZ4p4OhcZtDt0tD8+WCfJLMxIGOYRSh1BHYeHsAMDGIoMpmq11lJUBV
aR+YXRaNctH9KBZwBUdrh19oYNw7jeTbLgSb9/pFNo/vxX1dgPFdD1sFeeLbkoi/
nUjKW0CpDsN5wa9AVyTGJnJrbLKsSiP79OycJitkHMf3DBqBplQk3aXVgu782T6O
OYcXwKzuAS+QUnERjO+5YMrztxsuMZExmsh/L8m6XpUSmCle0NDwKbfzj8YQag21
7mYlTwTZBvhXxDeFRGM0rpwPMqse3LwmBKGlY/7OSGB+2dTpsrPOyXPID0I48XRv
1MGcDUXI9stuMNDNLJ337cDieic9yJgnKp4J+UCujuc4ofaxzbh31+yYcatB6A5p
onSy2bxfoVt4tgnSZ/WAcbaW5khzytdGiS3fZg0wds0/VnwBgnbgv0+DT8tjLfqd
HZayuBa8bbEofPkJfqBaIHMcFEtgFJCrx+zbU0GYlLFMaNyOplfW4lCMpygAnq4q
S8WYF34Nke070UhxDYKLENjlXgcxGEo60FDAvId/7w6FN+3jgP1+qq2aMdZm2iXL
v2tUYo8cpB9iTENjtIEM0gZLiUuVgX9yqrjHLK4M6C3wcqRZJ+sUZozC9aYWqfUw
1TpQawoFPmlPgDmCkBQh8sUzGRpT6FErkc9v5Oqo29gyW6uKfNR4quNpWiaiHsqx
I2oLXRb0RI7+5jpUjH3lQ00hjvSFHBke+X1Xouz5mjULSGH/q6ODENb/pJ8qe/bZ
PVF4HrRSZFn4rcub7iGLXe/lskCBVARMMQGjkOfchwd1Kvfu2FiHUGDX2eqwZNbc
O8KFbfrrBtizsvb17bNIOyMYptYpuLxWyvP0JcKQQxmW4w1lYG4KG7Gwig68/eEc
cTa21HGWU3lE+zg21oMTXFOM5sIqMIiIDVVhaCu+mX0C02fg3sDhOD0nwhCBIyVK
Pj0bMz3AfRid6kNdI/pdd8SBbcXraTIMpBl3IC5nK1Ii98IDDIq7qP3m/hzNgklV
qb0rj27/2ZYEA9omoPZUGYTCfI15BfF6mt+JnhW6NRvDIp93V2NHGGO3g9EUb6+9
WPsb6om2L0RPiO13t5G6wUeNv7sX17pgwatzP6pof6843c7CG+BZhxNkUTSSm5kV
h5evzBoEBGtiovqknaJwCZkVSU5XHYH/b1ub75ZGYCe3w2Pq4mHt1Ej4MD2ChSGp
4RAjpeHTBi3nf5VfPEkQdZSSaF5bLDoQPfSo49nHa0LzIiPlTI0ekMgKfaPbaHcV
EYzm/0XZ6Ln6Rj43NVHq2IpB7Ej/HMGk9wxeUxtnMI+RVFIXrNd67KADJH3HRX7U
ZeCKFJEzgc7h2C/AF8zU2v0aF0HvjSy4p0+ek4zGRjhzO+z4oGZ9Bzt+GeAcgdFi
Gs0TejWe+5DSzmihwTaRO/vAOhkThzhjGTuyp0GO9PRn6KPTCcZpPA/z/xM073be
CA5UcUJm2tnnHRJ2cV0mBVMGQEyj2oEYcMJNKVaLfZVTO7R92rLcUHt3qEdu9FaF
bx11aTPP1fy+CzGBSQQFZM19af6XS9TW5BNdLbDcp9ivM9RRkBrMwcw7tFpXDPdj
Zow6X+/QZ6MasXmeYH7CjQqQMcDMxP4h8o2vBvJfhMUelY8prX5sur1F3IuDFq7Q
BN+Vkv5/SiFcsAyP7cw3h6DogPghOuHoNQi6z+tMRKzqirKLuaSnxMJvCsyM03QW
0CRUxh6GXhBTNh017f7xC0yAo0vfX50GdEoS/Ucu+ESbXZGiDCWBQWfatqxb7kAi
q36FQ0vjOyvZsyK7T5WJnlN9QesQIQM7paHVxBKME1dUOD74y9r0dsDtX6rFyS06
jZEvekKG5tf29D1CMlNedHt5/4Y5dHYILvP/idlx7Xbfo/4kbzVxbduh3VDZgx9F
fqoOu/p/DgBUPuG6DqFsDDOMhwH+oxzUA06qJQ4NQEXuqjAqqff3oWs53z7qpGER
l1kQ0v/+Ad0LfZK1Jermmc/93vEyGrCZM+EFEVTDfPB4GhZR1LupbvDmh051rRz3
bkUjLRbxju8pBWNz6h4aNvL3jJgDCuuPoT/PsYVHef++fwK1uvuzS/3Igv9c1WQt
7RKGchUw/ADLjaUVEpmSklvWFPr+nL9bULz2QVZkZWgJrI0YJ79h6+aIfVqfd+hI
nhNfaij7WNzj/Nd7s/CHS8nBN0cNbOuNzo5cMmaHiSFO/l9BtEJ5jCgtN2PNFCox
J7BnzZwl7iGRQ8fk/OFGgJc/2GrMEiuxZLCsqd/Ytw0WyMifkRRQ3ID0bTgJPzv6
FAtyHUxjJc7KHJRzeKoP8+VrYaOJXCp0Jx7ysXZweyjchisZkZFsPsxDN1BdTiss
Uig8ovdSEnofyvl55gi118fXqyPoDstrO19E5jIRc9/O2H9fBSRyfmIHsQs2BfO6
ngqVFR1CyklPI68ZLts+YkkSoe5AKoECEtSdmeQa6IcLalvaF3i45nRihGlB3Yzk
W/S1JYvXx2qyBOBTJPiufGe37l1cgIV4e9FVBwsn8zlJ0uzEHtWyCjEi0SsDTJ/q
Y4TSN5K8iJ6H+BrnHNcjo+IX76WX4G3LgqJvmekF0PpltacnOhTdNozP+Am2NKll
5suf2tHuhHws6CgrfxlM6SWz43DzNSuRE0e3b5j2h4VVvgsk/Z32R3QHOvCbb1mw
/I3U76q6e6TRTYSvX7YLW2k0pVeGF5bITZIqLaotbBfP1FVeKVhxb0uBZ9AoahXL
mJJgFuhc78e/rYXLR1Waw7NrxogqGTnCtV002irA7wpcH52KO24HQD9Lp+6Jh/Fa
vPahZsrj0RgB6rv7GQ2MignQx0t8FdOax4ewZ8aOarqiC1Cwve+7QTyzIWA4MfWX
oztWyLLNb2UAlD2elF+Rs+AyenPJe+Fgkptn8mD/6g24NWDDxFoyNmoUvPnLI1Cy
IJp6MBParksww1g4AByNaOVwunXTRkbW6xyjfW5xZGuTihB8UHTx6MqyX7TZb0YY
P2twBb0czNW8tkcuiSIm3whfoCoqbHX1iXF7KkIdT4+5+z05/KzyJwUl9gvKT86I
7xcu7SXeUWqQp9IJH0LNaGxeVoa7VKmUtsnqe9+KcdeikQCCSwIGXGjpL05WU0G1
cBty+K8+BYc8TNgtAMF5YUJq8GUbkcZ/AtakKLLNTC9B+KKLG3ip/5tYkwoA8Z1l
63ozl4z4C/9oIjB534ZOZZX50hngN8541REB7ky/VoCnP53oq1Skg809QAy/rsQe
PMSXx3NuepUwgtZAEIlpUT3JRUSurJ2MyTspk6M0oh/vMCmsDtKmi7s91PGbUk8I
7k0pJj4rfxafmyMAt+fksSC206lkbMupSaziWXcfcQF7fy53UPMvSdMppwaQzMlG
ENTbT+q7LwAnHRyMqirwzgPjgCn1XEJEX957PCQBitTrQWDw3LRoW3jgM7u99wt9
aHUozZ4gQyP5xl1svsjHYpnABiWX+inPJc6t7f+yR/IwJBl8iO2hRkHxtoIxFnHY
svFxmfUOss3fbsUq1CUgCZPBrXBr9FosVLnfb6CjCZsKK9IjazhtgHoaIVMuG/uf
WqvZYjjeeLp/Egxo56Ws95Z5ydmdxX0ZlF7fT3C+1mz7wDqxvax5bi+0Igy2Ue4n
kpfqzHAxNJMGsmFPIFaVe8nhozU9GzQhflilJvAaECyrlQYaxwnSYPhh3ca44kBr
KO1nk1k3kc7LCRyim/22CwqQbS0WUxkno0TBRzZX157RfD+0fVwwRGlE1oCA0hjG
yCx6Ka7hSt8Vaw4LjuaSzcynLMCB3domzV9NSHQW+Q0XWH/VACLX5wudZ1DkmWlH
1HAYMIPLrsio9JubOTBN31GhSYbIitEFAnCiHjnFkRW0hMHKJPC5L3B3sxudTILF
naIWyicC7IlTTMDlci6KTsSmvk/RS+ku1OxVX+ppFR+sd/6I/VVp8HP7NmANreAC
fiUesYzQwjvxH+vAyUuvojuaWrwknkPxYuyySbMwG6b7LZsky7xGYApIrZ25WaqS
iS5hnDJE5xXY0B0dMYccGElq1xOfVk6haB6szoK6TLFHlKrzMIYYoJsn5cwy42qT
XeSDaXlqlrmCXw4gJu/aNcVdpa76XZ6h86qzKc0wrLLyxPLn/G2O9QM6Y887YHtw
QEKEYbvE7918uqGVzBvaZCInuZHRICPp239+ZKWyG/+2IY8mewCe4esFLPJSFEOd
/vXrAl4mc+KnkTy6Oo1iNkfTlmJsqZK5UYcGujRhfHB9KptvdKyFOjSZt17KidwP
eXHqcVQ5MKU92lVib+RGXGn1d3MEXmIILiQO4zA0aXc2WxmyoeL9K3Fph+29jp53
CdoH2ygIqEDhpLhR05F2gMatkHfVb0tfASfgTmfaVtviDAICnoN1AWzO9P9O7oGW
z/k5LBEqGd/xJrDKRgMNrM7DO+EGRqfE/tTCVzhNMtsX5PppBju8ZlVgYD7zHByX
0eRw8Dzf4DK3+aPSTPPKwVyga08ZIbxCDJjps6SpZukR91Z+cw8Ewf57NEYagfHf
E/8rrTBTSBF1NuoM1H2M5rSVdBwtMihM59R5IU3wtdAOcMHb0RALLCig/XtQouco
SRojPDhPtjXN7wbIRiW9gV/w2DiodYvPedX+04dxxR/GgwDKxw749VCQ1ElPbVh7
V4tt76N8Vcae6o3n98moR6R3FcASJb74dJrd76drlPUb1qgyofVfcq0KtegjQGA1
5kyDfzLoVwLdNHQLtACnkXblUEbnOUzS7EGCXzK6m7eCHLp5pWZ4JZUvLYQ1mKH4
wMcfmbPpsZ/PHAOmOwx5eWaRoLGjJF2neH5bfurVAgdFr+s/OP2Rf7ePaNQDCXyp
VptwY1n7f1piZUo/L7Yi4TMXM0T3oMVPQZZoObTieEJhz6NPNyTFYZbtG2vw1uea
cDbQmMLgqfnhfNc5LQT8QpyZvQRAMy4ah5CO1jeYTJFXC0KK1NDUPz82oD3DexQM
A1cNQX8w7Qpe30bnqiCOdeykTYs0m3xAhyzHtZto7Ei8/S0cUSFpFiANFIS4h5tD
DFHmZsHZPMIXsYtJ5OXM7nbTZOYMbseQ833vN09bscPnPQTw5AreG8uIOJ6doloH
niQ9o/1d1Cn6EF7Or5ATFX5e0TMfymGvOO+wGB64Wggh8Wzb6MYFMyl5Ey3Q1nNy
d3pSYRchysv7IRCCtqXV7Jqg6vs/7WWP5Fl+D0SUjU7UWOZ1Co2wXtCpo6PmQ/YU
9LBvlCg8Nc8WiNdCSzcYU6W/f3hTY5wJBxe3g/tAEDavn6kDtatmhS8tizTBm+Vb
flMu9LOzrxbrIZqaQxMLdRcFVdriNFh7BHUAL1iAoGzKF2oRTUgExoZ8YLly/FeP
zjHjW+G6Ctn53vQbNZ3E5jM4S6gbM367ecHml9lYzRkKR29EoGpf/+Ql3pBGiptV
lggGteTGc1l6pNuZcHOquYzA+jptJYPirQTk+0OzCu6xE52KV980QAHJnIZQ/Chj
Hm+q1bodYZjhCZ+kSVJp0/tunnpyiizb2MWnPItIcsv4sGOvyuAhTdtdEn1k2JuL
3HB9Gv6U5bte8ILZDRwj4pDd4leyd2WqIZipefX4mw7xbGkhQDp+J6yy4WD4TEfE
6lKZkfBi/dr7HCIuoUbzAOVSmpISOMydSELkD8nKuIIV+7DvJONC1bzw0BDSt0+o
XziO+gfWSm1gwri/lhMOW2VS9fMItS9AMBvqj+CCC7iJuFSeILbCrEdAnvot8++Y
PpLe+ZNPW5zFQPCkHMJHTQLi0bbMu2U28ybNBxZz2hWYJifaQzDvTcDesbFHmjVI
0eJzgLsObGOii1bMd71lH9vJgl78+5VlfY+K8b+JD4MXGA+bKCkX9/iatdTBRO3p
PgjymZ7esVNBgVdrVJAZvB7zGQbfzX5Tb98xDwJ4ptfnUGRz5BmWmnCiAVScuySf
UtVMyVe0/NDll1onKvG3mm9pkeFt5COPa9J8vrLJS7aW7UbEwydppDsFIuwvjqGA
QijCUsvwbo+vW5ZPVltACKoF4Eyav9rsRWbVLbOduHKtT+65u4RLo7XuA1WH9BvZ
MYtAD6pODjvd6a/isdUt+WR1VvJd7da0bpU5tC2kL7krv3zFO3SNejmqNaBUZOGa
X8nCWYIbThdd8FBAX0wcEd3qXQVcXc2yTEoK3ihab4ILes7OmeZfFdVNJK2LkLcO
6NpK9AErtbEUB9tUMV/sq0mzhQmuaMe/kUnmJLv9W+a0vHA6S0x8c2V64tBhuM3w
72nPTiPVaHzrz02OpSk4Jcka+w1w87Cnx6LG9tRYgJ3RIREwQbbcZG+4INKbE3Jb
6I+knP29ZAe0Egko0Ap17EHQDXCOzMVoqKjdyva4ariVcbL8mjeWDaHcD/gvHE21
GPIrrhA1xDk3a0ODsmdelmFd7sXP/EBFSHFt6OIop5T+eyMhUz/r69z3NSJ3GjUK
T8ixNzlaOh8B1/6rxCNrPWDMAcSLBN4LjTBhMuN3sfD2KT7xm6eJUY5QGvz0jQZc
kP09JuGmPGizs06jBUmDo/P3sIY5q/CnfRvCMX3xuZ4DIQK7IKhq0SdM25eax0J7
wUB0a7QpP2/bQHBvI+c4PlXhQyFnCLXR5ZYtTQr1Z/t08Dq1kU+cr2IwCePdGvY5
bQlRknBt2fVHRst1TAKaxXL5oqTwaBbk7FPPZPc/SvLjmEvD4ZYHNnSq1qo7/b8X
KNshTMOJjfA5yeMsxPB4JRgBi76/r71lgqYAgBnFKW35WYiNm09p8z+JA8XqCnbF
661r3k5lStysW6urmAZh3YC6Xmi0unM2onvD7dbRcuY59KbPDtUDjuqJQVEdD8/F
gK+J3PNJ0C5a7NjA08V78LIVM1ARQkwiDFwWBIDBcjI+XVZdGjOeGOP9SA5IZOw+
YO0gfhVBVEyem+OS3+PmNAXNbL7EeiLJ+3aBDc2GZ1ui67NWeM+d6vHpbd5ibl4o
uPOKut+kzeBPyiDuJnpN4PdUk6kCY2EuKXJ4zeqXC0wGpzyE3DF93XOjiYVISFOD
X4grRVxH2wMRZZAGH5YVar3hniChSmOXdVSXInOIvTj6ZW9APlFfShptJaQdeghr
bbH+9E5HEJYIy+WmUPnVcI5C/azC1KwO3kFaXoHCq6sAmIpYTMVywkZizLKFR1Jk
e8b+g6o7p8PMpG1SqwMan0fvFKRohsjfs3YdR+HfwI0qdyLcKEpf7oPidVjVAgsN
bVpIBDXCW/UduBieADPnweB+X5cQXonAHGZk1CUjVP0NeoD8ZJdeQ9QQQZlwDxFc
3Naa3Z80cKOo9wD+5TF7cf0SlwYeyn4L/bcsLS9AO/fTgyE0MXm5dMzGmv/pn8mN
w00IrHlN8911Wdwxvaq09nixI6Zs9hEVTjcG0I9E4s1ZrlLetUNVDHO2fLiYQGF0
I5uEutcIu7QU4JsBzIr8n4QYXluWUrrKv6JRreQXMexCQyZCJWtDY/omRCadSrvZ
pnQCodFOTxwOB/glBVnEuLYBgaAeF/XtC5Dcbc4BkTwwfVpemxBsaQZHAZ0DGQ7w
TL2f3+YkiNMZP8F1cmd5+qWdsDma+ZiPjbDNrQjES/Guxz5UzPoAYd2vw7qmpbPZ
L14U95ddZDPY66kvtjpnR5a4TUMhgsnLHjIRyjGeFS0ERfnb6GXA3+7SMtWx48+5
MYqdFzmzHeK0pMaiclsnagiJewEhRj1D41yIRt8spZXniil+2lDN1UNs/MifdMip
j/TvudSy8gAIpKts5MMlycoZCuVtI4Rp5n8yH8MOsvj9U4wgbk9QVeT1qATReZzw
Ifb5AN8+pYBGKg+D/3AKU6astTOzC/URfRuTLvhMDMVRk7M5V5dWGSKzFdrsffKU
f4maK+GZ/O/l1E8cwMv7hQKf9iDHcNDaEGLi+V+RFfDaMEIoChRag4J3hc1Bko/y
25DbC/aIzTd236Shx5sgOrLPqgfyxXv6ATZeJz2gt9r3HzQBxWfzaUAplHGzgdQO
n++5SjYMCQjZ47obWduERdBDAMmjeTfL7ql/2Yi+uTFtmEl68OBo1FKOdFIqLmT1
0Su9nCB0x0HDGmcqaZ3PmZOEcco1DySukO3gObBj4sZOWwc4ML8dSWpphJaDioTm
Gd4c4VYy/39MtQc6/lcSfc0zM8AxOEcF288MvlPIbB7Cb9PCjKVd+pJrugG5iJE/
BbE/2AfGfhslFOv+685IoKA0kHSqAEiTdpr79y056l0wlnXxReKfW9dUVjHbYcV6
TUl3oginNTjEKKonePA8iQvqa6DFnwqh6n6BqB5bMXwQXSj/H/afvqru9St/oNWE
imBjR0qH6uOXSp98VMSQpXqZDHV/dgtgkyxIGX7Mf3FEMJRs0FxRJlqPSv4cCGKv
FUtBrtokPMCyjyT4EGYX9km5+Eevt2RsSptlCnIy/G6hy/c04T+IgjqcXxa8aoTi
iINGbJxGJzVxOzAK5LjUD200j5QjrTbEBGVW5qR1S/IMr0kD1oiqJwTL4cpVxvwx
W8gwq3HxTLI2zPK6fGoaqWnO57I8QCWvHMgZV+5Ki8gG0ehQugJlTBRBLZtfVC0L
I0cq1kYXZu0tBkgWRK7doewu6zAIaE8q5o7Y2GuGD5RR5/uEH5CuUTigT8OjqPrh
T6m8wUdHmT7XM7tET39rHpan6rWiBvP2MKDecyRvOC5LXi0XZYiGCY6hY9+3gf0y
zDDZC9xrVRpA3vo1X9mGr7/BLI6xGfPnRkn6k2UKpN3K86yB4lx9I9tUwDHWUKcI
OhgKFj5n5FPyPOyX8+B/PhmfwW9f7uBPD1yzuP2gHRvCe7UtnL+HZrGPR7vk16XA
jLpqXMHUPSct8rtK0zzDoHmuhF1A91XmVvCRl7kgVscustN1U352Qsz0FGSY2PtX
1VE75AZMiam8Z3fSjC5Gqn8CzBmsHml0+G6YnkPcCDhYOIRFKVz9BVFAZ+kJBeUL
mlYuotaJR2Oxfm3rI90SsJR85ei+ulTPgFD3AAVraNE4zoE2igwMvbp6OH2xRvIN
kioqO1RzXd6ZehfHngjVvKPVZS5D0yVjSe9bEmHB+gMdQrTRoUl+txduDok4MNlz
erSqEdc8CzFE3Jx0XCi2L7J4ln3ZhUYyGIYkI7AAFimjhgds8hFK3DVLia3gPKrK
k3FXRbyHkuTEj/G6SZ706hHArP2iqc8+NInC3tvOOlKtJP2vk+su4dqyMZBcDO16
ieEZUAo0eE5bYOjYRi9RgepAcfpMUS+LGhXJUN77hLdRGsT1y2G/CQaT7eSVs5OA
Uo3TRBC3OMrKyPTdhsHCrRj2XdmVcYqp3zCSqpI/14GconC1QIjiTmyPSUSq35Kb
B7aISL2zq4COxIuAkJLfry9ux18+7VUvBTgjDFridIqZNVQN+CPRNl3vvObFB/8B
0w3YvKg4ZSCvoWsrqiu54fe8s44PJtAWDZkHaElXKipa/K10zfYPm1j/j+m6dpwq
BCz0INA5blZ3ozONbl540BM1/wn13edCiY2Sr2H4OAaDKivU+QcZhXttxctFCpDt
09Lj+MHb8bLS11QFqCtAPm5if5I44xPSjg/noR7XowsfCrisXNz+ZmBUyLAdeeGu
foH5KWCkwbtMv2cdMfMeXHQY3zLtGq94PAmWadN1WqgCzksa0cWeYjeBm3JMTkMp
rXu3kx9f3YRwCvldzRkN72hiVthYIjLNeks/Ck31XneipYioxlZLmL9q+hKqgSIz
SqSaWL0lbqWs0qaBoTsC93siEU75kvnVnPdVlFFuwF7lPhLPtnZzJN+b2Rptwj2e
8ES9FDt/Il1Mc4uxjOrgq106BHj4vL1e3S1ESVCvKDyKCYGCcPthUQ0E1pcBZ0Ld
I51tO+8IPE/lS9aQFY66fxknYxwl38BFORaRCfHhQrFzc3yCzJ0DZrB7S+O0TiHg
l2HhtOD8TDofcr4zWu/an1NEqQornNfNKXelDJyqamnrMJI5w6714/j5FZn+ll1t
HDaFvOI9bXNyFiy3UMJjccD1LfTPxvEpWkcc/JF+gym+E9Eza+q9WDBIRlU7MC8Y
adpQUPHMTsirKrTT7u7OXYURZ+BzO9yjKHp+022c3Zykjn+RsV4T767PiWabXPLF
kdyYJhADCij17+TxyMMRNDYwvdI2r0x5RpxLB9c27Mck4o1ecRXej1LoNWANpYdT
0WMiMhkBRmu5atBjNCC2T5yT1624SYHW8sc5/4QAk8ifUmm6iH39K37k4tulKMol
4FGoy5t7BsEA7yerz1tZgKaK6+JRkXr+FgUmUl7KiOk1lboLjJ1Q6XlUSQBlopfd
GBuVfo0h73RSXGWT6gyqh7qGLhgpHy4LpXKMWvknPtnFCSOTFbJCHd9o3X3fVss2
18j0wjJVsJdHgpYp8eatZT9QZXLL9UDn7h0g0clJfEX0aVylt3RSkx6onJj1xueJ
94sJFMGCCjzB+6Q37MDhBh8MKuJs/A91+T2GTVXFXinFN4BplYpl+4p0WL7wVou1
tc2WnF0CzYonCsgMiEeJs9GgI2K+M+xCFPevX5rbtHZdN57816lr4SdIZzRJWnof
MftYDLJPesCrLT0Aa0OXri+dSeJ20fg3wP+QSnxOF8sM5dl3NBdsrW1XElOwC9oG
M6kYgCaJ20od47EJp4JAs2ZbtO+djMxH095rcgvj2T9+HzLMdVXCiOq1yVVSsH8I
8n9LnUCV8MqFjBInp6ZlDBeljyZpzpyj009a7cR4yo9SzjubMxJG0OBf2MKhjJDq
JpPA1jADgX5FFyvmpCugKpIiD3vwk/CUX4szoZQLPz62ubXsnZl/YxjK5AjFdOL7
1tXhpEKWicpUxqBxj2FByCTVBa57cA/gbrzjnOyRbuITZoUo/cwNxPSoqtKmBh93
4+ez5SVoDpcuJY5WgVleMfij6WKBZ9hUCRjeBQS/T80kbIaJRsGEUTxaG+rXmdki
Oyaz6jEbyQeOGFWGREtocX2Ki3Br0RzF8Pz/qQnvTNkuFQx5lDu3HY/pEjWpufiJ
zgt8uPf/Y8VyvjQZiay7zD+/HBlYUveWIFNHAictQSqdIHloi49opxXbsoWuV885
fFW1RiF0aflheRLCDadX7UdRBG9LFJmqnlZeJLTcHN5RWEBn+uQK242qHxZhJhD4
WCdpEmG1ft50oXMqiFsvUOjnB4A4lAtlZnKY2rKGnSIv9qWglfFwHnMs1h/KLyp4
Yj5cSmAB71WpxFCcZdJ9dcDyHQKaSk1+IcvJ1WgKCL8NvoZm58siDqpROGKlNZsF
DHKX4rpa37wVkYR5W9e43o7CpYnkGz7jSd0Kk4dhna5GBXIbejzRZv5EbGwH6qec
/Qo0tmlzzvF/t9K06Nnv0rPRs6LscqeBf2HeGF0VB5VsKgjWGgqo9qtc/eqzXXhu
JTVvLfxCA/tPdxixx8q5V/0L+JhgbuBsDD3jx/lCNMHeYgWsuF6kJpwC3jvcA0NB
ev+PS5avWKcWRRQ5VIV9PN7PGZ4kdbHfm3zdriw6PgyCIv215ZDjdPR/caPNL3jX
N8X9z6laIF4dLQuO0IRIkRBH3YUUC47QnRt9ia8Qi9yYlgtCf24s8DVJmVJOEGlV
hQv+nup6YEDkudBjIIBHi0fAOWjQVDYOmFDySrvTrVwxR4EVi/4s450efG83viL6
PqIa9Ff6t+vOCOt9pRcARU6grqfVyHuVrepaFE1pNnpRxA/tx+NKOr9dh4uYpgD5
T8pt5PApJEgRSHX22ePOD++rfrW5IShrlDWVuY1UpH0FFC5x2A3H8/mAmrnYYjIQ
+auhUzG8H1xulPet5oqd8phEJ6McM3PKPwR5ch51DJdDuhyvLux2/SQF3w1d4Mri
a+ox1zvVrEBOfVvOZKen2eHLw4BljL/ONxI6MIgJ2hh1mhgo8sj/ZVwi6iuTTUbD
lFvb/IeP0RGRqpXGPeqp1I05Vcb5WyY1Or6ii7fDHsGORtjxso90lfIic9vPaMQs
VwF3svN6uAmLIEiSWZCwNRWnqleuKR2/+lenunNmdZQBlpcRLHq/ofatuAKur3Er
NbZQFq6WWUiZt8yNAwMjovPKZ0uE09A+eR2OkmpYHKU4IF7N6UCNEYaV6Iaw/nHS
UIIhsWhjxRXqoHRgmbp3G4u6bWDIMmnORz+VwmLK0Xc866QN1JmrZk9o15zuFPHn
S7yVPEZOV5i7CrKaNvBjBqFR9KYmncakiWBRc/tdudXSsmU/7vb3OeaoEDmUibcq
dmUufDQAeqosV8bMjRhC+E60CKuAyuiyA53zF0kugYkhl8D21FygvIgJj9+3KG3i
s5jleHzE0V1zYcqu3ua+zLOLOu8te9MavMZU3X9PKmu6/pwJT04QOJPsVrQZcxMG
AdHBwc/Vj40TgrefM7pjCw96yV6cvuR2iabIb4ob2SLCBj+fNIUjOrGVAgRxtLa0
cTOzJV+/k/iOSTimN7yo0GJmTsvQSMJvoExEMgVKidA43ckKyqSLSAZ5YYCxknnE
3bRf+0RzrcLmFJVLVwGmQuOeTmPyq5IT2DF8hn2xJ+j30KYhb8X3hKKhUXWqBMRX
4uzI/E7WvTlQC0wcrh6iOATcH9ENu+XHYgB0trWjTPkcf1K4+QGjKt0Id2eyE8f+
ZKGgLxAJdQukAR01cRiutwzcR/ACnnkBjcbK4cs1wH0RTE9JI1w5a9rHgcXiDDkV
rYxCp+yW5wq4FzrGHn9lmFVy2okoDOftJo8Jsep2iYwT5k9kp007ePSGfxG1k/BC
77aae12ZvzmymqCYElUnECaOm58RpwlVOsEiYbBNujcCRX7Cs3uDPvLnvmHYlDfW
bJ2uyxJP8qxc9Vr5AK0lw1fh7xGEFpDdCVriktsSNJtW404bEawsGv4FWuU0LORk
HZMqmusn6RDfdEzVzXKJqgxYvJp6YIMrGhY1Zp8xQCxXHjqO8v5kfS6pFxNcoW2f
aDYEYT3PbTXa/TZtqzqZgWOdOii2SjHE3XvcIiUJVBFi6W+ABq4Qr0jcE9Cj3SQR
asnhC0TffwZ5EnOxtfOjyec+Ne8Kdd1uFiFCDkXVNDWy79K0jZH+UPjuQDrRulvk
HdAZ1+7snAFbmbsM8M0lKNqQCyWPeSLhr2EvzDH+OrYodzhClmGcOKz5FtAPYNFf
7f/gXqlWDNYBo7REXMBrPXNDg6YvVEspTjg6LrwUP3b4YQXFmztWCwW4BjczA2eX
OiG87HE6UiMTA15Vi8HSw7EhpJJcTASbt8KlB8VhL+gIiUbgMJJ7Ytl7HJiORzH6
ILd0IRuNKn6DGFEYFaV8GqqndqyPXBtWBybI3eYqS3Ab14ofAP+fNB5vHAVFbck0
GIMEvocDEK6OMpnMW/pfGMYAzivKCQWERT3pMdv8PQccrGHqPNtPZYWm0t74R2vj
WI6l0qPprfQTnEf8wlSweSuZoDMKIMDJBbnX6SvWdc+VLk5kPxA3unWxLQusEbZk
XBvKgTIdx2JOr8nypU/uNr0evBJOgvdzJ+y0ZQy+SMhoZzyEAJ+c/cBOFmiukOiw
AZoX4Thzw2suXWiBEom78V0E/2ppKfn4x3+5pA14CmRE3WP8kd72j9xdWDL6Gvwj
fhbj853oNoT7WOCAlUHbRznkldyIZ9dQbgG0LCtaPb86yPtZoH/e3+mrPU2p7qyP
Yw2tFM6iry1bGxd/EGd1eZGndZOb7kY5SAXIbaYF41yKrklrp0mEAv6FP7VM2uWk
S0RhmoutNvEpKqSqfMayDNvdL9w1cO38+gCB3f/2reuVyRQTtu9L3oo3p+6nXo3R
wbtB7lgM4mUbdzQq9yRUAM2ps6zty5iZwxx1Llkj52gMvTz/4rzxzgYeaevLBeXN
NISEFFhYP2KCdk843V2cwbnpD3lnDmQAUxYgW0FkT4phAlJC/nH5/tHjFmB3Kexa
uCbZ0mkbvDzUWgxaq95PwO0UAuw577A5f8qzJ7a+ZJ+8QMfL1UtYOaqiAhTryO0E
pee5TW4tksXbaUemfXOX2MDkMRUJLjf/WJgKDgvskUO1b6Vdm66mdhXiG5U5dBxE
mGUIrfseG/wyLjuBCPJTVEkQAVMB2166CdRIWzazqE178rQDaxoU1vzus2F7e6/G
HE9B4yQY8pAueVALKsQAvVrI2luz3T0/+9Xb1szC0kHiTiUQFqQ9OCw2d590DMrC
E/Wh4OG8AOzzefl7d3+HgVeBURcwiQEJNyZkbzEDB4L+LGIUnaWiGs97tWNrmuV/
7lC6+PklWvFNezOh/4IwPeluQTtL/6kqR6DjTvCoG1UUbm0hWkjKFIsPXKvwlGT6
avORKMlt2/L4qiplDvQ6aEnCaYbpub8xYtqZdvbDqjA7Bp10p8W3cT8gMPWi3Ae7
Ezd+lhAY3pkGM/PniiUs8TllUWHN63qvV0aH2OwniAw9StOQT7aDMB+03bCfqkox
7W3oAxF7I7WbaKJnh6ZT6jWYvc/RvX6uOIOKiyb4KpyqF+ug0C5EFmd8cWO/znov
ujx+EXZJvZsS3pFe3KnD7vlPqknG8nspM0gAGecCiaSSTnUU/VvJk8yu0+QeX+O8
dYkQ859vp/RHDddn2n6bfCN85rdjnJI+rgPZGpgCfWztBKdrKpUzfSTdpAeTwTkp
c+yjcA9GWsXMiDU7MIGoLFWw5cJzKBWfBhzIpO6RC4FiR3vUzmh1LUn+pg0s9DLj
wFBdjDp4GGi4ocWDl455vg344ndXr1Cjy536zj6IF3Vxks4uyynIhxwXLkUPb4gU
EsaYIkm61CeIWfoW1YnfRI+MBNPR9X/1SNwUuyJnt0/HUIwQshXOLauCVeD+er/M
S4LAh/FyOC3NJYcHebIbZNr8wXX6BkCcHVq8tYapMRv+yKhmlSJGorej1VuJyTV3
rPAjVclkkDoYrwHUXPNcEEotoUumLnzmlW5M43fBJG4kon6qWfImrA4eCVo++YMV
Cya/5z3/WRH9xY+cUtSCFBTzfgjAiAO+QVwjOZq9N0de8yfqLkQL21sEnWbXxU3/
aKYigT+SVZ5PQlqCrlPE6hOZnEaELprh8jR1DwBGPj2jJaWEYoYNPmyjTTGRC0WL
JxebXxq2SqszbE+E6U4Kh8Ahcou7A0qG/qxr3HxuIrtNIouyDI6iU2lokcU878Tm
KJ8aKmMDrXReZHF56qERac/ePLAX0ckQYY5OOXAx7ic8atJb4EAiEOmjWEq/N2t7
C1fJwRZ8kl/xo3QZjn7Mi/mbctMvWz37d2KWH0zrjHMF0RDfpK3502QaW7VFimN+
g16sWXLJg3PuD+XAIeb23ZmNxB0CHfL3Legdlh30MOo3R3Y1SyseIs66zbdIBjLL
oZsTPo3RrsKOmy6XgTirLXWj4poDD978T+W1zScRmoaLauGG66QmFU/Lvvf27ixI
UefTJeY9TvIbG+3e6uqFU1eSFEYwriShuIzotMl4+Q3yGM1+ZGEVlX/qrCaGSA6w
LtgDE5arqGbUkbxXKzZ/rHi1Mi5wABGMh1mCMtriUypzIPMBDkBvdEA/exw8B4NN
7vRQ2UvwNvoiSciIU4yJ6rgkFfZ6Bwne0eAXCCEaIB8qeZg8HbPVVM7Ghk2BekXN
wyZX3nWEZz7P07IwVzfLDrcjPdnwG9wTVc5O10VWaoadt5tagcHQD/DtOXOW3YAk
qI4ff4+Bevs4qsxillm0myYssr4H1nJ2iQOHkXNDs7VMhm7ZFILBb9auU+L4tsb6
b/Nol6w2h+mZxo40oQIn0pXqZYQP4B6Pw6OQsd/8lrGUGcU7QseRjLUtyP6j0srX
O/2qbvTe6cSBxk9r+rjmVJmWlF4EFd931zzUf+073WYPFl+zusU6y0O7V81dp0Kd
n0m/WIz7qJXXkUqLKS4Kt7m6AoNXRL7zY9NwZyP3/MucW17DKccgCku5LX6168dN
qxktNfy8Ejdy3gOjUc31EBhQDRGM5owE1kmISIhlWXozTc5AFTG1GYwGP/MkS+8h
MHwCXFv1kObOutfqM9BXXlSrmoIDTcOAVUtKN4vv0U0Yd4lY2IwwSJrhoi5BktsH
PfoIgTo22iptp5sL3W/shNLffs1HXgkzkzlLGjUN9mY/zdCnQn0jANr30czUuihX
77OIioD/SAHdCKyR0DjmBOt5cbqfnzOB4gFLFsYNb4RM9NqkNBP+MNyC3h8OiWYB
UpX2HBns4iZjpbPclBBRv7eQkJaT/WRFcMp41s0BjM2+xZy6D2ep+Vi73hDEjhPc
ADECcI6/7jzBEqcEmtTsjChZpfsr8+OOgCEVsamDZVY5PBW4TDQKzNn4uyMJQqht
hKw13lZo6jy7CBS19M/PGz2CU/nUXwx6XVmNvsU99HZwIccS6f+4PmLNqwMdWmGK
EX/51hTpAhCp2kncW174XxYQXQujScVZossOprceuhq/m9AWfthyEWl1/zzMgH+O
iKb+ugkGQcCHwyHqPL2BvvFt/TQaRXdN1Rh44F+tGHeWBk1zneUqey3t6MMANKrV
fWdA1k+hoo4Wk0eaJNuHcRqA4tplsBJMa5fdl57cVG1IkBoowvPWz3USe/1yQtt/
+TvL+TLMK27ZYCpowHZYoaZYchPkYDIPG46Cr1+5x8ME+KgZ+pAIb6Zg96tg0fv6
leIstUL+MvYe++PpcuoZeVfrn2ztfig84XHizNKuTabtymcmjlTpD1aUfCrMsACB
E/Il/yTrW6Y0TghzxL/cxskvIRKxFhRHw5zfmAzb3OrFT8jEIXchY1ZfjM4rkPMV
s+q7TzTl0t2fyjAjI7DcICVGhy54Zj9d3Fen27TDNZBMv3ArQ9k07N4ix6NzKGVq
l1HL4Uw1u3Zow8C6i0mrUw63vbp2194etoG+eud+cq15yBAR/p3NWYyfUB5WNOkg
RjgflMXAiWIz2ISCXdwrcpY75XFIf4twBhPPOrKuFsSRBqkBlQySroe0LncynsXX
dU8lwi+kM7oFYjUTgaOhbH+8kbOOvbmO3cRsnIevgBQmWPF8W2kiCsFACRG6VfN5
Wq31UkVptKcrOe6bBkdm4oQwHv7RT+z/cgXbWgTVqIJcIDw11TQMQowms0SB5QYS
QQcz6JiphgiCjp1evUV2SCej9vo/y0KXqoj091M/gKKrV1O8mEgJ4gmgi1lJsj9P
jy6mRq2+vZogw/LJjilc9VIcmrq/5uQgv2Tq9ywyDsS2HbDMLKGpc7asc5TJYpwt
6aNBG3uEpeAUI8ekpe/f6R8TkABsQZ/jEUoBrYqE3hyNIb/ziEBtvvqATV3wO9VY
aMdtj+lM3AXX8IRkU1XxYw+NOY+YAgZQeGKYY3iplXeHappEor9WUtjMYJoilk81
zSlM7d3VBrSdi2vH6AjeatfuK0BcgIQ1zSflFhDlRThkRYe2cqdklrBKDelrar5j
mGF2x4fmJgSSz4BE6XM66wJaHhv4824ZBpKeRRMz0FHLq3ZEdErrlqCuUKTnZm7Y
gOskRyG0GGmYpGCIObgG4IhAWQTTVb51q5nQ3yAZ4zC0wS7Y6diAC3ZojrdnQcHO
0Mgjn9/IGotBO1NqXcBHCqaVrzhLFZNVVvl4bocI9WYq8xBwfItypwaTU2tWG9xZ
qVXtWPcHKOARwo+J044KQUjEBkzO67h49AbbFR5T5mwYDK87da0d0WNYWx7DtZW9
6nqpsodT+lhXs7xjKr4bdbPCAVN9SsyH6APyxEYmcdPPmwIf+4XXGDB0QkQuvz4z
9kr7BFfGO7bYtQ3QWUELrkZu+wIuAe9d4MzGfhKAkcwJ+wAZNBe7jI0u1iLtBrEj
aiowIPW3WVVV+679EMF9UYYEhH7UXEgMRZfQ2S3sOFf06BWOtxs2xofGtDqqXHxx
lrF9NcE3WkuwcjSJErQMNJjCLnvx8Mq9tGA/dVqt0D5xhUb5EMDSdfHuscjJAwkR
zYrCPQzSXM4o5Bq+vBa1SoCrokt5NsAVnE4qoEhL1e2uhXd1FVsfIuvdzIb0vjLu
RArQbSJDHRlKjne8dLrLw4+5hK/F4YnAfhAbWBEfHWC5vJV/X25oPuX6mhy4PdL6
fGoNaZipnE7+M7MNwvfD3ssJ9OmtG9N9cFVskDPv+GOi/8Lpfg0KOWM7scU6Y7y6
vpN1WzX/6uHfX5Ohdd49cgwyX3p3+VqFEA8ErZyYpxcuawnEMNk12LzwKGd7g5C9
a5W+c65cTbMEDzGugtxR4K8Ov6rZ+yDrzQYzKVVHv5f7ZLUktcPhuAP1di81ZYr4
nsiglF6vDcrTBW3fkOwcMnoZP7UEorM05d9tIVav1YPrpkBoLQA16MFUIHX2h+TR
fs3EWYgip9oPjwAlrRxm6RRhtBDl0ymEutPPiBQZm77asm6PsttqKG17l4oQprTi
04GnhuZhn2eLT05W7BcaF0OHd/JEu/7sZbeQEhaY0fek0CpJHGgYnufqh4t+yRRk
n6AGptOAKvmDMS8gBY4qWZ4k4/7YIIXPzLWgC6xZYpw3IjIr0WE/SRU1TamE14P5
Pjegh223hyLtVc1lfJVVXE/GUpganoIYCwBNwfXYIp6IwXFOdFeQX41nw82P0tCY
gvgCC+rqPWLy/XH7zj3CiPxoBR32wjABaj8wli4AwJwcYwztGrC35fD8zmFdfhG6
Zpnt2JTs/WxkK9c9U+h+E669qhFRARyuQN2EZueRVNLFXPKYt396xOnwMrtuKREo
4vAdPFVxs/DVjLZqjtbFcdv9zicAJuXxONx5BepqTaJCPJ6uwBkMYFJirMe80V72
5gAQhl/LhLKQXee5bZlN32fx8K5xUPex4q+Jcv8krCQbLvcDI8eg8P2+21mn4wl2
pzVbi1t0C0SxvYqngYY7SUAC/Y5Az5VuNN2re4Wlhf8o4kq7UIvZNFvx5nyKddgG
rjtQvpQMJseA+zW1NQnvrwfEUrKsiTThQPKOfpr71o8pSEtYb2/ET72vXIIjZ8K+
2mwcC96bkxXeaJbCDCiIKqVSQMeV8bT9Vh1u8ffUStUWBNTFFjw1BYx+krRkQyT1
CJW+LbOcoddcWxdO39WDerqygWxoH6t9750qfQgLMoBw+fnKawP/3h8woZvVMRO7
iHHL7adsR9+6/heAb2IQxVYVCifl7PBTWSa3C1vf9E4LQmBS+zcXZiLJ+hPf4f7w
0CrRByHL6b8khF1w6u2L1x4n8nTJVyin52M58jOI6dNSrMpDF1jy7ln+ZmILbdAI
Zfm/NG7gDJb77QmPRFx8d30GZ0OT7GBpjvB82iYbH14Zu5kfWGdYzCXKcOp+CKf4
NYwj/qC7erlLoiixuaXQGLTq0uNMVtkxKWPJgO6ukdR0lICvYtDqS1C44syM5K2M
mhKcJqDcjg2TQl564pVGknrl99nA7lOqwtg/8NcG0575DT16IV3QyeRsBh6dHNOD
O4iPYrnhI0Vpi3Pa5wGE5gBFl3mah+yfwGv9ZAcUtlubCxhXbGh7w67ZllxBrr+X
cwUui0q1Vq5WeW7HWLtKtUub88yIIzHRmOE7SQzBUNCd7iuG04nHj0hd4tRB4Qn/
+jhOqGD/0buUsCqrEP1ijfL6XMtzWgXzgtfB5LxfqEqLjhrp3xNrNQ0Au+1fAvnC
XNYjjivZ43Dk4azEBhAZB/evs+mGbV8LHmTlUHKvjd9O0NuyeZeEX7JdeC65coJ0
9QJLNn3qA5ZzE8SycEq9bkeXML6XDsaILMqB1p3Cy8Dfit27/OF39PMrcpGnwgpB
vRMe4lZUdLOpGOtytTTtmKvMhI6ANiSMTWrTZlWj8aW8uFSJuFWhsoNlGmkcSJoD
xSnN9xLPCkNxipFV4ClLomj4Kk5myRSGCWcorVJtKjcl4HcBGvDxs73FLiuKzn1j
AKcm+MxmnRl79yVzu38bvlpUwgcOPCuCrT/cvgUgwY4GNVWADY9Mh2Qwt0YyRTAk
0yXHZ5rpsH3IyTQA1XoU3bKRxlDhJzA9GtQmd9Kyqd8knvSST1niSUrC4e4YLlWk
z2KfFHgWghkQB5RPgk4D2gOIGpmN+UYhJ8csq9eQM630vEFWWHWgeIKsM2zIK8ND
yVMM0zfi1BsgGQL+KaqIJsIDEetv2vs6UJ/7NwD5QEe2Mu2bjxx2Mceru2vQZJE1
mqivrWP9ASpRdAHJXkV2yfFTfTsEEOF40qvRve4Qm6/JwXMgfFvYVDPV3BtM5auZ
3oNeESEVnKq23ajo5w+UCyQf0m/JZNEisEUB4ia/VMO9S335EBHIK6uEOZnqdIAw
s+FAGQPowt6ko4y7Cx/5gATC1ZQlvxEivu3wzqMEiVEdUnK8saRdiIgY7lpUOB9S
+H1NgAF27he4tUPwILmlZ18ll6i6Oe4jZvNRx62HGI9XPJUONQjlStxTowBmkXre
10NgH2VvQ9NP3ee7kTadaPYgw+kuK0n9D1HHlt8UUI30nYZSLW5ejQjNZXIcjf1T
qvsGujTk/Xvvn183WyBncx2NYGe5TuwLld591RILTuiEBVOZ/eQ6Szn0X9tIvOhw
iE6e9i7oSQgfUvmS8jdONa5ZdPcV72Dhcw/FRLY9qjzyslxu8bgzCFGDtSLf0R+m
vxn+PlaZ1/Bs6FhWc7NDJ3v7JundfQx6FONurMpObwMNxaxfW4FhaIUfgUbg4PdN
i9eaNNetWRN2FBYDfX7HRAgO8HdqD4EJSdadvP/5POlsOhXZNpwMLLFwj/AWvCem
vP6+Hh/OrO72iMEsHuMdaXoZf/rhtCAHbpFNm8CnKpoDBnOuYzBGyWJYs3WPzLb+
f4F08U2rp35I4ozPTK2lcvO7clv86576cXeEmDTMMgvDqI/B2P8yYiE9nhkcLOQv
2IxWb/3FNp5XW7+ig6ypipOzr9GW7FJ4KWNN2xhKw/UlViE9VNGOxngISgAL1MmW
vskDcZ8FAUy3xr2Tl6Hp2v9gczWJFB8HYoqUJa69ajKgUZm1IjgiwP7EKabI9gtN
Lov505VMSuteKKjCcAogAFRSuonLWg0PqL1ykxlbDMf4xCwstRfmFDHtCtL3AUDG
i+mz2dDsYOPUHVcHxMnGISLEUqIXVjWLmanRI7RG4TQYBf0yNzKKUgKWgD6+WTKQ
BgrPI7BURqNepjACCc+DeiuwDZCzRYkFL7mfBIvRlVK5EB1zrVKpijRmyCO/ybco
Luto8eUMPt5PF/qe/+VKcsB/gcFT2U9S3mU1tWYrg+D9kdOOnpbR/RfEKmeq8pVX
NueeDizmCtB23wNrH0ytrWGqNvcM0ChPhvL9Aq2QuLr77Jw20BKE6a2pAbJyYyIZ
nTT4cykLBff9D0NL+IsX19yZL/RUprcEXrikJtawh8Vb/OEt/jSj7YRcOxO/FxgI
jlstNNh8liZuxerqYM0g8LtQv5CFqCZ7T4ULVf/CC8nPjoWtl7sfyWKn/fJEYXL1
SGj1UgcJmzU7A6KWLQ9SMGnqtnYXW8v4nwOrOkpE3RX0OVJ2n6/cFAjWG0D2jKDF
gvrQy600/bnOHiqbg0kSDi+wkVutN8FX2KHeFBTNg2IbB7RIWo5i//LdKIoQug86
skEygf2BtwXskKsFJMkqxZBUpCFvU7tfFxGQ3CWypJnYY1IwXaVs2njHCYrGesdT
bxXE2mvtiFCGyE8dyKhEc5PUYFrUvG5fyX1ek6G+n67piyLsPbNgewVtI3iNs0SU
qeRasYUv9sji0EX5byvSrPq4h0RJcca1Kt2hIPjWKeLu5vvzvEFiSWn1rbrEEldi
mod06TRS2XnrwwX5T1JO5yIV0+sUjk45RwJuu4tYEi8azchmRWibpX/9TRruiQfe
68nflwIbzSg5ae143RiaPcJuPzFnVEFHew6DRwlqaxN8dXTWPHqFq9fzlbTzBz5y
FBQy1pAMTPwy2f8f2S26Iha8/3w6BktShCqw8KekCZjt1OqkNKfEVKeMWbLlYKYJ
boz8JttitYVaRlAgcSObQv4urDiyCsYdYKdjz9gvohT88RjdHkO2OeoEyVo3HXqG
4NxT8TUQtGbbia497/CQGOVYSWmgLRZZZpX94lw7WVvj1LAf1QPPv5o+PtJ19/zw
O9CuYeKPVi4/RPr05rdV9OANPXSULJ+GAOyn0GI+vOTqx2Rr1hBCAJsp5o4tEzZP
2NUmF/4XboDp9KO+0+KthuxGON/WDEj/Hx18LR7iM8Jy55heKHoUi5il1CNPnavU
wnmENIQoxT2ls1h1aU7ueCoZ5zDGFa463lI/7eL/kTf4ekF+IsktQQ4AQKyaHDrX
iTY8MFAMd2zPG4pnZcmu2jHJUfEnXPfzbGVw9X/yMJOrdvjxbCj8pER/JHDNdXCG
TE13oas+gIN7YfuvQQ0SWc4yH9Ke11no8XB1cRRwJ+iASiuofT6AjheZeM8j3F5t
GbC7ex5aRgqciYRDpy+ZtgiNXEDH+RxN75TlGFHci9TteZ0yPM1L6B3afOSuafSy
iv0idITKO0apQtSiii8luH6cqIlRR20LY9Ze40UPOu4PFse8l9G7dt1wOiYQD2C/
7apsQtsne76AV7g1/ffob25X9iKK61+AFO1EzrxuaObbUqWqnkRJ7Bqt1JQjsaWB
0r3jfi3o8YzS8jD3brYb6suwkmbhh9EQ7DupR6MhAugi22MT+gywcuGOQiw4u/Dn
3PcuL3zGoj+5BDLeDUsTjaG3hkRu7RBxLOVi2ZxmT5l9UhI/a6T4o7jVwPNJYzv5
tMl48tPHqgIghmM/xGHa+oaZjCLx0pZ9H5liGFZ+sGnacLV2Yp8/HvJQqXNoWp5w
mdWtlON6dXZNspKW08yN1dVA77q4tMnpU9nmlWOdOptiE1hbl8iHnrL9fMX6GAif
GalWlZychVhIcUdkvAznIwAx6Yf/RFx/UiMVaV7hmncOUARi9M9C90bTQ9UZBnMF
av6h8FeTvNuF9S6x/IFqaSYcvenMU5gwVsNYQfJ7i5WRRsu10DtKKopuo7gh5q2D
3GKnGo49Gy45XMKwL9hrpyW5+B53SnAiWTZumsmXNCnDsEPaBr9mHvN8OcYecDnj
Pre01iLTs0xaDazglMUcDowTrNwXe4nTJ2oTuABxvWuMaXDRywEL9qkvPhzJX9Yz
KYMaERD7aOwBAxL+OLfve8dKMr0J7shtUSYlygdhWdXq+PNYhAq1cz+bnB1tqVQi
UHnU1VDdTP7dkMhtAa96W89ZopmOIo0X9F6Fpts6v6Hdj9zjf9gf9OqYqTR8ucJe
V3l8/JPbm1kUsUxdIGkmzCok2BI5vD7h7m+s+Ss4Y7iRDWuKWjggkF+FZ2r5No6k
btMNF209JMGuTPpaJdgmgNgXxaW/fNgNGQqBC8FwgKU3jfRvkwbnFebZljEND9LF
0ikUdduRZHaZwR9ld6bK1QN86Ko0GmmRbAixMz52bE6Y+nsFM5G/xhn5r3Jg7asZ
hgbCsSaWyQvV9pG7gIAzMkuxXZDlqWxYbyxuCA5Kg1NhL+WOVU4uFxl+COKr91FE
BRYC/z0EDwYQWogdlPdtKHBriVOUiZuRL8tSsZiNFcLOO48INRv350/0n5qzbFEe
W0Xn3PjNcCIShVHOlc0F3F+x2La6ot6ewpLCnsyaveG0u/ki9Dy1VPN9GuB5rPtb
KR6XNpR8QW57psWA+NsMj4CTXDdQFcO/6EahiCMMqN6BVi9HbWlIr7SX99qTCLpt
e1J6hKe8eJGSrXJybKwaSkL3StqUNOHVmuVRLrrpbl8LxbybXPNyVZFOYbFp8iJm
/igWzETyll+Dd2GzYSZTOM+RU350enaBFvHrsQku9fm002tWCKLSPBgSCd/ZQroz
61RouLtjWuUyBjcdL5xPNjBcbhQcJ6jpIEYZGAS1E9a0WtzQTx6HEJK6PWsYhLsa
JmyezKAIgnRPt8ksyKZe6Ejyv1idWaq5iecEpaPPlKcq7aPcDK302pna4Qx+cK9O
jNSxa1QuHVBiLTyB93qY+vHpac+cf/yPv6T2MiwBBAm9WKDSpyZWwwG/xhbA4lcE
tawhW3etw8F3liqxchhBT1wqk72LLicBQJfuLF2aAZi0ldeOaH4sLcVqPZN7osRW
Nxiw4lCOBHfMhBOKKO5TCbb2Qh/HW0SIjAY98oHGyXBBRkHSJGJlmIyp/20k17No
jGh2eq53jhU7Ga35cN89dCq9nLNT7Bn4Klme+SqmJ6iEjPCyKLDSpZZuflnt2uZ2
4bWEXKLtvYyD+MJbAQ1a/4tDpNORrzVPELbtjPYklxf/oS78DL8Urm4yIokzQtVe
O2oD6zL9pskcLBF9nzo1pRZtBwNVYUBVTmWf34kk/h3cIS8PcFYLDv/FKPOYmdgB
yhF1H3ptT2r0TgYJVApDvqn9yKHPLAoq6qPdn9sh81sFJcJJf2yEHv26G7QSyU9y
9oIGUpxg8JjAVlZIKtHNw5y5wOg4R52aqrfQESWqn+/M7l6NAMr3+xyIpxZlomBq
J0Hp2YO/K+mug/E6oxYnbknWP4gfbzsUJI6SeZjedcm1wqU11YmO4avU30PZrDe2
OVCANr8Sf+BvGsmvsPtdR94RuI7ejLRlMwZXJqjHt9HBMW8EhrYX+M51OX1Iyn7t
Tv5gHLSBzxugnSYp4eOkrpD8OIvgPsW0pue0clynmrKBIcNR4u0OjsfvcHvGCRBy
F/lcKJ5C3YwsaaodxrmWfS4x531UnQ+QR+KG0eGhbiXDxFDXhPHKil2JayZ0K2e9
UzmjFVMSphUVg90JN0+5oKCosRrEf4zO+8pfmwEn4ZO+b0n3xGoIMrNmoYwCgA1A
xvIYy/PfdOLFsDsxFizLDkodjCAidsuJ+AiTvgBBs8+88jiUeoidXW74v9bX3T7I
8alcYaMbYapEMGgDQajPDxtOhUgDa95yky7LngKybWTKM4gJ0vcUNbfENFeNxJxb
ZjBZMUFvuLK5EpNmeZVjpebLt4/fOny4FucooyHxs7sv384gzyLbowK0ubs4Tohy
ld+WUKcAPliVMhazZLKc9EjJso4D3kyChqanbsg4sc2DiamExY2a2Fut17OzOApF
oX1+l0cj9y2xJAlqwfQbgtKLP8z9CqsdBJ/WTAP1Mu89iQJkblwQC7C/QkspZ79W
G9W0yZyqd0V6IUenkGmJWG50KFLdKgyuBNS//+Sff+ZbefxJEk2TY/WUBGQab8x5
lAW6cUWQICTDJ5EiaKJ8gtkj6NPxEppSZX/gdSU81DSH1Rw1YraCSmp3vFXmx11h
jOMkKBsVkh6MqefFhuoLlVUkj4EMNl+aC3xHaEUm5xsnS1RwMcBHb2CigLT4Q6Yh
ih+jGUs9GPfU/fNEbvUv8JW7COnoVdKBQfBRGm37WuSIPCYtmS7RGB7vUriYF2Tc
f9Vg0Un36D6qzgMH5gP3U4t3rk89iZNtnvxBdBqkmIabq5oSJCvZ9zZrlm9Xp9FT
GFko/uZqUAWxH+XYKMetbsLgX6wRgdwPzeJOJt0Asna6WCqfCt/kdRRU6nE4DebG
NyBjplJsOuo3Xfm8agJI0iVlEa+qyWy5ezPu4pYE6lFXHiMJHSW/CJZGieJ6HZ3f
rDMYRy2eFA+mEHZXAO/I7GnMtLTAT+OZKxAT4TgtDX8cB5pI3BgyU9GK5axJdL5Q
stgVqsYoVejgYoS6jHKyRXKDydI6/igTtb5dJxKN/x8gOLt4qDHUZeZp3FEF3zrB
+zzH8kYB/j7/UsuVQShBZO74Ye8aP7/kC0dDS1yavcy0X7BKRfi1gYA82+CiuNtH
eUAuMHHRwnp4FFZ2oJdIlbEr5y3/j83edxoeRVkHApTfiIn8OmFWionIfjWRCskX
2JbUhJfOsoIwDFD3LLKTyImd9oSxDUHuMYWFjabGxZT1wB8a6DSdm8PdYxIVJ2/I
yyvmmbFupt0UifftD3HpJd0c8YQYVR7UK0kho2zQsVA0bjhxD7WzCz0AC6vkqmb+
CjAl+jjc6mB30R1WL9ARnGrZQQkn7qbLzr/bof8mY7TZcnEJo3CCvKCHX+53G87K
S2df5+WZL3ljnAXAc90QoAfLMfLAXgZOJKUNYapUQgPBfdp2nNPpJD2e+iLTt4wR
GQ5WeAcEUU9ZqGh9TbczqsNp+viKHpHyAGhB5kUXPXZjmNpUXK7tPwz9fw2zfy/8
cIexskCZqv9tFaJlu4muo/Pp4rWjtoHeQcpbe4OmP8kjMSeeXp3upc1gVkjQ/UGs
ISFqvCixXHFEXcje7pJwzEe9RjjDxr6O6mkkiroK/uckoCBNgwSDKs+buJcyrbtH
ymBLzkBwvrPCHf0XtwereBaWMXsMg/6hlJUTMM3+JWWs8grpvNP3Yw4tjie6cOiV
Ozil2QUdFkqHdGbQn3wE8kP0lDWDQbiXhxQIy2g56wqIm+uohRMe7i0RdYDZBiY2
0/xo1uDptNMKYMtbE0cnRcaCVS3fqkpkW1CM/vEi2vVMgd5nXenSlHO/WVZj99k7
uF86lqDS4gzIJszyRtNNUOt1Rv8tUfv393YkE2DRtZBmXKoIG40VtOvyz4dwetrx
7HGiNADjJXFqvTkcCPbua6i30t+bhUSO0GAGLxOkY2HNNUE/PU19vQF1JPt/TOMw
o4uhMz6OPQ8+h7IxphJcGuoa+EfWw92FivRf3eYiRghLwq6nODuI0w5nmvPmDKRM
djSJMFYW5JyDFwE8Hcu59mYGUOhaLTOIkNpxvyBC52BBs6dkxLd43u43EH5excPB
tPfAthUKVc6RQeDa+d4A5KignNGzEQMPftLx4WqLdgZL+qixUk1Yk9SYdiY7Nmgc
4mgP638vrhNJczyM7G6MU3XFF1tNjXEHQN4v30uVaqPwLuF7fDeslt4O7ouNNPGx
RLtxhTupK5SUC9DZfDEfD2RFgXPKDT8iBSVOMbN80Wk/+Evqpfk+8a5Tb7YiCH7a
q8NGrSEOJS5M4YX0vD/+1FRO6pnvNlj6VY28Pwnr3R61v8iKshCJkx9lqGkCYPq8
ZAiCPNOIgDKStVz31UWAZhj0og107v8PJtFWyXJhiBj1mrgi0S7wCGzH2tdk6ezl
t83W2peX61LpR7PuFZzLicw5OP5fEY51x3oCf9nQPKQ07k7PxUqufo3UehF3x0mG
Q/m+NQ7F00XPNpTh9dpGvQuhaJs/isoBXVFLyK3M5V1bBpDZNDIeHNKxzWbNzKK0
63TcKf+OEd9QCe6tbxc25pT/PG4HLoDkVa/nyeH4AM1iAMHJ1v0iWw40zaVb+TOn
zo/W6wpmQd+Vc73xs3M6MUiSuw/b2/IYCdl66agWHnc3S/i+hDEg89xVHNHHG2In
XT2l07mi8IbuILCkFb1ulg8pN8XMoi96ijbRbs0nYckluQYtFwn4L7BnicB0lUDL
BQrDDLPvHIKwotSjVprTRseqagsTYQCPS/aaijxcdZ66ZRe/IRhHzk7i9cyEGrss
us2ZFb8JOGwvQDjovY25k3E3NXYyUbOSeb5MzhBwY2hReDLPNV6m9RbGWKSPAR2c
ByDO98VqQ1WNMUw2oEzBsS0q0E0j1Mr9oglXxKG4vU0ks/aXmDLFaxVq3+OuWjLE
mcRLgU+tVYr5qrqEs7K3aJ6Y3nwOyHo3+QI1AP64zeetDYeUTb44W2ypAMV9dklp
7yQGcTvpozs91CaRjd9twvvlMgsbSd4zBRLQ+iJnKFwK/8Yqvpnp+xK51LEvwpnO
holYFzyrQCUeFN25R+vk7C12svoLNSOgPNx5/FkzfkPJeIimDhPxDG4Ks40mb6Xm
QFVDqJzT1Ji82bOzU8EgvsacVsR8diVI1+KnCwoOgeCvK2UDTiqQyVxiIhuJMCqb
i2iz77OJFp6T/gqTYSQsNVXcbKBQlw17wOYy40SH3pNc41oc7HeGKTNn6VH7Qvd8
WZ3kMxINpK4r7Bv2bO4Q6Ka8q2txpJekOZhy7Ie/MtnREEGX1pWqatEa3r7TJF5j
MuFaRR39tZWu+SfsxgBydQPz0SmV2s0jDv/nTVy+V5md/KDgmT6Ikbqyl1EDZFw2
ciuNJsYfz/MVKS6N5cN/ISwPutgFFvmWRjRkObSv8X+Zg+gCnpkIrctor/EZ64gw
GGjoDQ8NNcBoqe5ttYX/WMqcn2WhVwusPdSb4CTWoZc1t8LsrIpmN7uvnKIqjBdO
CgWWRGYj8ZqKrYMRv56g2j6jVAh4ggg/Mix76FFNaJuCO/BmJp7oHlPJBB36UmTU
Dn9yPmi5YSjgTXT+/XZQR7WrCE12hbwzPMu5UxxoG/2Rg/V9kMXCBtwD8J3tiV6q
mL9Rnl7QLICpl0S3uO88Hvt/kwt3PvjqYwbxOAVS64ZRJa+SYn1Uulybrm4ZkbOC
fP6B6TVrzoaQ7vTQnywYWQBtMfTJaqKo/yo0H5YfJgSfQEIg443Q/RcHkFyGRUsj
RA823I/Z0TX4Wy3YHUcnE1fWRuqA/fXghkkW/KgjsFEF8suaQ4PrY5ISrzPitVN+
DF6z/NH319JT68UGAj4Q2E0xzn2jxEBVtdVLLEB2mHWqBnv6ZjB7oDjjInAEEWWM
kYHgyz2ty41h3URyP8J4s1MeQf97Z91D0cew/EYNiUwmLq0IiRl2aAwtUrpDGq3M
mHOWPQNbak84xxRHFcITerfEWx+CPxRVo9HdSGASW5PgPXy2p7GfA3Sa7wCO5w74
K886MHjC8rjg3hUm99DRL4UOsAOeAiSxdSy6XOvzi7Ngu3ikJWV/OneC7E2ftJaU
rlNr4mOmCz8g/soZuWZ+16p2FVpri+fTXZE0sHZvGEQqvJTaG87xi4Hg7dilX9hY
4IhSH8VvJQ4AaZBA29cfZ1Cw4UE7Yvzmbgh5jQGU/HWLc3FnS8dAi291OOdwLBaz
zi11Z16/mH3JP+77qok+Sre9DGhIno7cByVUBJ4Mw3FRFG48eSpbcPKffMhmmM89
XEdMCuvjrhIYWqMn7StvgVTmviwTL4PBy56COH1muYJ6l/sm6K9XxBQmo8vfBvMD
EAEF2G6+N6IRimFGmPXwbXYjU8pwzV6mMChIwrrlQVd0e2NYG5ml4zm7WKpndfKM
HM8Qy3sHf/b8cDdAtt7sfKm4zmI9OkU7i7quyMBQedJscGywdJQA5Mimscn6by1r
E6WyfHuP7GMylPpnC7FjtdGrax+dMDCkOSLeW4xsK0RGWOzoko27Chzn99M+A275
1RqPcoks7tOcFIRT2HopREQ/5P/CyDyYuLB+UueWj41jYNSyAxYeXicux7kg+7zS
vgnU0VJZCS0H+WjD7RF0kOpKQym2+ThLNU+ac0H30WaHYEuFktsY5oyGwns0TKuL
lQc/h+sHJ7Z73uSKAS0vsOveZK/V2U0o4SowyXLX7MozIjnn/zJ10IhsB1jkmAhG
I+oJM+IjWpyg64WK4X1BvpxdCVcYSlpLl7AHlKlF1hT10GHj8+zSLQoodwFOpmsF
eKsx52GnNuqruFbSH1cWPyqZmkYg7XGYXeZ3cUVXBaBA8UaL8mEI5vH7/GMtI2cE
VkB4DaE6jck51J8efEgnMuGoftT//udsKCEwv8vUqE0kieCl9M8HHGKzEeT6l2W4
9hwk5mvvSUIFEeT4gBDSlNGx9WMVXbxqLbZ4yVu1hT4e+SuZ+F9qc6Tui+UuS47P
2Z3fypHvfXXyfYzp+ptnb8J7I2Mg2PBqTRfr2pbXPYpjwmFrsl7M/w5n+H8Ae/XW
7DP33HP3YochQVGjjOKwd3oyMqp2JfLa4vWIzXHjqaKWoKVs4kKOY2ttMJ/4TTgg
JNEoeSokDZGJthYgp1cJXQF90Nw5kKX7a+l1JB241lx/1hp7A3kmdVd+cFnGOLoX
xgAJzyCwDLO7Rspm3Mf4FC3p+Uauh7l1oWKfJ0YWUdyx946iNelchUnMeBVB+Wxq
vSOicIxF51JvVjTQjyJM7OgyFCUgenMlyE7PrP/YfHUP8JXS53tnoPpHk3fwp9XS
1ip3NDppy+tiSkf5J+AwNqxPOE0KfePQmN1+56iYUDdIhE6KpySOInrECYGaPOBd
LlxjLgbwGZ2sFpqRhNFHzKB0pGfcpgyQ9pwuUX8mxczDMi0SW7gXQf9CgYj77U5l
QgHyJIj4cv3QYCqAqCLwZQOHUO96BvSjhjGsWC0RSvm0Ce21cXSBGCk/dObGTgUF
VGlnq7ZYSYTrRd6+NedCPl0DERd9rTU1/+WUmDHOfT86hvTFqvP5Pi8/u1i981P9
TxUOFSzZO50If5Rvf9CvShKI7WxSbtae/VxwZHlEXgxkIHE+pWTKCzvW4YCANrRt
G3B6Hb4fMP+HM5F7y44UFtcdVsqJ9QyzCnivzwatFzuWtwTzQ+PAgRTEU+21KSAi
ZYV3nbDxjmJK0mbdEmk2uDtw9LC0jSndqUOPkve55GMDn7HQ1UR8ea0IWQQznhoW
yMT1hrLMmtOlQf7LA1JG/FBjCQHx6ACvaJ1gYfan73lxHSjwhAEOdSDsiQCOkOMt
XFLzJb9BXois2vHe0bwqIwgnXh7+pGxBgVBmu5gw7RK6aIjZtLtTENGTeaWSRSWQ
dsu6ckLGTJMkLwZ9hSJSnTQnTNppIA3vaY8+1wZcHzkmad4nxONn5vhIkfKlHnxL
aAAIkDyldpl/HBlLmKJCXFeWu+7kstNL+0p9hHCT2UKv9Uc5mmyHaa/eT8b8mgwZ
WBJ+aYlSMpBOFkhxX8Qd12zaUX7i9mSdEwdjBd+zbDtXFYC4vjPgbl2LqJ+/K16C
vi3W2VjfBYa4aQeqgpvVFFyrt9HmXkQWGEHZwo/EGhCq0ZoEkDlhyUWSU+cy2N4p
TWeC4AkD7FIt8IKmHPwL2EoOGhUXmzixDGMXS8vPUnoar26qGDssVQY12xwkDsWy
FtPrWwNDxfyJB7hZTiT6YdrwD8w1mmTWOzmIV8RCCKCsk6iLvPcbd+325vGAekUg
TSk61VYGoyrf1Ey5lCfKvF0pmwHwW3pOu6+mN4K7G5JUVIiC1IU7nJP1tUaN0nix
NzCc1Cxc04/w7AJZHbeea6Mabx+KpMXsWgyfjHHu3q8Ibcfk1onysBwbqXLKhYT7
JdWXoIJA0WZDneDMZ+ILnXH8K9ZMcSL1+RGyexIONMqY9XSugFKacBNj9g/t8Kfo
oD7n+t+YPxS/64iFIwu0OL9gRpNUkXVavAHRjddg5YZgf+cCcdh+pl4n2CSb4tqk
GatS1SqnaFYp5gRfaqJb+o/b8hgRltErbN8zSBQ7kaZJSXg8BnkL6m7OWKS3EgMO
/VOUOp8XtBoQegcsNFFZrQBZKn5J6yN3mi7oSGQTwASWWoek+u31WnUSxAyClxSe
ZCBCwgGrwCQXhYzLjFcVEnWavJM6H8TcnVhzfLkJRyA1KpgCFbS6dXmgbKWiw1sH
vkcZwctegWe0qbPtww3FgzKvOcwCS74rZBIeJ8tXGbWCrVH4SE908wExuxnGVCjX
+PjG6z8zgxGgTKM9sNOzbCTc/AZMGogejFo3PHULMJqFUITIFGZVkocPxdRkXjVC
Nw+IITs2KsHh7eudt00yE6oeyDqJnB/oL7Z2yk8HXjFxT/dvcSg56uAoT8XbnBgU
LmLzbbV38WGq3zSNgnbQq+RkAG9UeXEaQCbGKgMGQaQqlOXA55h0vY6Icl/Skffw
2q7mALODpK1q8i3PPnQxFJHOUPD0l19LsM0ugtT7xtpkKAbznHDkuV88wKvoGSVh
mJB9cmeJSrl2l8CliRglyI4HRJy/MHy95IXtADY36jH5a7JVj+D7PuxZiAU+T2wN
NTwXsqVxjX63BUYrZiYUQ0+e5c6UeAKCJxsXLrFjG7dosA5ImjbmpiEYN03zVujb
IwQsVFHdPsC0MKmaslxSTYVdI+PU7dzF2bfpnrDOxJ6b5ixzPDyHXD4JAdsjB86n
zZJoFygzyOY5b+/3Cx26fUAF5FSfk1zeTV92FuavoMIKiaBdmVNimGOpTmxgI4L+
X8jyGC6/8x9HgZe1HBAAOCdMuU8pMK6Fp48pArEElBp1oAwKGT/Ew8jEDyiPI+/u
/Jk+KKcm1vfjEnXDE9kaN6dDsDVC7Ue7V7onRE7T5oJkbTUkBm2uIPnoHrF/QD/w
W2Xr+iXomVAPXszASv6i3loONS8H7a7INipnNcccJVzuKrfhqHdVMx18JDWyVrs1
DhKE6Q+bDUC9H4xJxSCMF7KpoY7ItMsTuPELHLhYzmSHPo5B+rafE5HrhsxRcO0j
jkZeCz22Rl6NHQS8FzjvkhrObVmRvtJB55yBMiHi0l+l54EZahbM9pO4naPt3MYb
0g6HZ7QYFcZjLkhTBkLGo//UVq6ke4aBW6UCo7xo//1h2J/UfpnIfPzoKpLXk4Aq
qGqaFd7TrhcVZESspkXOXEVgWX19mRiP/x+6MzhqX1qsfs4bHYPL5PK2uyX8JeJa
lZBAdmCj86d0CVPTHVaVgbYjou9IGNRT6o7qq2aEjv0Y2E6BEYhlK5eeDMFNyzJO
BQK4hF3orqu2EwdeXufL4KK2bTCXZKVMqjGWlUu29VmafIt+RI6wzxEDwl4a6gr3
SAdVMWgrlXK4z742QEdesmmLL+UjKnTQm+F+g7tShl/67iGxQh5QZ4O94gIL4g4q
OuQrjJADplm2ueElEhpEFg5DBsnhD+4HSkzIEicNfualFOb2AmTcj4x34tmxSqXU
QVQCNgzVK5L5nqsJU2yE8PnxLqqfDZoIz7nAi0h5cEjORmO+rvchAvgT6IJhj1ix
6JsoX+47LMMA5v+7YTAiCqBjHC2nV2L5J+M/NxTRo+sHpQxC15VWxCymgJ4+CV9C
PCARmowIQRf6nxJnQiUWKoRwbSSOZMkD1LB9BwIoNNFudXg4IJ6Vs6YlI4vnY9R6
zqPnX9bL6HKgnE1O6PpPjcMJOPbZ1TdTU+xsCmEAbgFo1KKrBfqHeQz4iCc1e9in
b6M1a2H+UYhPvs2jxCbz3eJ3KjmmuOC+dEyi1VxKmlL4YG7RO2Zq2TNpCS5rDd59
ujjwTA3D8n3DHC+/vDkFxFU1qxCgmeOtgQe0gcPH/OavB1thZ71PYwEh+EjOXzct
YIqyg2BU/NwBynHR6tPcCqhroBCcAd+zI2JlxhiIceco1aL4cql4lI2nTBUtR8HA
0SA80RSuazZwxAdym9OgmUjVWqD4Gfx5a6ZN4jbguTOzwiHy1yM7dmUCLQ7ssXHz
Tlk7zYeBHG+9ysBqfNFZcN8L5f2gZI7kMoUYZS0AL8RT4lf5iDeCNAv67GTnBI7w
TrMEy4K9pnyPJHBQV15Z9+php/pl4LgthxpCBGjxK04NfrJNJhzAFD6yaql6c6wy
gbrmi2GEY37JM2VJGFNC2H5q0SlKJ+7yEPFFICy0Q1wIWcMLTOtujwL+2ye5ZS1w
QAz8EG5RHHz85G0gR/bdVgUtQAuFC8b2OQuB8arrbTQW1ah7M22cT/t9ucxxrbFu
wYJ8x6SRIeez4MdQYwpdlYkayrhoFtjZKugQvxgcuYNeefce2MhqA2I2gVdtHvrt
fVnKGByPlvYV7Y9rIOWuXmqniP1EH2nMw0O3QjGnivV++0NzrXUbpofd7IGRBQyN
u0u3a03Z3B38KNie9dgiVhmFdUA46szJMvru2gR9b8/w3MoCufC0E2IGBj433P6U
PnNupboQmjuJgw5e1qQPJGkle5rUSuxCMXTyh/idQ8I2PiDkWtiM+TpkQKsu0xep
SOq+rSz9Cj8FkWnkb4Bzfv4EOAKH+S51H8Tusi5bk09dYy1M+wxzFEZmXUt2LsTX
ECNypLn54QmOf+YxhlTBkfQnapTIl73z7AI44HtpX6/IQntKqolR1UYT+LlArRc4
0skmo2ZoWZ8ce9noh3TKSqHHnNDrfHuEhrAz5RshdgtSJACy673zJnVKfYhQkYdb
VBxZ/u7PJfLv94Fn5a/e559wAN5zjcvwjtayaOO0fAD4dCdzpVH+iQB/l0LugzTk
NexCZ1N7hkjwKe43qnWrYpT7vDkO1j5VCNIZS89ayD7ohIFNRHc9yCKIuAv+J9aZ
7heySq50gFG0K7zDBmgmdHBmJfKKco2OLsET2ZUHDOYH/IOfcB2diMOLNePp/f87
PUyHiUSN68qP4uEQBhANrWgqe1WKuPpkI46D8K7XrGdqfl4JbjL7mCu6ozy+MVQD
DkKOgCq83Mp7Sbk2v64eSajmqlcK+hM6KuiQ0ic8ENwS5MsIjcFzfHND2m+OFeaK
4FynAFSnsgycT1Ac+B7hNG5KT3D12Xewk8wqy7cOvKzzw0uSNXj3j78LPhC5yu3v
ClCNOVxO8Nfpv2ELXI+vY52cOmwcJEMTCelKbMibS09s72M+Jj+3bA5mKf2jx+9n
GNQboz/hdDzSJBxTGmnS/zoqGt4yIbbBqU5s8Z7ufhkpONN+nQvCTwz487e4vbvO
Nzn6U8/ULFEIBxcLufxzznLwdQAbn8j6IqTKohPLVIW8q8P5xzbx+M4CiVsj+TYZ
18wN2t8Tfc9Ghi8+pycBqRXLoibSRuIbEHZxdXkS2IwGGUINEzIs5M+Xp8lHCLUS
j5+9hMEth5XpLk35BGlIL4wZAIgEK3UjUqOgt0R/Yf190e0sxc8dVORTMwBkM1oO
Bsr6qqd8fLIdGFgZ/DaKFsrrx6pZRZ3FBdJMMYzl5rDZNXdFYS6aLIiZ2KETlcqY
L1d+0SXKeWfskN1rKMJX8XF28jnpzHb9uEfcySvAZ1XA7yIsVFgsVuCzxc+0TAAI
0NALiKNi3yv5MclmGxthMfhBN8684MGzX7+SrMceCQVrfPYRR6DwHNTayPCcanXA
WzFOaIVNw66TE5RcnGKMn8ROmpWVDQc5JnY9qbh6Zv8OEnwpt79QcQ+6GpnkOY/C
qzYnHj0MgZTZaVZd6iePd10nsaELRG15/Fqk+svTGk1Z2m1h+Ja/aBbhhENvjwQg
8l9HAcUo0rb49E06n87hTsXA/iooXTnHDHmbLfp98SjNrpd2tpv2XMjvEYdDz/fo
WQtd6xsRf/dNuk/5enZjnl+eNLkmeqQSNz2gkKtraHfzOoX6VQBHbwSz1lFfts5k
H+2qtrpfbaeJ6oETI6+K3hk/WonQz4Y6PSiFEVPmbTCvWYw9Q3GiRCuxLlyR2kWi
SLL9EqMmmLFppu+TRG+Wgb9HBWbAiPYD2hKRPlgPZjxOK9q/sT4YXedJYANTHe/+
5Z7gnzezNjppQPQEkQFPHxEI08RX3yLLJ3LKJw8XAiPUCs6a/avPk9TyfPDt87nF
VlydoxVIHcV/yMMqKNZjFDOlvx2N5tP6TLwXc/Y4LzcLnAWCTo6wpZLOGq4U1Jp/
//2qY9G8YOfigASnPugtndLoYGKYE2agDVVmy1NgTlasPv/HmFWeQPgO/iVOlISe
hwDOe1j0Wc8S3ZGfLHn12DiUcm5r/FVcDqdnVtqWuTgkbTDQikenfNUn82Me6o0Y
ybuvyMaXa9HLNUwwo/e9eCMoayXpnJNkQjdJgSUNvTRWXKq4XXU8itAZrTZuXugl
WbKfZcfEF/PQ1aCN9btQF96XWIHnWytOczwZ0rwKVpj9GP5J2ywtRnEKG82e64ri
ERQyg4kf5InpFoDsBv7ZwP1quGE0tIIkJJceCfkrpANeUS3i4Estyd0eLxiN+lFs
Elcp2hnFHB85d2znmpe+dMBkap+HD0t4ZthKr4T9YnVF6VmdkFR71G/21iJUvf9K
dVrF6HAyhUe7n9lh9cwYHJ7ByfUMoskEagW+Lx0lAnLup/0Sz4ze3jGGw4Ia72u6
zOscMawaEeH1tF6StDOiwyR0gaOu9PD6nkUT56gLHFOfffw8ZyFFQ/QMxoE9PK2b
Bjqn2XFckJNtpvLBAflyoloLrMwhL+8+bq569INZhQkqDxOwVtUdd05iM1uxgJKc
cDAdC1AHPhUw+SHSyVcxVUHr4jwljv5vvuCU/Iv1s6Y22Gw2wcdBr0bWQaFCnTkF
Oo2WpLwQjTFsGwBO8bAWOhqemE0671yzhv5s4/Sv+6aKvMJ9rgRwybg1VCU4rfpW
u1sFTx9KIvLwoUm9yQ8eL/A53h7bF7f0qvHHOp84zpV/Hm8NBoY3yOHKU0ZmrlCX
CkLFrwGGewvMrd/r6U7HgIj3Vtn/X56p6fcv0hTKvV+62XRWzvNXiri/CUmVnqnG
jSpTXv05OIiLQjkzEMAUqmE4XckfOypXa0cpETdrCgiloX4yzCDBrk3JKTvYU+9y
aqOOcKKUuvVoHzuLvtn9/Eh/IP9LUmDEpppDglivwaWAlYYOTeD367VgxgLpJAQL
oGkMFxtCCByM5BFRON5lDJiaCM5sy4GtCrHP5M3yeEblGB7uEUGaqqTIUWglLmAL
LU1oAbiVVoCjqMdxXubGWmNtylG5da6N9jFVpjWvkqNHTr7oT2whf6j5F+YDTUR/
8myJl7Xekav9zXxdhYrRZuO529seKfZ2pyh63+ycfpNWIbTr49+adJmykfI4KQs1
heMN+N+gJ5/Rfu2lwnTdusHdHNB8Dz1yiP3dPpfQ58F/Lg3Y3wSlNj511R9jOtbM
axfiD1JXxmgLZgAZ5zYLY0j693dJdMXRpd+V6ucUs6/KLrd2n/tse9NxGROokz0b
CXnkfHb7941HoC5CMT+PFqYhlR2bX3nwdtHI5OlPBfQ3mPZbWzakc4fgEUkrm8X9
gP3FC/6utQImACpGmJ5r+p1N/2pAkvgkI2KTRYDy+IH+slDfJPivNXuBfPneLvh7
E5LZ4C0RjzQBDlyPDc03u5edEdZcOKwQ3p3qBkzE3gNZarGiM7C1pn3FCQGBceh1
QtK/GIEBaBBOMSGg/ayKIAXwi4nyqIdGoTcq5AnyWRocVRTyfXGPS5Sbw2wjR1Zt
ms4FsYfuZbhyx2vnYUoYvHI+uSKKc5sqPy+ntr13TfNhrdeIyhbxZkzNvY8guVig
ja7FtlOBrDU4eL5MZ+lgt2EFDN5rvKBb2HK8E+g34FYa+uGbWjxxnPpWLxhjG5H2
D69Zm2N3yhbU+Zp/nBFDbEgrBd3H9aCdNpwpWGBQmUfKgqqdVmZXKfSI/52Us4sL
YSZnTHlR4PQtahVuxQMXnzyNM8QsRXwq4/+r/oONTuTyCYyJ4xvcYIw8jRSy3ml7
LWvfzXjf13NLIBjgI1e1y5BRCIQDtCmBVtguto4z1LdvjMSYIJQZqetj5wfandfS
3tFgNfBg+6DJILquN29PZ4SbgF7q0B1vVk6KeYwL7KcT5EVc/+r4snSYTqr82qTG
IRCg7l5/ihKIiXFO0bpgLJDdAMyFpT5u57wj+HqR8q4RHqezgcy7NfqFSw3f3ZnD
mKp/rQZsrPnE3zHo2Khg0wtvfxScwuKP5Yvp/jB/16Ggr86JcHCD/3DNsgRU72ZX
/arDFPJhplq9vi1G9jVXTbqM6NMKTdtcRAeEBqwI2PA+tAGFy5mGMKo3LdBhT30l
Gy4EYoRtCk72COSM2ZmVu14yXOZmTJeTG0u+CtIt5zmFKZ0H7LFCAhdt7pusFwEa
lUiclIFzhJ/Q2jqBiJI0uWVI9bkgd44bLc5DNULyHEpkldf652VFj8Yd+LtHIA+R
YOE6B7xLqeq7Gp+X383yYwDCjCn8fbeMWlxN4n/zinoYMy6H5j3E3jHZ92ZpXBfO
yaXI8ADkuaIEj4X1oZDJHNa4dQIeC3+cELezlctT2omrXZ5i//ThBKxg8hcvQ8yo
ts3/OmyYEz5cstH2k342m3MGHe5ObtjUEV1mlHAodVMYGSJb0aav8vSz/d7eysDe
cMfzRWAFhwsvGe6wn0zvO1xWeGKGwX1WrcPaP55SVQ4pqHHKN0cD5F96bQp2N9pZ
/jQ/e6C9o4NQoDUL5bPsCmY4hw1GGWFp0pXz8skW6RvcT+NLA9Ocveqpaj72Oe7W
eQJn2WFN5a/2+5KdVfvrMqGgpd6Nim7oCQdsiyf0jMqsIzE4vs08H4Fvyn/mfJwX
f6GC+f92Cx1KFUv9BAlSnQ0LxRgVOiiZ0vyOq4xVQar9xPYNh0mpdA1UT2gqdX2x
HUK5FzEp0L8RdUFsgWgSZkYM1StZEQ9m4uRgRmO8e4+BnlH0c5lgGC8DvHl/IItw
X7i2M3EvHHR2AwW7A2TD4aL9g0g6loipH1ySa9G2PVf4pMUEoQBWAdT9nz6mext8
NOv4wBNZymP8cSQc9xzVjLQyqoLWBBMGxvdEP2InNGCFKzZtDukXoiJe4VZXzryE
B4/F7X4pdzF2PPuQO96RzUgP9ur29CDcNvdIU/cjWiE3sa8zik63DIeMc4hUQl++
fi52vrrbnIVHOnGgtN1XNtROFEeiskFKCkMn8Prd3nmjZZ3bNeyaM2uacItgWy1b
sgSO9Kt6KKGVapYZE1Rm5nF36AYUy9YE1p3KBMTRZCbbVG+8l3R6ZVNX7fCsieK2
NK/tQENrckPSeU1+/KmTcZ7A6XDz1bh9xsp0UiYayWUOT6CAknGZX//7t2FuLhbQ
eTq5BYlg43CbRD9hI2udGOy6fjqrXATewwP7QXnycBLFJpfttoE75GBNUCcRuD9w
M+nRtFS0e2kphnTgbtakSG0PfMdD2cSp4CgwaBlRL+mBsv3iUrvqi+NT37ZoY7qL
VWoASNWTP8FvBs3SY2/ynKVJFOpSd9HEshdDEZXAPxLN+RCeIb4MdDOUAC25LZ/r
0uyhj0MCLdljlDQDD7PMaj4YaBehTdHh8df+RR9wLj8W5kAnITECL+h9Kq2Tr4c7
e6XxlxTaJTNl6sSXBk24WokBofk/Dxkx8kqXJaGYR1WGlJiCZqxM+9oYBDLrQ3pQ
hiW1ZULTvE+fA4H/v/5IQeYX579yWmjhIwdtC85yqp/zZJl25SFzFGPAgBpt2YmC
2nzelnuMJdukvTR0IVMz+w2TelR1iMpOWKFISM9waLtcQ6M+eBvL4x3JfnmGdcT4
X2vD6wnoOYf8sajMMDHFOQtAD19oHdcDGbzw/CsDRKa7LXV3TE6uAJwZntuJa/pa
e8H6c8vzFUmERie//YaL2j26p47H2u9mQ/3lN9r+KoWu01ZVdbnTqHZ3sB28z/4x
EZm4cA1+WfC9waZCxrciCQu+5hEzyYzgf4GPJe2OqA7y2kQxrjTcTClNgfGv4PU0
VSbFKAC8AIaglElueYrishvZ3LbS4CqHYUM/kdg9DHKyKVo/+/nd2MgAkcJ7g9FZ
a/HBSWTZlFvEyFHMdDm3N84BFRioB8EWCF9ch2Nfoq4o5QIVj/m4pcAVWnrM1QbX
NWQtyLPKAEqOhzhijimyswOpC25bvR6wcDXT4u7s8dcUdPVXPIVw8Y+r/ZEH4PPX
YVeOMzAYaCN+AslI9sL7ikMQvIOv48TOlcWVVBXbzz2YmQZEn95fTYEc2zPmhJHR
JoWhxmKvtaHwO2+3QRSEcRgak8MUKdikqwDLq1gBWuhKBTAIJZwTFcKPpr/AJoQ4
C6lXoV0F5HQOxh4gFuc2Qq2eX2gM7ThuMUWuD0apJ2MemSTOyNMWCvLFYMOmc9k6
jwt9o/NbWt+U0RzPjk9AlbTBKrF5jvJUv5RY4jJY0aryBzgHtv4Gy1PBP/KUTPEH
FPoySLKfV51jlZF039ZFxVpClNSpFFG4IJZU4+ApFRY2NVMF5V7VnweftFnRLrS0
iRTgeioByPEW/2v0Z2lZkN9NuCSbRZIOxYpxl3ewU7KFswvnQctu9ISMZT2u9gVc
fCzrjL6eC5fxRyjLuDwqR/PO/BqQL4/JtoKUt7JSJNuDbyBnvZBENFYjCwZtvAb2
xfvVI/mJ6uToS/EMJb+An3IwnnxcMU17Gx8zzrIcL0f9kDn3JftZvAVkJdiFXRni
8p8F0F2HoOKj694yoPOO6uQdA9aLeHBFW/xbza3I6lZrtAatYQ70khhbk6sv5MdQ
WijT897AMOKWeZhGiMGJ448jnTqP0EwNIrsEoUSsM85tFLZK+zOpl9nwkvFmB5QK
AcziWHynsm0znWoZmHpMC7V8Tz4FAfJGyOJzZ5cR9be+NshhYCtC4usWJQoK1lAW
kw/An6uwN+hkPHqPVbJP/JnDm1gA8bpHnqB7HFO5+xPfvB+Th2KIzbM4QRFeYmbU
TQELxb62hV//90SRQzlRgfgIdLU16RPlKjZ31dpHgZ7dJymF8e96ktiWcFBTnLZ3
9bU1tS//xYPyz46wdndvOMxsx3IBco+Ni49JR5GHdo8v+9V9gSRqco3nQvGpWhcN
5hq5YnvLIadIg1fQgFXSSp1jNjDZMJfG3YXMfrmdUdJSqiTawq9BZz8TECR8jXgA
FX332GkfO1NnETeC5IoFf8uPEhFa+sbLovk8MpJph5fLSPGw7jpRsj6LdYFfZcCB
mng/8ijsixJgOlHvToXuTda6ip1j0hRFPFngyOFup3HSb6s7P2GnooSxzZDXzaR5
cIGEJNRIJ9tQVJgEQUUXW6hOjjRZRJNbaf9Tf2mbiZWFWhRJsCZge4Z4+Sg5YSN8
XdUsOoMfkEFUDSpuD3LORhi1AaaiIuGeUnT4mgqi+JwalrpLT2O1Wfx/mEa5QmUJ
PNYYIha09jPKkx2cU5K5iZvcVEB8MOmay1+Xk4/R3NeBAkqtvhilvOpV7BPvhCKp
1MOEzBOB3Gew/aqscC8xsaFqyHHzPIxOIh2sZeHlndWfZP5Xa7hjGZiHZk4WM1ds
BkBmxc52dWT8U8FR0cyugb3zfbSu8vD3xNiuBa4mKwcMSbk0ZiBBFcHe4Ouc86UB
j1fS4vv4mKORxJhh/8r00SDOh0Yf06hfx8VL15igXSa3YOVYaAYcQc4Coos0Adzj
cj/eRE6LSHPFlOMWrG/ydyI22joYQFGNCHSDgATbFfHoaGPKG5JFt+nr+Og3gvOa
HClKXknq+mDKSIKt/l/eQuQOB6bO8fQ/4NseAb8745cyYCuiWxT+sscbRDO/KCMo
X0zvEx9/uoIPaKcjpq0nwFRUd959na/ATeORktkM4ttqLPLoDuzmc8ZehZsuV6gC
rjilnbvHF6yuXnZgsUPegtbBRFAVnArFP2gPB0PD9b/22M1/iBrcPo48EJwFuVcV
Uu1EFSy6W5wWotDX399iXs79gmnAEOxDC4w60//Vz3hh1mi/d1GAaz3HBdX4w8Jp
7UwH47cEMSVhkjx2Z2VsUjBIMSRAvITCpgoQUkTb2Yc6gv1eQy7JM8oUXSbNTa9i
bfzenGccg+A0aFSwwpStjtYHTUwMwndN3Ee8RzIf22S9nHYKw/pdl/MYJDUBPzeH
bHhsi7N+joTL3hn8GqLeUrI3qo9Kl/nxbhy1+/k/Tx1eiD4O21OaX6jkmi8zWmkc
IxcaSa5OrgjCPu0qcBmxsRnTTumAWONtv35AINFTMkV6L2IOal5IbyPMiFsHPFcM
6vNrcjwtk6Zi2hT+cFW7jdJdzepdXELhRRHxKWQt29RuWU7uYPcym9mSmcpM2V4s
rUUPZvVi2QPyH9jXuqzyxlqBN7t2obsavUQXGtbsyfktzpKcmV2XUP9vL88q8ezE
vGNTKYvTDU3n3GkOzY1pE39P/j7BXG9KY9rvD4twFpCP+kiTJCBrtNzT2Tr0i6WF
qlaUHC6nemjPkGLQa128LaQu3O9iEjZLE6C+WqzdPN0enZTZRAeExYYca5/bwBw+
mngzjtJwf/Q6VtYK7XZCpoN/+1sPnd0V9s7Xvf6bibf2Tuy3lKgixAiC8jb/2JT+
nbT080wppLVvD4a3C3T2qe2scmqAv/vbji9D09oR+5rH/rzt5c2x5rZFuAsJusDe
Zbh49df60VMRPRRQuYjPMMgbVMIy7jYeFK0YxBcqMCyCMdW9B1M8ibc5olPJgKzo
nSNldmDHYcGYK5ElA18anlxguww98KaeAUVebfDP/o3LRcFs8DLoyK/7hwv1YblB
av7hzimLAABfoK6h6qNS3LE9iNLJNlsMjZKHb5YzLLahCGrVnw/UzjNsIEuNoPmt
iXEOgnBQ1gAQuBhZmCVxwu1q8vgLX73tK75vAWNIC1oqMps7oQ7Tz+FgE03xK39G
ZSpZ+lgvqw4X2Oz7GIm+/99IO75vnp87weRlhpFIl8laQ/n7MMEwuTWE8LDCuu7i
QfTDffBdSeQvKpcYRadR2m6G5LJY5G9ZciqbLnDgqNlwr7xiGTs9cmj/b88aIWXa
lqz3s0ecpRDILwUrh5ON4VqEVkB0h7TjEHXgANCwCUFII6+7LWh/5F44Jd+MPyTb
e3+sQKB3YQh7If1c/xOmo1r/StCuK3FZ3wlGHlhirSt/EJWM7YFI8K1zEqRj/wev
TSKll9X6VVb130iDMYM4UkrmA4B32rOUsk9y8ZRMnDT4CPRFk+BGizeoKAJsL1yf
FROrSHVU+IubBEQmjZVdgx1aKQuxFupbCj7AgchemwiHVvxijLIt72Ade7GpV7jR
PFfmaGTdwKliYo8zcxx3fvb4YoUctutmJR2zIzXHz4OyKUuMq9+R99jxl3jzI6AO
8YfaDGrPWdJLADbChpqGVVVL7ZrnZLbzCM4GUOS25P9eDzaZ6rrPbmYwx/T7Vjjp
Gh0+nY4/4N+yEU0rI9Hmr8x2nS1t1TfOhD/gCWTPzx7zcohgXsBbCHOXD0r5FtaA
IYhKQxtmWJNTyRbMatWhbB5UDsSAO1XSn1RdhfOvKfPpllTQJ62ck3hK7xqDVdTe
1UJJnjDMQmE1d3AMCDwERGiN0j5YGsib7pWVDKEJATt1UgST3fxTh2nj1InF+fWT
5vtTF2XLxL7sSj8krpCuKoxFGvPsErEOJE/J9KWNdBV012E84v6selMMKBRzhCNW
+XH1opvGkD+dkfPaSLug1fcNEax2sMmgbKqqfVEYP7X7qbqhRlO408ZE7CCMXakC
1zhNg5L0vrPN22a+89ANyfzcbBG/R/PuUVn1WH31+Jk/Ca/7gYfT6HWZL7kATfBn
lPi00/liwWHHu2QkH+L9sgzw9NdKGtf7payL2GnV7SdPlI5FczpFfVhMFbg4n1Jl
wBLWFZOSjuHpetbhFC9YJaHy7BzYT40sn0y+8JJSQ60ve5HjTKPlxICVaSqxKI4c
uvM/1hvvJFk8cfgNgphm9MsqY6T1cvI8J5NEibMJfKB2w8ey2/R3VBOezicAZOv/
QhzRqx1opuUhMiZGl/6C97ZYweJOr+80VVF7z7uIq+BMc76A9Vr/SBIyvFPPt2cX
3MbUVv2F6u5pw0QgTKlv3tN27/wXJWgnG9EPJEgMKkUKgvGZEFfgvBMq6o7q2ZH8
sHEj3IoiLwdgGwOc4IVr5iiKS+31oqAC6ed+ednezX4ME1JpJu57GhRdBI9sE5bo
3uX0JxbNtVPK/sFQtnMUJu6OTKjlpdXtZupkVg6BL8j4/T+I9eIzZo7JizRBxaPf
CEFwZk5MFCLQK5SwtjXxKz+x7JIlZCIYN/A1iD4Ea3jbnpRlIy+JncgvUPVqVkun
qMku6AwIYugwrQ07y689KvtfoAatw7f6wjM5Ofh+hoX2GhbKAujIU1/AyRqkX3Z6
mI2NukegqX4Cxfmlj0Ws2ORe1hq8iAxM9FcpVs4hR0vw0jq9SUorU6wPOhq11RhM
DvRbycm2k+HU4RpK+3hTy96TSscvFJZG2J7HKlI53V0cR4+ScYVquedEe7bNOg/v
LushjVlbW8KRTOu4cSKmPD8SfzphMHoBDsc1J9mDbgkvrf/TXKiMX3oH6uqTRLLW
MskG5SL6B95shiBHlcJ83HV+OViQAECI3RE31xFENibn/TPMJTttCQJwJ6puqT61
27wieIjo4jsWk+03P39FP91D2Lbjrg/QbyWSl7kdT3nI6LdVsM3l3E8jTjy5zjuY
Mvp0fA6znZ2F/26RfplZI3lB+M2128qipXnFqjvOFxiU0Qax4LOwxhB/oNV0mlVm
pSVM6ni42/QqzzBSV6rNIbgvy7fvY38GJv8Skw5gU8s9XqUgKuNOr7ZVqzb89emb
2w51itbwuz8CUvjGXVwDiaOU8NUOnoEoRtTF1EfGTjJBxpXfuk+HEkt56zhmHHcE
6wd5/s2WH6LPwGiBOrg5KYpeNGgr/nrGw67MmU7F6Jd9VKOtPkZK+LOiNqZBZJj4
wLoMXUEpHpzt/iXZGdW1Ya7omfBA25GdXfUqHEgZnjOiBR/7UpPj4fhCM5qPZqNV
1/loFF2jpTTEB0US9bjjQFOkccUAAKycmmyU5QIT2ydHcGuYzyg5x9Ae5SE3QtGi
JL2gCOUg5eyOaD6NGYOAw3IJdM2q4UfW4c3BmSB08YHCE3FGpNI/n97beqzi5ZKC
08ERHrbGkYVgOtLdSzjmjd7j2wRw909hnHgNyAii+NqlLAbZo64TxD0RDtf6Nu/C
VyiQgSWcZPwYchfsA4f/tAVG9MP7gfjt/+OSkBRwSXSnh6z3kl1dXOjic3N+ofT/
RpWwfBZ1PQJtB/OhOvXFntQY5Os2OrH6wAJA4AP/FYSXs/VB/9UAPOHUWlRg4apt
HazAuxbqIGnYPO1uOWAzU0bihaksW8O6MxT+XnUUuuzFnyq6GVznOo7zbHSBt7sb
iI0V+Zov3f77TvW8l0+NUpUQonWvMAo1JZRqLdSrEH5w4j4e4MiefbShipZqdi6a
76BXshHYWF2hZZzVctrEacwWX5R2ANTQ1QiHHwtrqhaCgOPlKtv9rq2OgHJv3z4O
FoLc8tMQSnhzch3BDyM5FaD4yTRCZLxqaz/FM92kh3Un8Wnu8UkARC6Ac+L+Z6FQ
e4BVVg9kdudklCZfWPOsC9Yr60WoD1V6KfGQVwSk2LC50FF54BL3lXepyRpQVQYO
yge0OhA9OyXcuCy3wARb1/hEXc2KBvzBt+eePzD48jZvGzi0DzfyduGG0LYkX9I3
VroOQkoSl4EWBRbEs0xUOgvPJR6HE5nd66zWtj4nGu76z3Ag6gbE+XuD5Zye9Ot3
Ne8Plh76Cv9lMDKpS7ipeAg19SbMCdU2qdw5JRbPHLoN8gaONxLnXs7WnVuJcDVw
lT0cQkW/wfuXyxc40YfRXBNpN2oUIeaLRmbDpQk8vRF4XU+K245SUsbnvZefXKQx
BcbLblE+ZrY0y/yqqYbEM6IwctCA1C9hVwSVpgrhDJSBAhDHD5u0LRGWRoEH0SYA
+UZwJm2gxErK1Q7xZQC2htTe2laEqIiumW6EtPYbIDlpwA6iKPAHAPUIL2ATmnMy
zAKsDMxvlRLfe2pd8D6IbU6nPsitsXwCSY+RWawnt7iejAShwcd85UG6U/udUaFp
pXkU56QFJIYg1yECiErantUA0sM5UhOWlbtv2jvSeWeoERrEyGXYCF4cQ0yYUPXC
fxtLcXqB8xxEn4gnC38d2NXAHfyF4JB81A5ayxeo+9xBNMXgBwsmyvsu/zNcO4V/
AJAuCnhNS9hJkOvo8reSaxG906TPxdk0JiP8ZMuTKuPUYWPX47cLPvHavfxR99+Y
61COOQZ+SenYcQOFSo8QNY/ZbAvAPNESOb9eHyD5kjUdPdhjWFkd9WwiiZwXA+By
cFYjh+JSvLEJ4prI1FFDKUUv9LcEylqbJU0t27pHk048Tunbvlk9NfuDR6Jf0/nn
`protect end_protected