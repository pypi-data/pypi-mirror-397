`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
bo49trehcslJg4im271Q373PMZb6Hfd6I6ioUvGoQ/S975iI7i2fkjr08qeqKXcy
Lw+ttOjek9IbOjcTSYn4p72ZrwrXRPKl/p6J+QKxCrIwTf2+6CxhZVWEYlPYEGgP
HFVW8XYgz7zFBMFcbZJOxtvCb0eltmNrAecK8cp5D0H9ju2VvHUUXEDPGYJ2jB0R
KvcBIcaQqyaVGL2dk65I16J5U/VVLaytXoLAMp3lBFZeQN0cqCt8sD3NTYRyy1DE
+PHtaJGVn8H9BjjXZ4eTl0zyzspuooa1KIbMWPcvYBRn2VYFUnsU351KtXMaLD8i
7YO+kU+Kf/5D25q42+tp723R5fgE4swQ9PIheLiv8Ao0LIqrf2y2G0Tj9mKmCuB1
m2p6z43dm2CyVM4tNOK7rCTF+g5P2LPjRudd835/9auE/qIw+Gh6xFbMkgOs3m0X
/sva/LRh4hHSdst1uDhP6m/DEtmPZLyJtLXP2R0naWMuFjzp+OYcS0O+SSjlhgcr
i/Hkc22ECduwImHP50V3qkVXUMLzuPRHCZucOecX933j1KpPLAq4R2rguPoPhlKf
zcm+ywOFI9zc0/M9r/Cz1eF5XcBt4x9Dib8QcqRvynGTnQ03OqRzMwIiOpC/Kcj/
WpTxOBFfQMjd4oUlHU/93/B9/9PJDrdFxlPscQRV5Kzyh4P9pITl9vicsYi/u4de
ypVWfLcXEIdf/WYt6p+ggUG2++/CKHLYB+AQxFln5d8kTC4uEVtOxPlCNSKNtV/2
5f8Gov3BoZdO+90S7hyqPLrGD9CchWX5g4gm3ZcaU0dmJmyI5KTlmNHc30gzwhZ5
qClYC1N4YYfk4xbaYHG+uHrOvlNzDa0JzysHWcTZDqvPvUeW4edkDdhABCVNPinz
AQ4ojtWUDCy8TvHxvXcV5GIFRY2y4yjA2dAv2rQZ7tSFRPPUQAHfnq5gSxEW7Mpg
y0nx158Pv4uPxxm1RAjcGEWo/WKM7GvzyUIESs0fYLyZmXvlbbhbIjqg1BLnveaL
Di+MWHPlITF4vU4Q8J015as3x5RYmGMEdnZv5SklJmjusPF6rQYuURLMrB0qKFPH
OAzOnAuEaZV8TJwXWQ9uMuUsI4hKVBtSpJA2l90uH8luO3yPClDqm5aOGf5z4s29
VlKCRi+pOctAVhZ9VQRTHt17VLQ8bZRJDPg0+YpyhX2s9nLWAFf5QX5yqoD1yAZZ
iuRLqGm7tfBBApAlwoL4OPktAe/u77rGcukl6KfY2gtBrgrGeXKPUy7CZMcDLQdq
wbFHJeXJu96cW+EHzyXn1AucbRkwDEYfBSwkfpsbu1JsGFiPWm47JSDDQFHauREi
VVqWhh6BEfyvlem/kVz/plkDtEjgMNI5KurMdjSaAj8kH5uPb46Ru87dLnIuAGIS
v/1X9jVWEYi5J0sYlIbGbQsRZ+uZHzRs85M1FLRlI492TN7S8QxLkAEb92FKFpsW
MaU7Hz2t+MW2B0qsIuXBvxFsfa6ebOPIwIDhzGMS20j877/7kiU5cAAymzIja2cj
fZsd3Dj4znsXmuthpqumOB7he4G1JcHoUtK54kT3z/igwLYs/EgMroxLAC2sDzzn
Boeq3GfXoXu/l32QS4CA+sQQrCniqiGVbJ42eu5WIiVMSuYv2sdz5MlzrtWu88b2
Utu3Fn2ti8U9wryitv4dkdClWeNCXH4w+Y9OtqjqXe2v2+tDnAIy6lECfr5dSPrr
bv6LnDRkL+AboBynSWlUC2Bt6ILbzKqizOf37OtkBB2Z31C2viRp31i7vucHafxD
LkAbfVNhZMLfBWNlm/UTNCcpqu9gGPLZMF0C1YhEDJt23G95Y3b5GlUi6NsUAEfO
9C4XQhfUcGwD8GYDhQVU7Ek+aciwUJgv1OkazOADTr5nP9rdkYzxQ5b2i19OVUYm
Z8wMl84jxs4hW2420FyRnGHHdDu3rTk3LBqPW5qLSP1IGqBkx7dXPQI1X4hWuQtT
RRpjY/8sGqUuWd85hEGbhwoqwtokqgjgEwcprwgijPV9aNR/WP/vLrKtFsAf4KtU
9t9YWNeAroI6sYNca/gOZMHoWuTfzk43uHcL9ug/6HZ0s5ONDjOVwcRJdwUtKnL0
or+jhTTEU7y76LTubWbtujscHNMnUXuqmZBamDpRPXnioaTbXBLgH6naAQVS+U+G
etJVQWe5O7/wyCFR5XgO2YkN2prACfs3ePCQNkGl3RF7oLpT+5gxudVURojKlr3p
HQKhEWx17tsywly8bvSi/7plGGsm0ac9Z1cktY6ejT5x14hdjZ/959WgnGvNf+IS
k8eYi5hxpbZ/76iApP16JMazZRyS7IalYojDMx3pPcD6JHAwQ2x1AtGiqK64L2O0
rfpDt/EWmhgzgrxXcMJVN0mH9wVp0OaXGyFA4cXBy/KGN+Cg8PZ2l2HEWO7Y5e26
+yLJB2ntrC/MDqy9Fzf0qO5INbV1fPH4N5s9P9pm3GzyOiTuDN0KUePMrEx4BZlg
v7AFRrR4vT6sWKHhdBAXWXyx4IHURxptJNhSEIwBo6dihU48HnpQlzw/Rm5HQG1B
J/F8LX18/Rg6OXIzG+hKuVDVNhxA+JCsRG1n+AT5lNwZjHkBYNTPX8hk4j2qdQim
C+O3rhXhJrzeDO/w22xCt8lnlBnCD/v17Np5DU0l4Oh/+Sy2/lfegYXZpDtD0Wna
6hUWUp73xn/0I9Z60hmkYtsF1zCSPUNjRUAyEZHUZ3r9hJy7aUIj6sok7BgiLqF8
GAFOcyHt4/xdd3vxFKgfwdbS0PmO5QHVPgE1PyrwGOPBZkms8JrFI6OYkRWbIkHe
+zaMXfTTMnBt9aoogf7xDItEvhw9Lf9lHVbICkqI3V873NY4cVAUy1UGi9MLllpF
iIRxTStCInRCE6IrT6bKHhggtMqB1PdFXqG55bPV2hDY/OdN3+o7AOxY4C6pxahL
7jJCNXqP3CRuYW8SCE8joSXaaDmIxLkwaqfhzKShxk8gxRozRORbwcI3N2+dMAra
Nlc9mDub+nOq6XKRNW4kLPIx4vBDDao1RiUsQNx9V1p71w0Wq2j6lKHX5XpLdUbd
vv0gxxgxt2b4WxKAhDUKn4o36gjBjKs38833TRFsEPZQNvhAtFiEvEPwCgDkpeNF
dxIl/UNh3PvTzQH7BD7+T85EG0K/SEzJR6izLXfeM7C8Ql5KAnNhXnGyeINZskwo
19lzJF3ukO8mzkhtz3gI0m/UqEWYFuUHnymfdjxlZf+f7fssDc8ummTWRJM2pq+G
t5uDVxKXNVUanE5UPmj0Ngzwcw2MQZIW+G3QXmnptZbrqtr11+rPW4i6Iy2b6jeE
4Mhq2Kd+zN87MUpEREiVIzQ9UHyPm9+xtDqtmUKGDbdsTza0vrx7/tQCp5aHhPU4
5VXqqf4lDoLkg8avHfC6fyXN9FKndAxWBHhXZcz0Kl4In8Hdyif3GL7N+NvTcvb9
mcmsyf1kYOKspvECWMp5Zl8P8vVKN0SwUwGnMhOKXt4P/ir8JnmG9IuCGTQNqO/8
vpp4K2cpr8Eze/sjvITWj/8KLMYvn2OCsFc6ESDsLXIRFsN4WQZwoeVtdfiCyDEt
cFy4DRe/7f3OfdRxh+u/rwnTNcLwFYPuEmqViCukDodfYv2Nw2TcPK1Ck+pDvnsR
hV6i3v/AnD2fknN7MNwF/uommn/4XjdrDuejpS9nCpaKw8XYM8/reCRiK7sQMwtW
vxvU6DERWLKE4CqXXwUtkeT9WegkIgjICnm4Gr6gWblm5PI3BAb45sOYyOLVyyzv
BRsckdGFdN1z5ORDNn+/zA+1nuCOVBDfHs4Hx3MD5QWGDaIg5R+uMuOJZYMCFcDv
YWf8kuDOu4HSpBO9WMywZRrDSUsdGR74cPhpUt/5lowdtN8iZlmDWlhld8EM4sbs
w4cWlScYnIXl8Cubz/2b1m48FSPEi5m57VLel+SY4q3dZbW6qXwLj78YWgQ69uDN
9Jv2N1xnL77mm5fKZC+zDt/EtX2A9KpaEO4Irx3Xh6z9LMZhZoeCIDsd0HQ/yHJn
95BkWqPORwiw0qOpjns+iY0ji6RAvAELAzfmkoKj7pmNzaMFBfs1TpUuSsdS6HX9
i0ZVmQwaCodzu1PN3loar+ixlEhsERIVNcljwTE7rr56HhA/QMs8BxCJs5RTqSpI
6VTJfuGDWiVsV4lJIHLlhTGweGGFosVwbq0Ytvzsu50g5h/L0B4flr+42bCynPJH
xMZfiMJQ8dESU0/lxGanEoE3fnSqABWLAtEUOzd4da5SCKpoSOu2GAoJObv0bUWp
lh4hiayS9ZgyP1cp9hHShPxhP6MhXGbTgSgPhrMWLhWodWYtuwUKZVIG8wkx6nng
eXce+HxbkhoHvw5PyZo0eZ3Z56WwqxfG4aDFpRmcB+rsJeGNCOlpF+108gSBhWhL
1ULp1W6rnSAAN/Tir7pgyvKcqRA35dedznY5BPXBnrLBe8lzVIzsjFLGe3XnDC4H
Wm9ysX5uIB2Pfhg0XxxqxYYOkdzJq3ZvEndl7G9nXtXzcj8GygGvJYAX5g9GEpIQ
uXy5bj1IyAq/1pAbCjP5d1216/UgeiiiDPy+f82aZFhB8OqN+stWWpiilZ7ryF+f
Lvey5tJqfkQJPR+fRXLGRdSkVIKIGQxMZyuQLScVxpMxls9/fgaBw+ZdbKi2tHA0
2uFVcPrEdxaRxaAXv2devXwUDYvEhEEAALVOG7QNzpv7ibT2SUor9GXanM+XecB9
u7SoboJwlkAKlt+X+09gnyoQktSftM77fSh4VRetQPw7Y1Cms/i5LthzDL+ftWjY
YwW/XroKVTpL8FKPu4RfyKJi/OJdUvkIP1jzRB97b9qk9I4bh//zXGp9u6d+PNSH
UwPutJqiC0jecmz9IrIRbSP64naQJhCPxPRrf3aA30emfecUIoC1gz6lsaKmHSmT
GNlVH4JHYo9Fdea88gtXacAx8JnHUzkfaPmXC5/zuX7fTpchfocpKLVNSPepPLxB
1SgJpsXf4yHarBhDr9m3H3qkyx2f3SjcPFif1oaQkvX4TjEs3gUrDQcG5d1pQayD
K2GE7nAGe6EUWQo1/iJvv1dzQtVdKu/PcQONQViyoyGmJVpu7KgD1UbWCihQ/mo6
KEoV6nhLhBAKuKoSV+NRGJCGr+JJ/QJdIfqqsSCC24i4ZV4+EJKqlUqr1zcFw/a/
GQCjcJ4N7UvYrc/Us7N7XcFp7JimDC9Pi9M14+ibxEKNwb2SO6qPvHcIg2Zk8wEb
fxbotzMsnRs2RYHI0H+RYVtzIQ1hmvD3kOXULVetHzNp3V95/VzHZ8+nM82kcGj1
7px5KK0wuUV8q+W4i4YdcP0gDCnd2X0mGhifzOnNvqreVb15rQLcP8e8lOMgWUIw
ajKJceb8BlStKBe/Yr7NO734THa6UdSlJYEzBqG/5B6yp4P6xvFiFbzNgZ9F92Se
BCeh2TTnYMJDpJp8EX2z6ZUKl+zVdR52vWL85JEt5S2KgWhsw/Nmmg58JBII0bkk
njfbpTwnhRGAAd5GUjUoY5sy9enGpYNmJmVsxxo//TJxybBao6T5mGmYxmPq3Wa5
EN3xsH2vHvE/NdAAnLLgNhtsrTOQRBCsz2GpmMoUBFoCU78hUsuyBpP7FQhVjVVu
Ho6lY/088ONdbonoDYsstxSIQqUfXFVLk0YcBVT80VUsZwH/6n2guoIwdDP2XsgM
mu0i3v8msJ52dvmi1AGo505AcykkjtDbxgqGH0sLK+aE875s4HcUgwVxpj7xw4Dq
z6yFwFXfylqomGpZ+SC1aEJ7/UFPoc9cIm1h3EXU56OAs/Lm7hiqV10KrtvRQrie
clnr3iQNNdNJqIvlFeN2TFEq6TYpRmt4h3Hin1K3iCJrUQFAGVSKCUwTEeSOd8Ww
bzGBi8Cv0NjkeOumyLHfoI/0JhZwBtnV2WYX133Eagww6lBhspGczEhvPuQaQzb2
dFSuxyx700aO3ac4hNNIXpYVUKoDz8aGNfZW7ERhZEm3eVHoZgcSjxmtrOQHUheG
nXTxs4D0x0+f6mGT1Q1V92YJminVG6bT+V87u4YGvTwKoarzGYiFDBr8KYI4G8Y6
LHHGqZdfopvnb0eoJ0xlDq0v7Q/bDLw6cZOT0T6hKFyXOVl6bDk3MOBFZRoHoPJO
l6o/6DLzIPZVyBxTV+vpF6xZXJk2X/DDZpqzyApp9cOnn1Ixw93v2sj+MANRLPRO
bte1UdL9WzegNGahG/pEXWDDMxPfxq7S1ijN1XHuPriqcmHCS7WxVVkr5T7JuFuh
6sXV9S/hfPvVvY8QUrn0y3tjPx8APhFDc+4fQhftFq2ifz854tHQ4iC3rlN/JYYg
boL57TpjAcsmGiCfW1pcAzF4aTPaTwRP98WD7DU1RGwG9JZFyNPl5DMyH4f9sYeE
nb2nsYjiRqvx2451ucF5bmn1xugX3KRXDnL4/XBrQW53wZwxYGANtHFGi9yczIx1
AtHpnnQF4TSKk5HHwkyEWVLDG8Df3C3N9SekYOByUb4BtW2SKSkfGuR7XK/RIK09
9CRO9q9kp8G3DAsEgOymU6XgYMmsocXETOuNgjzvS+BjuY3Zaf75CUhEp23LOQo5
`protect end_protected