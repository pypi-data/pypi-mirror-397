`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17456 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQDN/EwIYTUTpfCPqCp8BOJLcpXM+xVOhwoOgAqi5qTUe
jZkDJ2xu7LltRjMFXcc5vfuZ/c/YMbhXcR1KvvgHcUEn3eNInjsbHcqBMPztRN9w
lHKRf/yr+Ytr7ZbWT7E3Ghws22cvTH9dLnYbrs7ixNQlIyEizwSBqcg03R6Z1ORP
DD7aQY5MRlNHNsw/c3bNdUy0Vy7mYxpCV6ljvncL+2J2QAzxl0PMzl1ovnyAtsHt
boNiNk9F4vIpxq3i07/KKogVJbAPYRRJGCtjlZaqnCV4Vc9Zxp6w5DG/rJ3GP+UL
BMMwefBoK03ISPzbzsg7eV4I3bjb6lnlwRJBi3K3SDILERDYuXnQTHWghPYd6Hod
Wfv5Egf7rN5MJf3bsB58tHwrV8QEOQ8UtMeAGLc2yoftxzEkvYvnAH38XOMSgBsu
KXULKMf9i3JD8A1iEBuoNwQ4X0bbt95YedDDcw+BwrXFKKf5F9mpxHPZOFQvV4j0
Erh4nLFCCMksBabriu26V8kRXDN//NkFFej6YfzsssDv6wO8e2/nLEYmFch5ptdT
aI1IopCA7MkuBJoli5W79HyOnS7oF/J2t2Cps+8VRkJmbHuzGwcHmncL/mStWvFV
ytNArZMclucZQF+dizuV3sZemtVZJYC+hFr6aEe8kMXIGtUCVEKxK0aJVT+VQjrR
0Cn7TBZ1Cux7Spv0E79k3B1QJepF2AFKAzLQP8jIyUydpif6oC+K9ken5q6cuDP7
hNkQtsbd9CWfeIwiNbWvPmwfRs0ZHdT+WqsMXJUGczTWcRPxiTY/ZOMWjxSmGGfy
cQXbbRDV7YnoZT9aTJ3N529wDTTXOmDzlLaSNQ86+d13ZcofiVNayBts/JEcF8Ft
lgeiaPDXfIRekQOjV7dR2O1Ko2a/M3zTvoMn+LSB0yWuqCrjGUnIbKlzvD5uc7bO
f9DHZKJLaLZwTho/x1fy7RxQ9zUnmt3KAQTZlt/69MmEtjd+wnKJByOvCXgR7bbp
Pc56TceVJ4Sdo9FTGAdWb+FalBQtfuxEi/9bvRQx8bAm+2DZGWwZc5WHHHr2dCwH
meFGWqFasl5ioJLrybJ/SjG6RPl3VIPtiN64Ce7TlY+t1G66j7wok3pkrOlxP5gp
Tgtzz4io1/0opB2uEQv7rCvzvzhmg4tVfZIkDYHTgFtq73UZTwy26ABEZOLdJXWP
I6fRQhssiKVKKKS+i2/Nw6ElBokbdMKpPhDmOHaIug5n2F7XPGH95cxxXrVLvcXR
S9Ti+tphlfDsEaWuit04KT+kHIKmxdJ8xftAFhy+7PDNOZ1yalm/M3KxyYy1Cust
mnw/kwidVbv+ttMQVlRHR8N5WTMCaTc1ITy8QblqLrnfUeIQ1K61wka08VKKa1uO
e22ZncfumI0inToLuu8ugq7ulU6XmEkm5eQjSXPvYgG5ec4uv7d3q4yb6tNIEcbZ
tIe3njr14XI2JeOBfBDqheZYuh0YhAu0uQZ3fhpF+KIGN5yOsGJj6WykR6G2UEUT
yljOgFUMgE0UIEGOTYiizTLqh5MIdfyCssQkKxOEB1azux+eYZjFBc5sbI/6Q63J
LYN9A5xG8iwpzWKuk5DWwr/0RZD0KZgL/XLQ0fU8lHXi+Gf7f1/VroQlirEmp0w/
iPw2k4jFoxLuvSCXsQkAVz2AWzvbZ/hrATCZ0L5i+NGpTYBJwx/0H6S300H3h/Fi
gSzk15rubCJDuMIoJsFHSW0tD13FvWhUG9u3uA01EgjaC2GHan+zEPm8pOzUkAsw
FlfkLohx4XhGa+xhZ7NDruRqWJFN7XPaR2JdSuQxSm6ZW3mJvHqdviX+sBEUJCKd
yw8t+/nf9HZrkujCaq1SWNwRQTgdgPHloYzbtdILapozwA/eUuM+blBWhfJ2msea
kTfJgfe/tMHW2Z1AUKmGDaj/7KARYJueB9Ud9Na44gSpToz4uCZMNvrpOKiM9jAV
SddK/yhVZ7UaVH6LlwmtLxjo1XQgyfiDkK/h2peU82iC5hl4K9Huvpep7lFSNNP4
sm2BR10Oz4RNRhnP/9T7x1sGbYWvY0+xyLGGv+LFIakzpi1Uk2HZ14R2SZ7wh+Jn
gLsn0fhDTOBUMNjNqMhkGUVw9oW1iBfODaXlH27FW13CO4lSjvpvq7dG52wsPJVH
oN8yjFrjJ9U/4ApuhG00QK6xSqIfwtTr9y22CWp5mM2d7v0E62FoOxn69NitLUFi
NU0IVB7RfSHttHuYmPEWG3tZDmuDKqKTX3AE978k3bhjkKLP8GA+OnBVtF+AdOWr
xE7zd8xgfZfavIU53+8pnHmY/mNHVHo6n3vN8SgoPs8EGJDeoYLfSzlQGbbMTD4K
ePycrfuf8kXQOR7koHY02Zl/3OADZhr+nKEwjDxFxesgRvdeac3Qwg5yevNLxcus
AYWbaI2ydjFfWp8uyN3gNCEraTB/flUB2fRJXJE1Ly/+IqeHiFr3JFmS5bb2Juoe
8g5rf+Trb7axR3YEtuP/q4dEnlVK/1B6kAHKgq9TyseBLxYYvY17bGEKIEeeyU5S
thwIQ/8wf5T2oMM+5/mWBdUuZJHVtLSqy49uHzBCboA3UI9pcoNhqgk8uRcD+CnA
MVu5vcnqtvPqvLvHZPOCSy8RbERKyur75wKQOBAohU6mHXzuJArOLlaZG9AR/345
jCXBvG9PUJM9QYJaMSgiTvibEyoG0XDS4hW+R6TCeuVlZPJ4RVWsd5/yHM1MfFAi
o1EOom2+J6NSuBkVXNyjq52ulcsKaokZVND4EDIzVTl+uBRWfgHYcTI/WGnZetSt
JlolDXXWCkr0AdlSdXehKOpLNxsALhXpKLAJYRRr5UkgKpeV/tbtFiqfXTfNZtGY
FP+P9Bb0aK/4uY5GdqaZYCSdjqsCa7Ftyv7UQIyU60xvGkw2CQuNri04+loYedWG
pttP8uJLG9ivdlKKdfZ23Lri9D1DjzX7UAG7z2fCdkYA4fGEOINw6aPL9lHMPhnm
QFf3CkiXbXeOav7p8eywApyZHqvC8yTaWctzyV2VJ5gpGpwuF52Q1b2Bde/c51eI
Bbp6WhBFJMVnZM1ePXtTIM5YGbSMLeN/Wk2iCM88S5V6Ox8gS7Fys6EsGPT9HLAc
QPp0EoEXVWECVeX2wV+tSw7JifJHQ5szs/IyHie9KZrjJcPi+iLuLJrVrgdVH50H
C0qUvvkTfKB1d1yJoXKd4ogFRf4ncF6snynQJgQPTjSU9x4/Mf0yAtB8cWEOHYXs
ZNHW2hqnqIPkkHLzeBu3rgDNZKP+CHlQ+/52PCW6KikHzLSJjMJZHd/8+E2P+02G
2K02biwt+K0QjSgOAoKQhb7uS1Dq2CEF9yDmD1T5it2ZhkZ+OlZ1KIrzaZ7fneOX
S6LrxwNtKANHu9ZSMkXkW/klhWpjfBr4Nk6XUTdbXmi/Zul85LoptC9gVw8ZK0ZY
eaJ4avZDgvoRh26/8ck6coqK4tLofk0Mtseo3oaXqdMY2eglpMamPP+gggYhpUhl
QozQqvxxEPA2nGginAeZwEzg8aVz4EzOxUHMxRF7zlDGC12tAkXr2xMbCE7a5rav
4HIP+hyIevr2XV4c18KENnJiyx3+tTSPpF8Kk6oP6wL7EqzLemmNWId+Ru6A1LdX
aCcIzgfrRh/brAT36URvzKXMEWYk98/g0gEiM36gkgE3ffC46I4sX2kfiV9t0lsi
FKFSct9Rp59aeujd9ojQrkI19nO2i/XL04/UA8VLWm35QLcgbFHhueaDSuTfFIMP
swbDch2AtCn6wMk0ZfzSRvQ0OvYoYobTXQpTY8grQ1+MisHGthWbdOPTbUN9ym50
+4FNbSQeAaebIz/fznK/PY1LRQ+a4uZuswo2UYOmPXyPQCNuvQ3wjRsLjc8O6/cV
vOpgSzQs+XjLPuRqA3NM1yKoxuUtzEfViJjL0EOGI4ZK6EFJzJ9EUvNkiDldbtHO
S9aIR3sw2mxchkEGymvfawQ31M40+drelw4XmWODME+cB44iw24XSqX0XWjHVuqi
E5gRurrXJKCAsWfw5Fsv3pcOvE8rHWKGUistc00dRGVVc9jnQsKsIYhvLmBnHRt2
VKZ62c+oiKqbh11VgffnuhmlpOLUh+W9UU3ezFOPWuaTa/a7X+SQkztYapQYdJ9J
1MI7yq/II+PotnWvh5zWamg12KrUJJi+qvFGBEQIADW6K9eWD0zgKqjbK/Y161IW
8qgVT52NM0d4FLXrnnLCZ5VpGGm2fzNdsrZ6ucjiOtPILMtERk17d4/ONT8Z1cPZ
jAziTVguWpHHRh3Gvkwzubq6dpR+4DhV7DYn6XJ+QUYcmkRY/bKMQJZVW5Xvb5BS
yrpZOZKSqiT+1LnJ2UydrN2NUwsf5Z2kJYiOrKCWDkwbPmLySU0ELkMMjjwwMQ/7
XHzExDjSJzY+hSWcwUsS763lb9F+E1Nczc0sfShYVPz4XbO5E+GjZxk97LL0ZmIp
t3YBQIBwS/ByAp8wO8vWJS8M6co3ZcsC/7gq1Z7vEVwFxapGjhWvc0fFRdziwDBG
Xzj0JnyVKVGocPgJKkv6xcXddF3wB3DNX0p2jQmYtSBoLhHpr0D/6WKF2L3ao19h
3I/rVnF+cHTCS1+hsgFk1U6W1gHIq/h6J0ZtSBpZ2kBd6XL55lrkE5y5CurVK2m8
OwXpW/5lz/lfN9I7F8yVLtc3FfT5dNa8CUBUw/vHqP7zQwZIwfCNdMYBk68ZOyuH
FRGbq1MIR+oropHgqfGcVolddmkHc2f3Sd4uel+W4QV6AmF1UFwix7Q2rPYBZumA
9qyG0evy69KduNvS0a8G7cA0PQmtXtN4ZI79oD9aL/l7uXlh+zuGYDiciilwwxNt
1A7VVfYVS9QJIbuB0i+nH1HuwohEUPpBmgc8g/T5628CE2HWxGxdvvfDOUbemPcx
YztLT439qI3V61QHkzQxzNwsJAeQ0+T9JkNsRdjh9nhRG+2uRRvTfWzQI9u97Gcx
dT578D+Bw1Sbx+DNMwbNzywueo3OjVjPZ4uqz+Qm79Bc6hYXGn0bc6mcNoii01nO
pBLYKBR8gogF3sXqTp+9esaExHkw3B9BhLRuuAct3EnfPHSFyTnPBZNZqdlWNj/n
aNEcRWptIppdg16NViulZoV6U3Udq7HRz6OErGz2WUsJPltwgiwbfLa9sXTZR8U6
svTh/6NvtVgky/akWHIn1IGCG4GMoMkJ+3tDt+TalUZGb6WmLQ4TJVIlZO29Isux
1UvAS3XWGxzcA7MozJyaydGhz1XztRZ6Z7O/vWSeWe55gRtQ39oLrUbIawKXGvw0
XafUCIvd6WTk7pMf6tal5iQADb9wk0qObml8uLvwZ/7MJOh/d9RQe/3GiZAYUjeL
6w2NjkTmEY5H2rADc+gpJpocQL4HigJuC0oUiVnMf7U6D85WsG4TXDSQlF4Ebggs
7OW7PNW2YTIEtlCeyHgWmK4HeLhVcHG9A2OuQnniGac8KStJUgwrxdJIybPYEQMT
yLPwLN102FGdaJGfzDWZ9rvpH60eaflDVAg/qhWrAMMU8wfzi3Htd4uzOQHgdnKU
KZWhltjJ3wbByfu4LrkYaRtEqrpCKU/m0RwFlRR8m6WjWKCyhpRrPHU0WNmkvYRs
eim7ffgKDKKbZC2G0qrREdzi+sjXzCrUlVviVmGJZV9KpuVdiJ9uMWtQwAngpJnU
n8rmO4svWG15LAYezBIilLLsoVxgZeGCvaWbBEBsCef0efTMg3+KSqLLP9HgGBzL
BXL3lKr5XHCYlOyk5KBEDQwSUtGNq26EGmWEb/ETZAwiLMK83503K6867zYu+e4w
ZDfTp7ToleoU3j5wEdKJMDYfW31nxxP0WgghkztpStBTYdG9pNz3SpuovgGT2E5i
HOHQnndhC5Pn5JumhCV9llvXcBCU4lEWzj0QEy+fvEkYcmxJZ+M0W589/IfyWAYk
snWfKrxRQP38aL+1zpW6+Hk1bRKs/RyFSF8wAxwtCut5zFkNvddR58n3owkHiQL5
VkttquvmPK6h3MLRTyjuKegkn+CG3EzZ0iAhxaUfJbvsUmbvPKWAfoBO0GDFBmQT
Ts9oIk32mdFAqY5LKOMlcGJSb+XtFxYZgw3UkA+hLVBKplYk46yTgWfbtDOFaUdq
CnQoVInW8y7ZSDtFi19/DwNmk6z5mkIP1qNpq0BF102Ipp407IAqFFBlyPXHNf9E
mnxOnag6c+OU4aOmglwdholGWhH9+Q1m2l+ML9BM+EYCVQuEGSKJaEkmpfZ1rFr7
efjOcBzvts+q/Xz+ucI3SqwIjg4bHUHGYkJzZNslpEx+7N06xVzZa1vPg2yNbM5o
ZAIUPEMAfpDVyDGkWikBKRIg+v2RHDgYrVfv0ms3rbYpCCOJVeJppL6KWFdTxT0t
WtZGMiwWlipqWENWBGOBnnrROIAzt7rXUJAQoq8pLMqYHWzXzpuf5ILYRnxM0+ql
6UMwYCDhfr4ZTx+0KmRsqBt0YiSkyPhq+WwRZv/raIEkfp1X8iS57AEpzPujyO4s
bgPeKGZm5NcPddMIr0XsWQPUj/cYRlcfE3SaZlEoIqPsipz5Lm6IpjOvE9QLYFGB
c4xnGbPb21ll93MzrWefjT4pd5fnNMcKifQeEWbUa15J71tcLnvc8o9kBukelocP
CLTnA+G4R3mfXoKinK/YtIDEr9Spf9VHFWfeuvObTvkBr6mQd+L7913JTyc7o3KZ
wEgVu7lC4wY7S8uNEgXrUPbz7NJpNIIdrT78MVGBK0FNxUSiJFNtIuDopPx1h3sV
L73VHtUuCo9UBL5QQAcwAf4HEL+R7Y38Css4c9lrGagMZ1jaJfgqil3/rJr51zBj
UOPfgrniNnfcjAKQJBt9IlVGMVhBMuYjvOpVSPEqctwvGxXZQKxgb0r3cT1OqeVH
o4Rc57Vx1jTff8qG0JbI77XlMfxuvGsckhbKTzTmSvwqxDPDrm7Gb6HU9GXOqWQc
EivU6JfTIYD2E0m55VF0zzbUaGoTevWzV/mg4ujPA+fqGb7TtJpzC+Hw434PScIb
ZFe4yD/mV1qyFjyS2Vn378dG58UgMfL3m58H7WkdfhM1VieXPWfcgOgtI85Wx0Os
f8RyX/lIrg1WRC5dBHDhsBFiSpKtMt0bKMUCeKNYQQxDIs7szAX+fVcUiQ8OLc5y
+brh9ZaZQlMGl8aoIjtygVac3aI8wa5oRXyp1o2voK1CVnEHS8V0QBqGPzL/WZmv
yDCabWgi96ffAAvkdcpSA2kaWFKzTxf0EQ8Y77xLT1/YHbNbKpD1CcJ7D+RrUqQ0
CASdhOVLl17FG+ThN/XP5+jwLxAokM50N2X5Tw0cp2fDPkBysB9VgpgUgQNdCzTX
KgBWVaxq/v1dtPjqLEFOl1dmnY53CnHKYWc1u71KpgEHlQ1nfdWn5XRrGpoo6jEn
sQ+eZ5booIIRVhyjrzTWOFET3xkyvsUyVMLztRuUD0qg2ky9lo9AvWdljlYsRPF8
WucQT/sTngusd3jPnWLJ+734G9F24C4w18+Mmn/zeArTt7hUnaNka3xfM3Vfs3ki
hEJivk53ahZf+pF1iHZFvOQE/phFvQPemmiZD3uyy1qKTsxooul9SncnOx6SQk73
NoUCgOtI4+enVssrb+auYphkgGkCfpdxs4IOpK8vfmX5FTtojaV9JAqr+a5sZV7A
Whym8E8ht56dnr1/DYJO8DoCN3URpmkJJcDF20SrCyUvcB33x3jxDiaae7+0pvzV
tSl7fvQ3QZTnmSU5D8boDKqNQpJS1jCO5g4ql7r60HEA/xFsX7GYrCTh1kqb3uSM
NB7GOOySDTDPuiEslJwMeQy39qPmyZc1U7jFxWZP2dq86pbeh/wvL8rwZmaMerW2
IkOY4rUlVmxefJAtn/yT3S690ukUnsohV9kyICeNeQBV+EYTXNpCunV0vwPK5uN0
Yn0SR+R12RsVLVfAm9NuJLtMHFpVthIaGrAvcCQSzYfNiRbA12Z4t25TSTl/p96c
mPyVoibhbPdzoEAIzaihPi+2X/oW2u6GK+z91Hqzkm968nseM2L+Dm7MfbvXjYna
HpHiOTkuJVzxcKSgWvg9cYCWpA6iuIUrU9Xr3mPm/AfaGrkcmQFZX53ca/syO3PW
8KAMgMjz3URZZONabmylfQ9xxRHBaUZzng8Mlg93MCvxYSUE9fECWMneFJhKWB6P
Mbkf8DAFdxOu5qsSVNHF3OANQSDVUc99u7JSfZaeuyXWx2jCpT9K95DquSDisiQw
eg7gIapmaMXADbeWA4MwycGDw/P07HGPBX1dZyCIwhK3gE5MsYWeWHAoAesw6Q9W
iJtkoFvyMnzHTVu2l6xsa/34kW1VX5tvrw5LXT5cC534Ur2ogR57oilHVKcgCtxZ
HbCkXRI9mZkBOusuLwBaIVq8fSAj2Ru/yAqaQ9ZaWwSOzGBvigBoGDN1o2PJPBh8
HBZlnz8iEcvqLn8zqP4ubZyvVXdtmO5INPSPlz2NlFAEmVmzU1U3gtfuCGkzmQDo
a/lbBt8zJC6Ap12eZEUFxuoSicnl3tpOhr77zBQnibXRZ4wFOaQd/4/BMz4l0I3I
UHmjQx4mS/3tMJW6fILTl25kktMAdebQWw/nNgDC0enyORj5uayM1jHYdYVrm5hc
gGnxArSXBXAGT9lqr4bNRqhDHebtsqi3HrOg33kbAI25KpoCYAh7m7uCQIVcb7iI
9d0prZDjN2sriKI9EgopynR1G6R8XiKp8p+6vcqk8CZtjAE9CTvdXQur6XoccPGo
WFZW47yldbP9j6EQR+TczRab4kCBBwQxvb0wpJwBAWLNPlKEps3KJUYPjnH8cfDA
rcfbnprCfuaip4IWNtoDwxQBFz3i76331dK2YxdrZ+AP4t9CuHXC5Ppat6BLkxnh
O8BbQN/wacWnVAZFcbq8Dd8Z0L2jiGuBqETtNuQw9XTQb+hdD2s5UvWBR0Qeb9UA
/ZHi0nAMabzsolBZS6bQ7+TIB7ZPlvb3JvA20hSPe+chbKLZ+bvkuUlgMlJleNGs
Z4B2SN6GpdTgerHqOUZCWoMV8ZrsPvf5o6CzrIvTlowUMoc9R+zS7KPrfSayyoJq
FCk36TFQkqrWcIcGuugmBTySKO9ne30oPgGZOUwahOVVPF1HjcJvs7v1Jn6l9EFP
KjfxQ7n9PMXNeUpj343xLju3t4lxWs/g7OEPIQYf3B1kOoxXTEr6akk5y3evhf9s
LTQJaIiqB7vsn85NOswgc6Z/wGzgnYJjpj5SGeB2S+FvQRqsRZZHmWLWNvZqSKNC
DO7jQUQHfDZkGbX7Cv7VL09m6cMf74dogsDpaBstRZmlKVlcZcup/G/2VYVoGpti
NhZZ53jTw3P5Nv8zk/LYJ2bMeFc/xRQvR/lEMydRBH87Pm+pCoFr75Nfk2jX6xLg
M6CBj7VilWuE2IYBNJbpp122ewZUFJYXqANNAyiK5M2agltXt8sQZgcbCFuK3Hr1
AJXJtLxcVQM8/kll8RDdIgq8uXSDGGInVcL+vmr2en+0K0TB7U5kdpOiEhtxeGCC
Kx2VMvVsLYk/i36aRjvNlGnMnC8ZRmpYSOAZDFaHXbeXqChWcs2uTKD5hpMANXu5
92TBT9yfslJZSe1KI9vI30S4+0FHNu+OIjdJxvLZp+7Mk0mj527/U51G1EZwxQod
2eBTPqFkJOnvrU4ADymKF224kso7/ADQfoTu7uasqzs3/S7oF8w5ZY2+OQs3NShV
pRxHh6PwTyc+RgIDA2/AFEPTn9Zps6oQSRT5GWXNybB82ok9TKWM48Y21OOvYNgl
pC4245jx1MRveR+xb0lv4PJrpmmm6ubnFxpkfELb6+jmmYstu5Zf+H4fr5ccGs3f
/PmD6qh80tdVIxdG0P55SMGirmIk44xHzCpggleyRLN1N7GaqtHJBXeQwKR3He//
l7p6dKFV8TcRIb0UagTYNlXn2pNDLLoJXCtrboa6R58R+q9aYEptg/12n0cQ6XsE
xKQGyPIDMZBjj/ezVCVuriEbxXgaz54daM99nRQNNnZ4VRclFc8EBjMZJ2sNQDyU
Jva8Kkr4F1I8TUGwnmHRYma0n2bVGf5uQqJvqWwUmNUkbnr07qm4ZoBYjksuWtA6
39A2VOiPPchRO9OteJTz2imXnnSa2lBisoTXMYXZSSL1TgKaSq4/kjAK2RsIPqzi
4QEUEsEByECt0x8euOg4fYZ3myBmXsoYlRANusHOm7H2D6EwZ8uZ7oyYokLbfURV
uGolHSVr3vcN/LuSPW3KVYM1Yw5ecYSgO9BiqKzjzNeDen0j8iErk8FHE0n0HZC4
uioCfAjAS1Lox7v3w7dd2m9eSruDND6AlylwShl3m5jYp4K0s02eEV47gqDiBDW/
OgVWsnWzvUEAOQoPc0AWVRWCcNuVsRAr4zIeiq0k566T2bLAqwrdS2SkCOvlJaPW
rDS2eX36weFspViPemTO9d3RA/+R4VGHKp3bkzPUkugJnm05ko/XDZZYicxqSw1z
TLCGT78FaM3xIDUgeNvCKixjtkdOxs45Uw5EWUfGNC/+XFN9AmG4S77UDpt5b6JW
Zel0WPYNAZqKDeduor4yhn1YBnmyhCio4pZgKRF68LqV+FCD8ETqaCZsiX8gvh08
D6PRlsBWKaazP1I13+qgqh73kHMtylpFuSd1lCoXG54I9bKFi8kCHnYxV/g0JiV9
2Af/9CzIIB7Lespx/LghEms0vtPTIovT+NwuHFX90S4Vp0RafvUM0O+JXp0kwckh
S0rSR3bNSMKYB4kYRyZhh9kWuHx5rOUYulYXwskJ1XoMHWq5+UxsD4tNTdocOmGB
AtTMRhW7uQfxAfA0N9n1PLvddB+WGCvGsJcC3vk+i/93pdqnwmtVv4PVTmNxXvW0
BsN7FvjfW4kXI1HrUYrSs56gXR9t9VNtrJhf+nCiEEUc4Cn+Cw1UgUHJNIWsilYP
cvlmwQXdmkLUZbRgjUb3zcVqEAQUp/E8spJ2x8gDUy+NYBAAZWv3uln/a8I9O5f0
RVB4oo4vm7aQKGllVdAW41/fJ/IfP4Ld9p1HQna6FEDp4DFtiX6kQOZW8/aDYd1O
d2pcwj5m0ONC4TxBU6+IustXy4wJoGko4cJ87d2kHfjMy8YYTwdjIekoc9OUwbg3
tR3BglmGJJFtbPOrle4mZ4H6iYSJYGA2rYRsgCGSq7PbhksOIhUpImjylWuxtWl8
lcFFavEynuPAyDXoWwDQF66QK0d1Bau7ioIRXrRB7nmGFr6xixoudJ3Wkby9+XFO
dxrtNeHG+eeI3fwCa85QQQhNQSd+efjHg0B+YUpuKe56wOv+sZLtRO+pXcEefjSL
4GA4K2ntA2pjQ9dxU87UlXnADO9fQvoDEirjRk/OxcpRZY7lbw+bBocfPuQGXrGN
796O3o2vKjePSO2uD06EmsIVF0VvYdBQ85hc4WKqfUuYrAQRDKX0YVpFn474KP8H
bnXX8xIMSsTtUkGlvM2ZKmGR6xVGqmwjbpfWGERfKYfEzuLV7wlk0YSMf0ADzGWV
MIw6P2TwrY+itQSL7khsQlCYecRBM+YM5Ioc20qWV/2I4iAQlo0hRI2SxZYg+sOe
aFCaC2/K8l+L4Ap/xARXSMasIaPp6bwcJ948cCziTCtdpoFl1Xtgfkb5QfZqqsJb
o2W7q7y0ADclNgSply6b1rMrBiEFBb0UI1GOub+47+TI1yE9mG+7xFuEr6X/durc
I3zSHFp8aLPWiLqlpGVjI6zsp39D4d0IEGsbIW5EB+/YKjt9pg/3iYHpjC3ismUh
o3bZkMQb7rLjVHykOZKJf8AR4gSH9dFMniX0hGvhgRm/qVH4W1HzBMA1wzh9zGec
a7Mhztzi9oxHWn+KSoPhIUOjR3JNYWnHoOkgvblmdbYcyNEWNQvLhgjwkyxUjM9D
xlawLGH+kNsn3G3ZcyUgNGGJt0/tFw6U7bMNZ31GxgMcsT8Ij+jMhFB4f5JKMo7E
T42JgmFIb4cO5eekVND6LQAtnB6+o/4FaUi+qJVszaC+gUYCS0tL+RG8pnNWaH/g
6JkDvb7uax6ttjRX46SLG+9KsJgpDZ3/OqjuB+FQ77UIICEdlNWn68XyPMkNl3yI
s1Amank9QoNEsBD6yy4ueqxFZPHOmyTcMr6bZ3OFDcLHUJNmHIPH146eMLgi9gGe
99KccRYxQNR6lhufYzXL7bJc3W1sgCv3mVjXcDrAxlZmVoCnqTU73QNV8/43lIa2
yvMBFyANn+Ok0E2mRjuy74kW+G+TjDToC1ZMLdpGHfzORC/kSG8CAWF+LBOspnSy
bIjkeGrpdumtmyWTVgoY4S7s1tW66XBNNHRtZtzuC30t8C1ijKLTlQ/3ZslfV/1l
uxY84fd+9DgazCB7M0Sk3nLRPWkgiHKYbWOBP+jLV5tcuuA8B0w3z4erUuTEV5pd
BoUzau7TiLimLvGRahCukrbpYfOOz5pSLDDI4TgMw0VnFvCMzE4cY1mPNZ22nzX7
O+2NRsBbviL3vvdHJmgijDZBdEw4E2N+h0uUa2oK7QRWi08ygTuiarNA7abKRkrh
HzkVmW/icK2DJ+sMxVCWWmUbdAXy//cAw7NLvJcU/z7FlpfpiwYWlsfYLziesfk6
kvI0Xj/5hT/WjG6K53xOehj6yKMcW8gQDIDWt2dxQiJiX2VngV/WnYnFkiM/77WE
3j2zfaquxlhnnrGXO0Wm19g3k0YPvTOYNDoLZ5kjQtc35E1LtwJ+wgJqZ8RYJCeZ
2t9fVEwu6ceFoUxAXDxIlRO0BSqbMbVsOjVrmRWWMiouOLDQQInYEkGmjEmVSmmo
QTrr7x6xaC4wJJJE3ypUVNJFdhDytJeqUhU19ghtd2EjnVsVyZW+vu5WAn6z83ff
A+DdfNTBrI0XHUEbsLXNAv8CR6uNZr/UyY3zxm6hWbnwZ+7gAft8S+xg1wZeqM+W
G1tx9BCk7+y7mxzRj/k5KYgeBAbklt6IvURcPPRoXo1whT1tZTwIa1hMSpIvfJsP
HrH6pWxAEfZ5WGlovTsj7qAX8zYnGVApD6m/TRBTuDje1uY8h0067tQfmibBGKnn
J49jfg5nJmbnT9fHWG0JC5yV8UisxQWEcEpUaq5PJBDwKj6MRLb3DNsS93cMLUw9
lohNp8f5KVQEPqm2uiD2nGEcidMme1GB/mp9bTpVgkOwOKLL6cVa6q+74y8FIiP1
XPobos7pKsMxGGTbNpHMuasxhzard9bFYvzrHX1ZYWBiGviqIseQxK9tc6J5tOD9
vuZE/n+Iifm3Yhq9D8FJRQTRlFRaoSA6xR5/woA1dELSxRUc/t7ZJu4Z9Tngebga
Wmg9jQjgQoqVGq2b8ahD80JRWB5TXnULxIf2GuyRq2TWkHMqtwF7tagZ7mIkQm1x
vDC/Ivlrq7JItILeFSrUCpxDY2KqneVV7bai1OokRUtf0nVgIwnQHwYoUs2Srb0S
gzaNEjplirJpjlzEkejkzwit0OdHOA/pAxbhKDTXtAi0j0xsjpEQRNHqhHREmuB4
77qSS/UBX4/RliNdUzFMg3qR5OKzOGSY0M1H1eg1wT3AMzfJkQ1Z5w9K85HeOwte
Q2dY6kjtiVJlMfoX02EC/NDiNV5V6ceKxrAiBsYHWZPX2TH/6qCg0T1fuYUG4uJJ
latYYoFfP38Gde+T5+jYPaB9EBuMF45KnNwzyWqm96bhvsv3L5TtbwxCQoeDbXWY
x/or4+AAdHBmf0Pcmaor8MfXSTWQJk2fC8b8stgmkgOYcs36q9utqdFcLu4ikKBQ
1QyYu+txKInUpTf+VBsDJp9C1PzHl+ITuefNgbmIASFMdjc+0Eehf8J2dX2OiWPo
/fGnAY9qOTl554z9UWVOLGDRrAFPY1aixs3yu85ySEvrmBSkeDcYg5T5gf2PiHIm
2PdXDNznJMqsKAn3LudqRU3MG6Ppp/Dng669B4XLp34oDelzMFRtlUKetEo3YTAZ
Htw310Y4Zegwzqx+Tfm9haB/AGJg63UMkVIqSh8l0G5s58R8F8FGMZm0AzG8GlQl
FGUIqRqxgMyRhM1wiVu+pQv9HRuByp85Pn5R2wHjr4Ik33v9+qAp3MkdVQ0am35z
8M7k7iCubYauchVFlkwV4VF8skCN4lP7PuPqwvxV0iloNMa6Yh9b+0w+dbrF2ULQ
dAftzU3guMndH0Q17XlpaiGR3s6nWRfTicgo1cqP9B0Xme6hSPahNwJawO8o+KLw
sRzqh8otylcVYe0xMGowr+Ba8mZx93MIoDJiZTQgwBNqJcPOqpboezUXeJbwR8rJ
Zcmtdmm4ipht2ce+SIn+GmZf4czotlOc+9RpUWfi7i52UmbG2NL3A92la5D99fpS
MV82p/3kFIHwCb4ZXdVFGiM1m/YM675GM2MZvik5NseUiYZmXaaScF7iqUu+2Y3R
byS3e3HItrctf1UlC6c9s11N9wAyAUbj/UsNPRFaZgWZ6MyVTB48p3Z8pVaBbNit
4k+ZEjEh3F4Az30xNrQ5T8J2c9DYqegLadc/8QR3fNVsNNoSdAigck/kCdijdHvL
c23+oiAceoFrHjGKxJDRQPQzIdltNerg03eZlg5or2d16tP5/CYkYmBYl9FD+PEF
lw23LgSllcv1cy2x7rNKYe1gRK5WKAbHaWchfY8YT0eDzPQ18qsHuKJGb9dbNEph
Y9SP5cbitRSjIjjAUsubXsA1Gw/gbMs5/PCO0R3dBQRZPHYMB7ZrmbOVoKAuZFPm
l6RiVqcaeM7X2dJOaZVt3Cd9M1D9AoH4v3PJ0AmY8eho+wtNWfQmMs2+njFqp+ZI
cl0bFv0f6Ro4txBLpmfKzjwJOrdUlZ1YtvjyPQ4kNUwvN7D9E2mwDN63bw9IdiWo
o9wq7vwe3YPwLOWCnENDV5Av6VNv4LNmUZarNy1UvacUT3jbwuwhfWLUmPZzGfEj
VyxAr7SQIplzdlXEwoYTA3aiHI+6nV1HMP7AmK40dDAjhuWysUgT2SI4s8KcjOdq
4MgB1e6REw9egBbUOJ7XFEklYpvr6TjUMBzweLlc8Cm57wjOYkEXkWEvpskSLK3s
IPl9CpB5sToinzWLtJdEcq4pAq3ulUCCy5gQuFxCPGNnkaoxqoCaMz92txmihIC6
GKcKN++ug1uokzgOCzBUytveIvYQRzrWi001aswB2pd17N4RPbK933bTN20FOOyG
pUpkp6y69islC/w8N0NDlYvpGmqfBED7dpBQZdsqf/c6PcfJAvcHypKVLJv9xcvA
I5/qXyhEQDyR1u9qjf4ktKfGjD0fdYazfEEYXGK84k1pUksMX42lBw2UF6W/nlE/
PqAKFzUjIPkcxNxDc1E8OGZgH8xEHfq1+6NQE8fDdgMYAYUwuQVHHTOLSuCPoKqq
htSTZmw4J6nBBizqP/NMI2PSL6BRnYBA+0CVueb6g0nr5VCWs3uhE2CXKu/IULLv
Shw9g6ePgs+n9g0x/7bJPdFasRgnKlZ+c7PTrgI94acqPqWhFFsAV50391RCrQyL
NYFiqE+riceRy5392vAycvPsPDrqBxVohYZbU0xzqBDnCQaHXDTVhDzzwXf7HoK4
EUT3uvFgCwk/f12tOLmlwt1gHOefi/Zu5riJWbz56qPtelCWp4h3IbFSsw+IflT4
/ir3C+MvadUvL0ViLX7lA3MSk07kazRadKMGhNo6oaC0txWMRDuMaoCs4vqw0LrU
0Rxa82RuKhYXdQAbuPgJYUJDqJokJJA1ZLdlmvsrwOEzN0JZb8aD9GNX+oq3J0Xv
IdbOOH5fNc5dKmxcgSeUrc1+x6UA7YrcNQcPwhLLyez+O8NxR+YnezkKMSf0aSEn
Q8E0T4RDd4Ykw3tonqVWbovX1WYfyGjoND+SO1FxhTvYebHjHPZFPv7mJDvpbAeL
Hvv1L1IB5Pv1Srh0rsM/Z3c7+09E+LZVw8iHQ8VCoXhYQvOU7AgfmUjoB7P3VMFo
vrNARRGADBtkvG7s3oiNcgYg99XKbudLRLsSV7e9uJ6r+Pq3iZxENraSWdCxzThE
h0Gq8/lUiGUWA6i0+Q8HbhN4C1WtavC1qmQ2liTx2pfNiEmLdAS6PQiIE+hSuRrE
z1Exyk7PTSwow5nSaCFlSOGMoPsR6FX/u4lMYjNIt0l4/fSPUwCAt8iaO+C2nJiS
lUd/BQyooQWuUPQy2p2ZbAz6dPhBhXq7omcZUozMMIs7QN254n3lzAs3XymlneFS
d8RjfMXwA+Hl3WYbdYuekyKWTbN0KcQ3fSnUpGoWPjjOZ7xzyRy32OqFZqZytxvY
X0SKUW3b9LT2QeBbEdIN7ghSOYV3zDWaXfRmiHu4qeUZ8GCXQnjHvx3FlwECFk0O
NwePh5NplWD+C3ix1wbAPT/vj5Jvbsfhy3+piyGU5pv87PxNJRy0LkS4X3MjYhk+
uyfkIhafAUMDakNGOdzIIT6MCyp80Q+tXWV561fi5HvyILSlqYpbzCpYI7FjAbbc
DENG3Ef61+ESOgEvHAV+QrimePxE5UORyhLfARWY9xEYoJO8WVZYYHR3hJL3PqEZ
YCraL042Glc6OOPjCdxJO2XuN8fysHwl6xrHlzFMDoCa8dR2j31ny3Zpno13HHLD
Hr1sCRCOIVNZU3k4VbB2RJmiL/XCQM7zr6i8tehxydiqrvmJlrkjC+xXjefZUEzd
k6BPccqxiZwTcKGdSR1FkXLIjCCDESUUGuf3KDL/lbjIVY2AeXPXoXTE8k0JbA6M
tSH+dg9VPl52N+M3tjbSrD/iXLRVAQ5zO9GXgkMJIIRDBXZrNGwmhNxvEpW0q6EZ
++acxkY17u8IxLS6Ve93y3NGzLWJNHZ+eHys4InIF3rCxg56RG7vYuIZxiUPuK/5
pmMZXgqBaGtVI5L1SPK8kFQFOxFOSgQ1+jHxvrvMzdgc5U5QGdDNxQYM/Cz8q1a7
IYp7NNPN4cWriW7MF/pziKipA94Ly8kn7SQRN2h+kBLy6onXsf+2PJW6ho3FGPZ9
w3yiaN1cniO7n55nPvGNYg68ngRk7XQUendGM07RIC3CX9mXNrjRFEq1qRPRrP76
vr7TtfVUMWaWSDNCCVM59pXdGDmgzY7kXUWhpBtD6qwLQd6IPE5f6rAwVfENOgx2
cVogXFS7gcXdcnO9Lc5hpbBs0sfTh8ssDSM3oCI9UZ2WLH0g9gbFWtVzGTYG8M1R
QBEyT5EFrtc00xbpmyGEeRgsOLLwY1MEICJ6YfPx9f8In4YVoEAK5Af4ZDAud6oI
wmQrvBoQeYRZOnvJHVlONGwY0RPXWDVJBfTEI/JCb2pjgZckUmokMsPIEpNsqHGb
ZmPDx1HuDVVyrPrlwuEn5E/fbfzqb98MFpqPbdJee3RvC9ZO5S7Dsgk5BnpYHpSJ
eMDCklxJrlXfsBXycVyupQT0OmcCMTaOB592uGg31lv7hR75OjZ09kAdaolJlUL3
UxNL+Z2ADYeVJR9nU0/uHSenozYWQI/oE5R/lMSp+p255XFhl356Jl+ZHGk9TyEG
LqMpT1+2fT0PLMkbSg20a1eJogtFoMd6o4UqHIYWBdwikI0wjh5WKiKvVBu5wLc4
n1yvyJhto4M2XAYssaY2iy4PiNmRis+leSgoDphRWL3EDL5bbYhAzjJeL+mmz0AF
U5Dypg7g1BuUbYLUvobgV1LiJd/nx7aTJu6TdE3isG2FvA/W8qBd2OeEZPLLQuaI
E4xqETjeZDORG2OwBeSJqFpSEg1dwkfmaVCyRa/Xe+7CzQtQSuyfsL154mCh1eNU
u7Rc8az2pZN7I8Z+DXcOOQNICoh1SWCLFWB+wxSRy0miHX9gVX+T9MUOF93rnl4Q
4YCfTtBTEZaeSzKF6GNoaNhcpTHl/UI3EcnNlgzOMu+Lcze+ueamETH0/XP2OWsQ
Eikf0Cos0spp2uLD8Rp43RJBMvSOmnehyr3d9KDyCQtFFLBQcsLZI3NsUELcEQNl
2r19uaX2jmZ2XkZqf7vKH+KvkhxbNFMTrOYCr0+M9Ug3xy1ccCEc+nX90za/YSTe
lezShGnAzuVzZTvWetnb4rbj20K0ByU8dEKZoOYZxuYxdZ+TspPLE/dUMvDIXpkg
LRb3xtbjnxLel8ibmH8r0sJ9pEqSTs02VHltjZauWVIO+623Kd3L2XDo3hE85w27
Aidxk0T7cBrPC1MHcDkL/aF1S4ieHYg0EllrEHBlf2LjsEfHlsASRLzUot1ttStD
DTib4qQjdhPM0JbtmGuhZBIMjoobR6YhVMjEU+641A2lxQYZ/7WnbuC67FghGEtO
61oqQNjqh2XJaTwrYWZt9i1lA36EkyUfps4+pZiRkH7lGQEOfqdOwF+HEsdH8/Qg
g7WA+TgNrpdH/F2kd3TpSiVJtnMvoKuAhJMK2Sr3KvaeCgSKgZF1hBfJ1rhXP1RM
evJ2FIbKlM554vXWtjRWODQiOAVYy9+Y1jl3mm3uAJHYYPjpyWaPNOQS0qwmTpPC
1yTYHoY5BnrYby5tDIsVY1wJUJ4mBKMyZYI3pvpHkCCBQwmNXtdbtEyWjd/tRf6y
jO1AhTNCJGlGzuATXRxGWk0GQ//X+TO3gC5Tiy2wBzossy44UaD414z1Ew9bAA96
mz72ibjflboDbOTNDWH31aDq+8lP7k7jqIPr0bdRIjwBTLL0/k+dGyxB/aGzF6Jj
LIjKXve+EUPBYyTTKsHMDtdVqiMmnCbBQna8bRIzkvBmqxDS/EnoxsVRAIg8vRFn
Ei0wn98GyzZ6qNspqlABXSnB+W5fdEMJIsqeyzbUbTPxLPL/hw1DN0Pc76t+MART
wKCGxReji0oU6E3B0Uy/ksv6K8z8s13WKGFYX2NQouTKMCo7xzLdE92RVC4HaxYd
CdbTAtyOz1ihxwBF4E9vQeE160zGbLi5xXrC8MFa7U6gCRt8kB0i+o6kctCfcq8t
6t6eXd+Z27A98TONNybm1wRN0ZQZ10No8+lIz8I/dXvUAxle8rpmRK/0f0JtJriL
1v26NluiXMQvVx3UBJxsBs8XWd0mJCfd4vogRUcrbhG8kFq9fBa/G3Vkm1Pio0jj
dBD/nuQuW+Hkx1Z7bFJiDQukTTtYLN5M3s3cgebozgLsnq5vmahSRhSHcjcdEuwg
mtKbx3yQEe9K41UIf+39/fNWMABUC4L5wmaMjjjDna1BUhsWws8XaRiX1NQkF6Kl
RWs4XnC++/o13RQnba6RR8mEfJYWE2SWTLVDrB+NUoNTS0Zf51WYHQlTbz5Wc8CJ
kEYkdkeLxhHM2imNHrsw2MB1TdG9N5R5cluyYj5oVzyRfH2EozIbgIPk1a2X6y9E
5wcEcV1p80TQSF/fq6UNILIX+/bdl16oo3O3uPnDIPE6km09SzyEOJm4wd37WSBF
h6j4/BUBcvg9r8NDeff69JB9E5CCfDrxHlLkYFaAlFCvCqF7BGWTie/TM0H3w7kh
Qy0FlvZn9mubx7l1hn5Lvb12MpNwHLRkmV8hsVFOGSG5d/yS6zjnuqdow1UWFXmR
MJ8GGtGObziSVQxAjXXT9YOmF/cjfunDwZ0T+350Ewp+YXQsVIBzQgZGfFkk5ZUx
1eBFcEBtpHczQSqwZqlb56LbwMpClXmWuRfxarHza9rsaMqYyGgWhUDVHFvcNmA7
nhOTdaUVCfhpjkl04V0U+h0cD3Vqc30kq+DZbdjeDRH5XF/f/cKZDd2ZQPMhUJwQ
HhktDinkJXGOyHoRDUN+YK2JQZQoQ2YMElvtVATjxlHFOnp6O9R6bW4nckjvuZVY
T4IiA1w3oLjm/wvb41dFTqmQBQeAp+eVB63xISJmdB3o5E6wUsuYViqv3cljJSAn
9fk0ly3yGgszRu6LCw71L1E6OsHwNJwS+E97/ftHo1RMxBtuUxh//W3IDRy0IzsL
LOCao2aRxbuIgdDTyAfxjijegaTdmlZKAG2fy6D6TsU6XTrzrCzdCefOzMSA6877
BISl/OxpZuHH1p9lPHEzQCHrH4QrG0xQzUsLcrkwKGsqEkHrOLqAe1U58vA27VXr
84zgXBxzlwfdVE4OnqU75skCjP6fGJ+bOTHTPcMZ7L8PgqNwo+lyDemY3Rq2tnWd
da3MzBCZIHyIt1+gU4j2BUOpt0+hqelCMMT9JyaaenCs23V/pwXuzeD+eQQJ6T/S
QpThCQNMP6/lVJTwhWlFzffqpODGZvy4426NFfmavO2y9p7Vg/wkfLDVgNifZ9h7
kZOcGsxzcaL6JD0YxYg3VQfPq47QM8NZQxmrNmnMAYPz4NXBiqoJhLeKvxDRifiu
17rbJ8dxB0NuoLH3btS7ImubYW9mbaAZcSijdF8oKbn8KjZ2/+a3OOpiPycV2lPo
KG2Fk237I1YxewUogCMzk3S1p7sjYWO0hkw+Y9LwjWEL2Yg1E3n6dmRtDZYswRTd
KmLlGxLv2/yPOMnTceXHo+OCVbWLT3UhlCFRLHk/edUJCFTgaSQHJQzrgrEexoCK
p6Yi86bflmAxHsxeKzxHx1yIwWGRd68d4ClmDa99W/MfI1p/o+s3WQkpdcNfCP8j
9QQf3ra7kfDpQGbh0jiaF77a1mkaQH0u46fqrODRCDOElaXjVrJdI8QL87ICox38
rbmaCC0V/NrUm1qEYn0hpFX1Sxlr/iVksubAoyvkxdWOBKaKKT2kvUEgN+rVJPfG
hCorkufVR9esn2V5peoS7kqjNHGglgADhLma1S+gtRNpU0nzZq4CbgKlUMwlLEQb
/rNuWZ30HW+ejOdMIx9oBL/wWQj26YmCwrvUvC2/LY6TuncqHWidffI+KXMnC+pq
2wwwk6ALZuTsBR8SQgg89jxIEhvf4nZk98UziE7D7U9QPH7kwxa4Ced9siwCywkX
h3PCs//pf05dNa92Y0e9SPfl21Ugchm11U+cv4EfpGMwO3fsTROR8r55Rek6qCBB
MeEOmH8luMkoKM6LN3sg9jsr6yiQOUj/sWkTWEVP3SWxncZfyE3Kl/VD42AympZJ
mhPGkf0HcS0MWZ+q0mgU0/f6GD0s2nzF1FhkP77uOuEy9r0TzkjVLu4qVBGF7uxm
RJHPNmzxJaA2FukqwrWt/JDiJPlxE4lLfByKrJtXE16r3GdOflnoBnUUhPYh6hxy
jDRTWn5c4PVKcGIfoNoW0kc3IZ5e7s70oo/MgNdCuS6V8XtKhi0qusRT2U3QsqyD
RTgSluYB44pwE1XT/3twtccpLOOE6NKB58AtZrkwq8a8l/Uga0d2lKwkTP/Vw+DM
oWNW1g/qKkJRTBNdi8RvquIcuPXDE+hquwAv/abBVhul9LXA+cWwuinb3Q56xaSh
12CRP0E40l6Z8B4hZnJcTVz5T2zknkqXychG3j6FAL5nI8axMWOhqDern7D3FJYN
BDNa73ZZwgnGXAZ3hGMzU95Ev3BHUSw5PDEGGGIxWamPuS5Btud3bOMNrBYUWxWt
0Vs0fQNNuh64DhhWcuZ5TfJBey1F3r4WbpPsb8P12q4HXfo1BGfgNMbz0VHpPmLC
xFq1ykjuGYezfVlmA66b+vUD+rrjCmVUZ8AttkyD4VzblqZvg2ad+kNiEEWwn3SX
160o1OvSsCUIB2bD8v+TE4YcnR9/Z6FUuUlo+dz8s4x3dm8i6qiB7Pa9kyCB38r2
tKbTgEsXbLEnJuyyGWN8RNNa8OAQaVdO8s5Cr5IZ2m3BMsOE1XApYGhh9BHMwPxU
PbWehSoHtzdfJPGD1nWlDuQlDkfGZADCgIwN4IBzbMx9JzTsFMEua2q/sDpge7Cr
P1sj5McJCf6iGzq+MATQ4K+5oNehwQJZqjKv1TMptzfqxGLOJEFaGM5gyuKUjf6F
+t5OI1iKZyr302TKv52uNRSKb9HVQComzC4jdeLIChR5NUy02p9oTo18ePcCpOgn
fYIZt9GIjFMrOyQRhIGWUbApaUcrAMQ0ITt1A674fqFhs1tNjDTtt0JBnPtfFSuR
EsJCsq40nDLlfxdgnYC3POChqapiA7qwPBxbagst2+jLDi7nQ/++grEhB+AcLKeR
b96wPhGQNYZd3YjfBGLv6DdoHBYh9QuagJ1i/zF1FOEz7QZCTYLx09aiH/v0kLsy
q0TI5HlQrIoQoP0LEhqa3gyVOIwYHt8RLZRqM/+VLixA9Bzy0NTOT880l1xIJItz
gplOu+u72Oh+hdPHRmDVPL9gqkDKYVmO3EbT+EqAJxVoKEKv4ROm4lSTt/alND/o
Wm5OVYXNHcYFizB1Sq4z/dOgfYChMFsdM++ObCyD+96esufbfgdaRXMTa0zRkU0d
ALzAb9FBVaoYU6iMT51g7JbY+P2gS5Q9nNIKFKRxgDlRAYmFxAgmHoswlwR66SXg
y4NcSEc09Six+psmI7msRS1VPFWWk75EJAACJAQxKxuJjw/ABqlSgdZ8h6T2pwOp
XJWjs9qfaefQF8DN18RXlWnTd/qFozfg4G+0z5h953zx5T4HMuE/Lk9KwRq15FTN
LeGsei3MZO+w5JGx+JHTzgc5L6LBUCOB5fndQbRPfhPNpQNPmIb7QwORTKJFlU6e
hJ4Kw61cnCdqZpg0xsq72YVfav/0cZt6KzrsruWfe7cRUl51FmAq6V6C4TWWK9o3
xloMIILqdWaqJfE2yVUyKk6g2cW3Qkc3T8rGotsVgZB2wlLpxSPv+Di6e6kz3Eqa
Q+cXuTqXIURKdrqA+m3taxFzp2cPUgFzwbjrL0JB/LnvRtRYpqVxggcMj2nv2U7u
Id4pgEg3MQ4iH0D2K+8DVxgai5syZlzb/5GT6Cg3qofxB/pJoBm4Bp1V5Y3fNB1z
hrAzQq1CegOPOgJG8efrIK+ijqGMM0cif77jLUEQYTsb7PiCwdDMt98xHRF6MjMR
u8rh49ujntwSORDgHD3+GwgFK2Wny87AfKcm9Sa94hFoAvrGvo7vTEr4wjc+wghX
4/8OvqDKfTWAS/R+Zcd/VscSJty6IbwQnYvaofmlpOUHxoO3cbzWq6lgrr+2Hw23
q7xNAXTHcmEu0mstQaiY4boBpl5naiV82Zf3kvFbCe3hLX8NF9rJUoNtjrU+gVQh
BBYA5GoXVOsl2ZLQem3qpAVDEYZsOGgd4ZMIxdT0+ZGlfvryHoRCDyu1csfYMi4d
sL1v+2mye5KpoAWRQeZAk1vxzMElZ73lT0MOOHKrTk17cCO+7OQMRQaqf3GVMBKb
3iW7nOSgPI9EYeCN9NAA5VA5W/EtRPzKANVxYjw9yJA=
`protect end_protected