`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzTtbmj88bRWloRpjb4smh5r4RfvLurbzyuZf5CggY4zD
dk9VKzlIcpENysjdUzlqd9cO1SGlXlZOcOis0YZGEwymj0aD44pVKNI4xPiC1MJf
a8rdXRtjnPf9j7Hez3aJ1/JdT/4jrX72C8Vtz8QitTkSPbKJxktLMBSlmEnKtOkX
fv5gxMMdfTm+u46VLGPvLGw0R1vi6/Kq2xsWZWi6I1btVjO58OZz+Af2OqelAYC+
F6OCr3acYiNLFanBU4O3MpkjpqqXMGoNNEE0z680OY5eN0HqNaI8M7l0pKeEmjOI
K1r2j7X83k4152q0+NzrliUR6TqqSdxKBNUOYVSEWWaIWfrDq3gfnvAYpz6Ynt97
cthfQeSuhfDHf+gokvI7v0JzjJYHHLQEcIh4Pnbt4M70jYz8kUp2UyxpN2IB880h
IjMPPdMiTEK4Be7V/7KJIwHCHpS+xWsWYt2JdBP/T+9RRG19cTJ+gqsouk/Hlk1i
fUNqLRdB8DvI0dZJlqUbMi6dbJDm6SF82/DHdQPnobjJX+ednGhc+tuRFFwSx+Ep
jfEftwoPVq45Y+bqYBVCFNj7ou77T3fy41LJdrZ3SP52za7XFkaaB5R32qJLy0ta
kyvSBC9uykCgQzt0wlaFVyeXZ6NvSrNxpkdFMFgrmRMCrMHd9GTg/C6uaC3MASlV
KU/cqGNGHpnTY5LRNRX8KN+eguKlbiIqC7q6h1UetbEQfrHZWmzQi/Gmp91M0bkg
7afIL2dZlg9ok68KVnSUN42mI/QrsTjYxzS+V67U8XfxDIB/qs6GlBmmTDYXHxLK
APldeOSvFiIASlGWr7KEgDjlZL3DZpt9/vswhm47469Pdzcds60dfTj5ZTuqwcaZ
sGTTgda5StUTlc0rUtRsD8ih2hjLKgg/kNdUF0WIY8to9ScDJFckShqnd99OeI8z
I/JGYgiJYGHbASnvjoTVTkWGdCpxHLohjsqQoyFeh/xL0wLSIHbp4pNMcYDBPh7V
47mTNDHj3S+FmXboCnDWXGExRdyrEhahCt1DePPpWrm5MXCDVhR6SeOqA4yqAKc0
IwB53RTE2oArAJefWOb+cyaPLagmmTEtjNDbl3KpEHm/7hImiTDk18DzWIx4b3CP
0l09ht0Qjn1jzmragFuMUVQZa+ybzab/RV5oF/7SQ0DBsR+xALo1SNRHXt0k/SMk
LXyrLqkhAqSclwCoRMLNYxWWNwB5S9ME9NUyAgAu3lM5VJci1HCh3fT1901JawPg
4xTCalRlB2AsIoOOFyV3yXgr6DCi6iGhXtM4pzRoD1zgdtLGaRWuAv1s0JvKBBxU
7UMNHJRJ9zhO7EP95WHcc8WaXuA358hpxwOptomDEyPUlc0BWFQtNifEplEa29HS
cb+YK/LQc5w/VtTJm2PjxRwF6UHemC1GmGjwhrCjBbdAcJsgI4QS1l/PFxQy6H3k
qAA5bmJX6tmAXPWdwWSmBPXBNq1FzQqUerdKpbB+AnwpO1K+Ivy/7HJiLIMUs9qQ
fLZTtySP1jEHybgKFR2VS3OmPJJNXrTToyGu6hwgibMq0QB1LcCLOkGAlqzGehe5
Max6rfaLvnbpI4lk2cULL8UWxHLlqYYofU7xsBjekhzbxG7XnJ+4Zlv5uQInYcZA
/RcFxEWySoqcxEwZKDhObVe3DbvrR+T7iMR4odzkYIAb99DKuNsQ48SmZrC4rlss
MVWsOA8cUWo1QEYXGr3utpMLU4PZdEWgBqPhzR8KKZvdlG23j+hNU/h8qm0RFilR
Nv7pcwVHG9zSnHuAMZS++97CML3TwQQQ/y1FwcYPm8u7J/Sz3ZCePyVI6fEdalGk
2am3PDk6my2Qg8zEwQHSxQF9hstgm+EL9XWlaSXi9IxWTJ7pG/fJREe5XhR2VMbh
Tx/+0DLhNvZfevg6HKZMxQ1QRZF2Pwa0WNW168BkFQOXRdf6tUCKf7cbDs/ZBjIT
c3+k1Ct+eTdj/yfOtn+RIIOy+1wgrTAG8Ogsi5xSTJB0+1BqHYqq9/5P7fNzjsWl
wYhw0V55//wnwvJYbYjnoztxsp+nR+ZkaGtdgHO2pF7KonyftyHYPONQTEmoe3tq
5jAL9XQCptEd9VtB9HGzzIouR8fPPBaWU8fVANF7sdX/uwV5FuRRVDZPnsMLkNeW
hrULyhzKQTh+ETlXVwRW18VuZnW5OU1S/hTtQWZn0/8d8A6ZfB2ng2ScpvQPiB5g
GSGvtZQ7dwyBDelmLjaesd+7AfnBDfeU/pXlBXYsCErByVIjia4cTUborTyuOtz+
y3WbZPgnJM1VqBhT2cu04bHA1JxIEFDkRV7nvg9jOOJfIjgngGfXW/EubG+Sz3ps
SfP1U1vIPkIiXznzvzWDqg1CDEVsa8IpKLqc4qWTxMoTzpcL0VxvnZRwXiL9Uz48
jv/YUNDwdiS88iHPx2HVVZKKqWf7jnpgGvRbhrFReXaHf9SHDyyRSbR4swf05lbL
iM9DQ+YOxT+YgFk8jxfp3B42BiLeUJoolZMWVZ0oc0Ve54HSrrpxfLS0d0ZVmg+Q
Eu98zvYEAD0R9mzfpSPbEe/cG+JFKz0YJ2n6J5SeyQXTAAbjtPpfP4YUYx/rGw8I
3Aa7xKg5avSpMucyhPzI52FZ/Guldv9iqsFNsJEvDBUXdn7NgroXE/JnmlgKGxHY
DofggIVCTWAyIl7TyVIliMadROD1FA/cM/G3JS62QAsYVFmYSTTfMWMtEcM/kvT6
0b2ZgS0AGz/2GQRZ6vdqDUbAgmAS4AN6GPfU5Dxz5loqoVU8xPSHdfR4g6zCXada
WGqgBAniJDU8t0gDulaO94MN7+8V5FwfcrFs7CwNuNTnFEwC496Xvvqx7jwxLbaZ
SSEXnwcVQ5ZTJih5GzAGc48MLXV1kkMdPTb3V9V8PZhCVVQnpt5saBduIFlGQAVt
Wmkn2Evkwq5bSMtQkmVzeFmnh83WMJKr5vx2pYIPn9S0n588jZwydtQpT6gBnmHG
d3Dmyun37TGqbMu/XY3r0Aq8cpnJ8ve7UF6EtVTNBR0xVtuUPrw2+yNAtoHbgS+X
U06PNu1YICnVRqaoVNffoyuczu3Ar2AjMYNH6t7RNk3+WjO1fyCQsj6sBtempZYy
GMBbwmkSbc3rUK9JQ6tf8F/VL5O2qppK9N43o+wPvBqjzo26FAGYIanh+CvYHERC
tFA4nfkXgCmCMeHjCAZroUJrJRHgOz6fjwhzqmfiInAmcpe13P7yLtIKI3LksHtv
oxMrClIeJZ1eLN4GOZWR81OuGKsTpuOUkx0RSmL/dFqRVoUS/u2GShxHd0tYSCV2
kFGxskmL4WMkDbogdjGWvPKZ9i1X1EOxBQlr0tSqFLZ5lP9jQTmQnbHnxyK/xH0Z
Wqi86z1jolDQtP55OOJBswD+fj64qoDzQRX86FqagGJDj+Irr1A4CzYIu/yryjW/
/cyEOs1uzlPYEo3NBnRDEyjOD8zeQUQ6jTm4ApoRKHTfGjPL9W8UM4iiYoIaKlql
On2HyA14OlNETUfDfxd4OSCV5TbvWvmuduQMegvkYwLJOl6uZ4CsB4b78hC1ikjG
GWUFHwhUO/asCtYtOe8sqjn/+pRXbRfFo4t7fz1tdFIHAmrYN9mMZNGADFpL9kRT
KBHLwb9j6rni5BWek2qh0OyMzN2wBMylso9jBQo/4hryexYwLquRi+mxufcI2Xh0
6GXgO2gL2iXrEB26qq4UZPy0xf/El+GXSRzWzSY8igZyNzAH7aDKCi5N39XvNoy1
SFfsOqSRO1lIO/+56CVa2f7hN28Zg1HYAO5qYrDhWtP1o8IdPnEAuQqmfHJTX+/+
Ucqt9XTwZ+FLkYTNVzlQzoUNegcM4AdswxB4fjt5Ck9WFjatd/wbXI3gzO60rTLR
tvPRpyppbtSamXnXTKBsNrndWZ9aCCXw/SgKI8c6WD1I3+bqR9hoEAu2g86IRO8o
xXWfBUG9feEGa0tve5b5uN8JUY86izrKwhiLaknK73gpsnjRCRCIvCUB3RXTLj4D
J+P7Zu1XCb85cjze1hBYeU1sGoNlx+YWqLJPSIXXbMlZPBlPMRd8Z3E/1d7sXBij
buCIkqRGSsMwoRenJmDkVekBPL/OcS2eBq7522XXxxWvu0yeBOBz+OAiQQgs5+ZV
7S5ri7O5VWmZR+rFd/B6cKpcyH2CiJ/modnjC1g2ip+K4YsHxrELlFvTSeLoTUXo
lVAU69dyZqyV1a2UwWm3k4CQMaeMwivayH0KKHgroUzxHOWryohKU/Q6R/GGER1+
xtvt7TOIW3isTzb8ygdgo/i6/d+2BSwOmY95tiCun49dGhGr9peCMIfE8zreMMhg
+04C58tDFoFAtXO/gLZz0hU1TZqLLBY8SVAJgCEft2ETBnzxLOdh64JhTsG8efM7
gEhdq+saY29L5ZMcTRGvCW2G8KF8Tc6I46Y17W0t6uD9geupNcknebH2N0vY/wKq
qcf3CRI4qwn4GyZPz2tP45Mhk/DWJz84dm3kno+R1Z6VK7SQWjG5MRljz3hoJaOO
27rxZgtzkqVKEXhh11hkimfVQUskkJfP3M9H1/6jQDyJ331YKB1qKLO349TY1pYa
3h04KpsrOe2YQzXkuqw9rOkZVi0U+xAk2EneOVvzRcObabpEN8yE+Zl/EsRO2WUD
8nWtvaQOPlhczeAkzEonOIeIk1htk3RHGbF2kHiPjPF0TK8m+1sYyYacmUh+3jqB
NDk6oRV360nq4+e9HjDjzmjPmbKEeWST9qNUE2ABHKUCRE/nkEN3UuysQKJyHXj7
qcM44G80nORAQ0o4dbrV4UlMJj2HsVblpStHC1l0NvCf5wBPTWVGndN8Au0cS/gE
BEuY1L7hltjD2dVcyHQxwDLm13JRTh0fY0z/NXe+DE7qr69OamVPLhen8v7rKvP+
AazUjf+mhEfcvfvDB/6lTx0us7EVRBobgTLJNlh+ShR0e3/q701S5D6NZCCAXRH6
UZXPnBxsztOYfJN+AipQTkh2/2bthLlkL+8J1uANrtMnswZOceTmRPGZde3hh22i
yQP1ImvG++q3KzMj8LBaZovjyOZBP8CHdYgN7owLWecS847ENFd+DIzr6WnVgKGb
1VoMtGlR0+EgY1vyBqQ68Pcy89lLUbM2ulNyMhow8LLpyoFfbS3G/6bssrmE+U88
oL3dOVhrlB/BMUqsHFmuAgWRIQNva3HrXRt/VJHdK+Kk3v6nEwPD0qUWLJr+bnXK
MdKBP2aa76Zn4VcQom2SxaHzEiBlRtdvyzLdvDVKgadharrdbWDhrZIX2Afp0+V+
N87IURIR4JkNUPQQ5LktxYjOVhJ4ueLPnGZEGNP65L85yHM50ZPnqZB3C61FBYDF
i+f9efNBj1txwCdrDNdYpI5+Q1tIgTeJ0CGOSvmhkyTsdKQi/o/mMXAFXKxCow15
1zRvX2Md2dJLyWa0eBPLSq5ODGwWMiVu+8G59SA0+2H/eWMchOsUK6dlwz1DKOIV
Ns5R95rrOwl8E5x8yflZqnLiMUCVaj3dl/Q599bUi9aH5zZb62MD62+PinT1DhwD
tAvCd+JBo+yWO2RIEK2Js7TjfpLZLupVG/V2DajUBy0Y/A2a6WVNQcoYkr9Jn5V8
rSaREIfp0v1D7FxWYiEkFr1XM4Ra77kMTw66ARro1hxlP4mw/9n83KQpCAimXI6u
Rp11emYjKs9qbNDqvQeRvc+munlYv8SYLKb2nJ+Tq73FqFDGA3m6rFulg3nQX8B7
uQtcLFEaW69PrHM2p5osY3E60EQ0bXP77h2CGmBaN6EJRfiObD4qaGf3pD5fugYb
VruHU+QLZDN6DYk0RwNyPDWiQbHuB3KM5R23t+3t2s8KWjnFkkxBLC6jSgpIyJH9
njLyIEbbvz3m6UlYyfwKP+fkySLODoK2qlve3RgyoXzwLSrdmTvfOm7hyp9kCPtQ
5tMI47ewl9oWFlDvzFKfYl05u+fvQ3Z9KETvf4wQnSfFQF56i74JgG2HVCBkCBEH
Bjq9WGgrTIZrmyDESoNzztsb4Bupn7lsqzpJJNGTHa1Z4RhKOihaF6a3F4HJ9Zdc
CpcpcZlTQBuie94S4TCmylbYwluqvuDzdwrOI2IZECQihkZEqyR2/ngyMDeSQ/xI
e7k7HjzJsAwRD+AlRuWHutuVSAFN/DC+4EGo4FAFgZnZ25ETDwgFE6Gge9AyE0hM
EfnOUK+qQd+Qp1YXz5TbHVIRGVyCEOYVW9L5EuSuGVtIEFV3GlnOvAROhleoG2W2
Jjw2IDgTOqu4B162RNkzl1QfAapJ3bW7sBNi0QIaflgJtx2C8CZkziz/i4su4P7Y
rNKZaf3PJsVCAUkF8rK1dAR4HiPMxzOWJjSwWqyN52AkLgqXLqQ3DgGjknK2cIQh
XUpMbUIklOuAwnKzbRMLiSyebaUDYfZ4kBpjA8wqsCqJ0yfg9LXts/bvvA9GWUdw
vKeZ8jfkqChobBpn1G0lEiNhVZ+bv2tVr72BkwLuO4tglphLwnyo9+V2XJWJGW5x
XH7l/5uW3JxdOttcGE8XhihXbyoiH3vw456jURp63YA/MFmIrIDpWRTcGQc76p/n
ZU+c4uLmoa6GXpQj99XlO+02hrZxfxWpBBM/qKFCpgMFyJL9XPMuVFDFovsnV+uk
DYAWvvWQYhinxBFj5GR4e7DHGryHCwyZm7g2j1+uxVns+gSvhJd81Iu04/hLb+HZ
B5wUmEh6YDY/G2IQsR9o9dNjsOeOQjoffkHfQygxdzn7yD6aqoOCzmBqcxdv4VGm
46daBsJSy5mvqD0yGIfMaaco9LrZrdJbN53vRY2oY8ug9PGG+Fm+AUr618Abo55m
AYNs+UG1zLsVze0KriGyMEg6mjJCKOqv+2ZJ6C2nXKW7vsb/akVjZBUgXuW0Ywse
xjN1TMc7R6WL5pY4zxSuvmNw4Qe6cm0VleJil6Q6xbKnryWClWRpirz5RoChQzg9
yQ1Ti4tELkz6FVFGvWndH2MOdnsmED4zHoOYw7ayjQVUP+YHU2hbFW4dlNi0FshS
XGPc7qXfNnHX0h98ASC8rkgKQup4oRHpYytGIkh6hD/cNtYirgkrQ2a9kq+iVsjl
kPYk6rqrw+sa7HTIyaiYj9QJ1NVuaKn1AhMZl3HaTNYYuNrsM/agGDjAByi59+aL
QNYm1ansXSREI9PMBLliXQvUnbFRmiaSt+MA2PZP95OqU8EM6dBlPvnFXZIQu6Sh
8ek5/HVd789nFjshiuqSBymHEhKFZ1ghuyhrQ4wv787tJWgcmj9e6HHItcrQU5R2
PL3A+ExcB9suvu74L8Q0nl7zlELDoOTYISqXrtkCDtqtKhG0ngxmqFp/1mSZ8EHR
pQWtrg8KkF5f4rZum8lASC7FCZWDopkfxSkmx8IovQsyMgT72hzbuYAigziiAfyA
PhG4ItmnDsmf72YhcnvxKzhqmKCPoJo7Uw6DNgtJLbRUwUVk62T/GtA01SEsXXJR
Jow6656yfTYZ5atwoTWGhgbS7i1pHewj25auXW4H0ukFlQ6thECMq3gOvtDsARgX
pds78tsWJYW8Aam0xGuE95Avfrx0ER/tgvC3Wn+J/Os1JnVEpKgZnnhRPXh+FCZM
cPZu9xRhbWImLL813yy/2dTK4ON6gN17180nIkUkgAYhjbFIcYm+05p4KdvaiWfb
G/XEXQ7KaTCLdiqPsVKkdC9cnQgAhCSUHv/we6k2UDIIowZggqrJfNjQIKjTqVCa
AQxasrMrVDmiKU5PDtAyQvhnbLE8lIchAqU+oF7LddNmh578MMYsEOr9vQXvdsF4
w8sLm4xQsRJTUUPeS/6KyFqXpeq6lZt3vTK2enNm4AL6yFeXTZS6zb3iCxY5bWG5
WywVjj10p1ufx88qmM9Nt8QKKHMOjHA1pd+8Y2gB7VUHVAg0VzETQfOLyeZ+l1Mq
pt6RDLIfUNq2O+IqUWqhylOZT6MaOdekcJNlNLoZmPI9ZnoUH9EtUpYm3cVTIZqt
x5RreIwbyk8BxBOU+hYcCrp3NBiK3dZNqOulXUf9x9lRMuifPeKKBKe0laAyo/Hf
9UMGm/KnwhHh6TROIXmEY2naDuop0mrkRiepwvarow6bbE/4viLJ9v2Evmr93Ljq
k/9Ka8H+ULmtMeMbFyH0S9IBrXUixXgZ2DsGYLCarjleN1f6R7oqRDdtTLkZXTcC
M+Y5UQdyArNDnPnd/8aMwJ24RG/f4QjTtjEv/XeqxcQf9t1QR5safMWYsoGlGgQ/
c+aXUBZdIszlwLRvHYgCr6Yklv1T2pDHq2KXVo0K+D9DUlwSN6UHGqYfLl1LcD5H
Yq5sGEWhK9wh7NtG52v0TaJR8ukc/BkYqXw5vQPANShaIx+Y6CX4f2zawfw9pjtm
/XHquYAuJv6GCNDhMJoPz1u98o7OTcDcMuyQTtRAAPQUSfqNVY1zfa5D1iCe6nfs
a53sord9QrD6/ZOHlxzx1T4SD8Zyr6H/IhmRCU1ZAjI3XSlBJSv6coecqFK60mc5
knphHFayMVcGDLC7Svf+vd3fnfB6mwsH81Q61zhInh3qSEdm6DsH5llF7vb4f3J1
V+awLdxI3H9bECFCxOSsrU6pft0lViTsN78VE7UVBokk0yJBDaVOWQm+I+781gZO
ieHISBXcS8MIAsLXLjq17ws+CHZLmosfDkYew8MIe9oMGpQ4WoPS4RR6Y4cI8iO8
4JpPlaQanoEJq6SMb9BMqcKWFl3hh542fV2ZPVxJUhHRAjbfK8hdl+s8Ka6aJNfx
AnywzwhnQZ+bR72eKFbjpjZ/VZxwxEur41Tz3VnHo3smI0uyYopQfSoTxQP6p50r
w63MUo1WcfyqAlgL8jd6RNcT8HRWsgoDMvL/sF3oQQ2kiCx3JcuPyKiAss4Kdf4X
71Ox7xigq1TNy2HjhYMTCoqNEnjzm0wA2ahUTKonUf9hIQDxYvpEEGqspmfvohNt
VQw+tNHpR5CV0fBg15DyGmCOlyfc3CdpxvhFdRM7KolWUJQjsBSzdp0HJ2e4Mbme
3wNNwEgDL52DoLGIw0GbYBBgJ1VE9jXdAEEkB8Bl6G0jQniTBY+9i66FhvqaJKoS
Si50r4G2vHsAN4yPGwuWYTcT2xeFbQ6ceXesFjgp9DmIMeVf8BourNf8KzhmfA6N
f6DuOeNIUTG2cdea+qubzP7d3yrHjaSxhRy1ABJQVezBwRk0vQSlN91etI/BVNZn
5E1+PMs8eo8Tzozx2yy7zrA7W6I87zJ9r0s1F5Pz61sMrUCInrvbSlcutfHyfzp7
qmFZLXvBo+cWV7fOx/ODMG1bSehRqIOO2AfvBOfyGn4/h/LOpqoWlmSgo6ySRujT
PUVdj8mroU4GU992Ghx1gwufjVFpsQ1Qbm5pF7SLWymzRVqMd7Lap/w/TtZ65ZEL
/5wDwtgySRk/wYk6lsHXVfYV0HE2gS+NGrlpM7IYeWP58StnfmnpfkFJwMNMYwoN
dY+5FjVwfu8nAS7g9Ui16uwtpyqHteSoiEOj5emxkdsm779JSFllaqUJsY7g54mD
Q+VYh70oFAZByZVXq3+PL2Etq+oMAbWpQoI3rtLHGfgLDDmrhci0gse/wba98YWl
KLhtWFPtbmEgvntqKlxV2gzDjDVzMQDoS6trP8J7KKLor/cDeNAQbvd4vUkfMZkJ
urMREioRXZz27173s7YYLqalF6cR3n9HjdDSQrabVr/mAKdMwuF0LsOeC0qg9jSn
EACcSJfasdMxt8RXeSqeoaqpiOhc92YDoQYJEPln+W8aF/VE87FZ42bBcIvk+Mwr
+glTo47hecNW5yzwbQKdW0QebVngnR3RX3zLtL40PsFA+AyVPp79hlzZ4RnAS2uK
syyCM3XkmMpsrfkKhchzptNEjmAnmEf/apkV7iyVwMzoJkys0A8YE7/kNdjuVxiK
iHmN7rTJu5SW3EIXhfTn8Ivc64juD0ui5qDLcy3kRmFR4DV0dWzXudQD/Dtj3n5r
ar15CqqcBnJX76TzmcehQBBnGthRzvYdmi/T/rryYyU3eFN/2HOCKzdhIIYiIIsF
/eaJLNLKrvryTYCiMFgDWNipzrnnssrWd6JlXH0pai0o9pTvl4DQpmoQOR+IGcYb
47ddEq4U1f6Mv05M3hRhbBCuNKbqd7tiq5dMEQXuh9Mze8Cq+QtEfQgr94i7kqtw
l7lgeAI3JlwnhTUyld1gsW+jCr0J2q/nsQ0VLwdDdXBE4ZNuLTiBSA3GAd11aJY9
2BzlzxmYxqLKMMDqXpFMy8NQ5/LZIkqSacUVsw3stKIvGvT8TM1TnZylenTigW9h
Xlk4cq+TP3/acheACC3H6IpXKlmNZuLrba3rEtTb+CxtRINZ1/GXAiqR/vmMK+Y2
hi4DHxvG/ZBpEIpB5GUu5vIAip83rxA18wBMQDpSpUVmBu4kWuSaqUW/EWezcz+S
aWajngVDBg1Cy4DBHHlarO9Xju/9dheO3RoHEbU4BoM/FHtE7im3LgsZw8YqXA62
gxiC7bjonRp5HDOTblxdkYT6JOArc2g9W8/kKRF/4MDWNklxDE2dxf1iOK3cwy8a
jAZ+lqL3tstTSCaef1I+EwWUL77EcjcsooibUvBA1O5XSEMrgjDnrQiWpLe276tj
nwAwPsm/8lbnZFiTVnz72I6V1d7dAhmTDOmhPRlNxSAxpreRJxA84YvnuJG1kC6S
vivJtKOxtpv0XqRWl9XK5SPkSlcloh6LRCnjL9RDImTRl8qLYPLwa7J+XRfofOJE
zobn3hQR0wFYEkLTohnxdULbco3zgDSuS+H3lkmWN6Y5gKDbbZLsTcvD7WCDkRMA
UcSN1l4nB56sJHdT973AiqIOyvSC0MhuRMFnjFiP9pT1lNqPvWocWbC5C6SA9z5K
DPjyvPcvjEcdJPcHYHbbJjhW+KlY4m9d+/phlVDCFA6Yp08WB938ZDPA1vQugCNg
wtIvXnmTmf6/u1dZsq6n+Ju/0G/Fr36SJrPSJwQHo/Eq/gBKFV+UpdgD5kJ9VgIX
Sd/GxgpTCFPjvp5/mv3EBUxNWPHTyH11Udw72HWWT1jcx+a+E3zvaMfYi4GUVN3U
YrN2L3QjZyQkDCdVzfRdWQRWdFN+y06LELlxJ+xduE0V4dtt6DrMEkFiLRlMyW3d
J1iDyMZrOKegMeqHW4dHg9+rWMcwQGyb8+W4nGQbmYR9hQ/YJKGSk8U+PkwMMJv5
o9Fjm7AdRjzTE5riJzDDQskwup9JToMcBK0rDm4oypmb7BLURe3Qc96+z+p9jlZE
SDH0UdkaHlwPQnZEjHMh2iD/TOclNUC6QHdUjJfZv5ywIbz1U2iCsSEFfgrkLP4U
KuYHWXVegFgrNzJkbjxQ4N7E7HwukW1qEKhq5o4PXp6Gz5/7ujQJ6+6ggIlCO72a
kZvjvbtLusHipfJ57efTHJdgSLMSRuWn6j8Psk6nN+7iqw1ANjtEHEtbgHHarBgT
uj0QxAqMfMidl8mad7NaXu1X2JtunjLo+pc1QwL66eOCEIPmdtHELxDLDu7yA+t/
msutXn2GjI0rhiXbrbkOFS1GatCavUBUvqMZu0aQJx04nvKXnG0u2yoTdjhzkk2t
htc1ZJIS5xRvlgcYQX/+gCJ5Vs1IkB7z4+tOjdhVR6CpxMLBS5Y9SfcRwD1OPDBT
cOfEa+dhwRFoylPANPOn6qNSask/1JbRHF7gdktJbvwiw29GRDlWvVNmjc9IDjXf
TFKGQg+0RwtagBLr29PlAKqployvd0PfMYnSuqc0oZRBBuP4kuxvxlX3+jVJj5yJ
u59N+cgOeluM1bL47WUbCcvnpDUMe1iUAHE4/ZDMhddsiZJzFmHD16dZP5X8f3vy
f0o6//3hdFKUVPK6NGX3tBiFxv8WJp7UlM2jsvtdEbLDrn9vyfl7BeUXrV/YcaTO
G/ee7IQV+3HH6xs3Qnws68N+712Wvq6C/bKzKQ35pQ3eRRwEuK/MdIZ2CRRmDJr8
wCFX0excvznbx7264OVNdZ5cl8jQVMeEx/TaRSSYnoqvGjeYySYDf5iup4Us3LmQ
gO014w0nwcSCVjc5XTcOIIpYoVEqgc8C66gVAcyuLVkCESjJWkdmR5t/IgnLtQDG
LEVKo1NHDLBMYtO604ozWBwr3dgX4tdHqLF603UVM7+fXuhdTwefvvkCFt1QOhSq
F2qtHCn5JQwRVKTiKClNyL5EwDz3+ztqe3lqyr7qF7uVyuzNeGlLootMZJIgdpmF
NTzSHdjjnYwDFP1Tbj1nrlr6RYw+gs4DA04y0Oi9Nthu1LFrXxkKSXF39eDkkgXs
rWFu8oFYmev09SvU5k9gRT2L4bvw3o58ymyV7XsjP5M5KioorrkovIZfFwHJYdFG
s1h92TYU0499F9b1uT2tiWJpBcybE1cUynL318b3DGvS3k04N1MLXtaL44pK08gq
wIsD+CBMyWW/yVqxEf4QLQM5KpCkpB8F2CSJmh6LqDwOjFN01z/3Z4aR9J8kV/Sk
1+eB9QxICT7PVyAPsbBB8hn0wJjMqLMCCfRdtqLKNVOX8ad067lTHhkRb5wH6bl6
g57PE8iz5EP3og3FI9t3KlKr4z+Jok4Es3fi/8RFgcjYL55DBcRqQpK/b0/qY3LA
SEXxelc3Q7hGPMMast9L7D/y4RalUajDo+JnI5MmG0nD2Z3kbH5UhuVQ/KiTk9wF
kkf1JnTpm4O60kM7MnltVAG2+bZC9Xl4gpXCT+kuIolha8X7/614ye0R1Ar6E4qi
aYYPVwVXVfennl+evm3JLND9Eoywtxx3gxvEuoI/lce5iop9ZiW7vsX7LDb5ukcw
i8H0FJLZtvdfLnhypihG/bhlrct/NOuZ8cOsXUI2llyFdmqSXop47hcr3nMQ2tBe
DExCcSEOjMETzPJLLedggxBPLrKNlEf2Q4IivoWb+2Tqq540aZx+dieqjn9hU1nn
CyoC6qjKCb3ND1IyC/w8+r0bUkS3qtV0b/eZ3Gq0yMs4J5UW203XqB1Sb4T16knL
1h2TVHrsBl/3H4IPjgsjQtGLd6oq/ZMj54A64XkBoaxWJwMyth6C+1/RFNe3jNiN
6TJOE2ITqmGkAbqu3uA6q9Pnl8lhftlGx6L311BJGUJyygns89gGG95KsJe3eezU
8eGeRiVNIhkuEOnUlgDMudFEha9NP/JVO+8jjQob1Gk2WEcgcYEX7HgMqLnR8m4L
XDnCRo/7XJ+5AJgwZdQTWXA/5bUbfgXn+IGfGPpxncEwuu3yJbnRpBVlI3dvbNDv
z3nRacXGijUyZgREDhjzyD4HMq8C55UXvAXPV/8y/hnI3Vlw74XmZDqLeM6oz/rp
JxInTVDvwoENAbbXTE53gbksRkzqa+Kza/3UROv7nOxyii87uftTAp7QQjpze+e8
TEva3Bwb9nJLrOG5JBjr5MP1v21cXm9JFJ7k9G4AC3HgOgcOCsuVMk+XAZdue4gz
CY5vcbVCSdoJ7pzbOxnXnDintz5VbqbOjsDjokrwqk9e6Z/uYUMPk5vziV3EfFRy
w0FY5iSu1HGOYZTyt7drTbTobYCGnRyDej4CMweh/trx7ObJ6e8x3I+k6Gx02bUy
OInaGv56yUwyU+bsavzVAhirIQNvUnSTqARDP+LP8v/nBy6nWxJfgXQrcP4Lmz33
EMoYqGZ/RpNPKmx34TRKmiuSordUlCUMokGG+4cr+hMDQxu2bNckEmE+J/ZrLjpq
+B6UE6UApFbAFFx6Xth99/89vP1yUf0AzxRDhlI0QnDtlr2VFshkmk2raXZk1CY8
R5eqwiiA+VeBsoL9c5OEp2fd2ZoAuq5HwgD+INC3ip/bHvjC/rzTiESlGP7qF/MH
C22iQgXdQyDpzKoXSFFY4W0a3YkP5DUvQuH1bXaCL4Zpl9oD5BjwjZGUkwWhLsNG
diyocTKDQiQAQUkkVibndtp/urqQxcy3cVEoFW0OjPIQceSKApLC+1HC/s2JwNgT
FpThCYgPIo4/tFrr2FnZi7TO0D1cO3sM6hQYRVWtf3MQ7qBOjcAXe5Gdn16tUiCh
p2SIEZ/OW0QKx/KP5oyLKHjsOn2eW0Q8oXvuYPy4hy576Iv+OFJy/VbXTDgemkWm
K2BSfYHYwoRO/eCVeYI2QUzBcZsVjzUxwEyDKkH2cHaCfqouTD+1hBzA5YdIi9fj
vD+1iOIpkjBrxF4Kx2X/czYH0LNtS3b9PZ5V/YkErzPA2obWD3IaWwY3bTSMDU2C
w6HbhXLl+EdXNi3QD8Ou3cuFr3f6DwLE1X8t8EODkzzSdyFDuiosHiON32aYPCp8
a4yS1FY7LggeSQd/Q+68yZg2b8Gd7+VKf7HYJ6FA++QysC9PrMBRRb7KopN3wjpj
9Vzn8OEBXvxB69kNNPrlZTzEBC8xKPSWy3Wm1fDy6+qd6csjI1fCiMGGQ5WBpany
hlBlrUhpn4KzRdyGCjG1aHJ3WPCJcoiag3cYO4/wGHgfgqzKwbhJbUaDSLwgY33E
6IxxGglCZnpG6TMvyfpr97gOf5dnB0bwcvsM5VsoFmsnsZK/pXMr7asJIM+qlKwq
jQu5ghoXTfAhtSrUnne6KGGc4ngjo07dNkZoPQQASrHq+JAiSQEeN0yzod+/l0Uf
siMeSHvma/cIlyMEp6gzLx2GQ7vsXr+nf50pAbUWjIwX6P4fC2QE5CEPzOGbwctN
0GT28cwe/AFPRuyQ66T5hfq6fokbTR3SjdTUttGbKm5w+Kb8zOU0v+IpK0/UTARo
psthSLQyMUISN0FaFwKVe+y71o2TN+CJ0Yn6giyynNfqFkK0gzG+S9gr2gll4xNQ
ji9SpQgvxNeGBiBb8LA0MyKl4ZQNqITfD2Ad4Bd8nsOpWXgD/F1Z3utlydb50Lal
XQxQ/yS8kg9/30W+vcdF6HwQbZaZa4RCrZhybSwwYETLKljjv/A811i4vis33CRA
pdTcCrnuZQ2aNpz4nVNJuhbIcUYcfmQRkNI8vVb45SW4PNHBSRqTE5f9wG1dbAr0
/vFEeH8UeI93pPxKFlqd1bawU5nt/L3yLkE+GxBa2GTZ7DhPY4ht82Yrtv8rCR/B
TKIFR2eepmpqZnv/An2f4e9t0uvDcxgFRauJsyyoY0+8qAad/mahN8xvyLE77CJi
z6aEzuBK2oKmFNsAn2oDn6lt9RJoJ4zcqJYSz1GqQfWwxdmDVh5o6I3MU7Z2bOMp
7jnGhmPmWzCJAK6XF6uA55n6kr5NzK5ffS90FgTtjBC67lVO7ddzN9qTstYjqOab
EXIuv8CxKzjkqe99v81Iw/Q0wFWwdI2UEUwMS42fiiZLjNo63y/PhhTmhZ64ZpOX
XG0eo0DBnmUjRBxzp+jG91dwCDWBGZJkjms307UVUh0/q2YBp8Rrho87pZ4/favK
JUusqhZoRLWaHYPDXS4JZBJFKwHkOZEuAVy3XKqBkG4chXhWyPAR62oRJmqX5cg8
ah85mzPVP9bWqU/NiltqXP5/WthkJeRWV/jNpnLyd71R6b1Cde5m9xV6/YIHKRqo
OcLxSqOk8AGq8eWO6KykKOWBR4zzNfNoBceBGzkRBasNEP9Sbd5n5U/QwaYYHTJU
1/WFhSyPB1U/6tSLipZTjLvClDIRCBNHeYun0Cfpp8huZgHKBfdIz1oowmXjWNJ3
UYjStCkhime/ltqrmkDQskL6Mwr9h05zrj1X29lvlm3/Hk5BboiUJmdLMdqgvIzG
kyl1aTd8Z4oSfhoIy+ibXJTnoKgbxvgeyd4MaHd+hlxqa3WExxlOQLwuaeHyTzbe
pLdyhlyG8q6Zp7qhroeeDqpjncnx2l4UcvgND6O/61L3kvCm/HKCjDv5pZLqEyVU
LUyM+4RsWwWF1Xs3+Rv2ysV7RfhAWfnSK87a4T97lo10Chbka7h/CUcA/JQRbVrR
95TbC0CeZ727nFjgeQN19o8MIHLaNONso7/QS5P6h+n65/nLzaSZS37jENTB7XEW
e1GNk2q8o685VScFJTw1l0GYD0GiT9RnRU/oUFln7yVcSYF6xUHLttpAnwCe3FW9
DBlLsgSxDJ+9eY10/HOhbAoIuGlu9LfKMZlIene5z4QopJwldfEW/FX1jkheQPv+
iE/F9/DGF2+80Ic2cMD96Mt8lQ1IYlKdxNHTtjd13CNJcQR1UnSRiG8u3zzxo3hW
HVV08Y+U7sBRtjUzz5qkLPpscP69YCqdwAGKb7H/7O1KJbnTzKR4HhcoAxViA5rR
g65FDXVITr1ma1MSISe8jDmkhakYyDz026BrSg36ZrCb/SKOsTNWxG4r1mdyWQ/M
bIxwuqGaMC47kUBQAADI7SBrNqpBrdCV+Xi06/5NLF3/IFNUP8yW+s0wVmzkKhvO
Vg3AH4I+pVbJpuXypLJMoF3pFkaN8hWAwyNH1AsLkcU+ybQH06Kk5VkiGJCmxjKr
iRu53x3F8nYdgfkFJ11bUQf2extvRqyDQfTb6HtZgUmasNp2Y66xPMNjPW3JUggC
PafV6soOAN99qBJQj1dX09oSC9+SEewVzAc3o8p8zxVt0axrWy9ayTvpkRWX+Fya
TeGFMj8GJsGMQUwG96mdYbJBU0c/khTjbTBZuMGt11ovVOSX/qGlQDIdKZNYy3R4
v45x2/pmHX9bZnRvHAuiwagVpk30Wiuq3NfuNOgWmqHPbN6m2jewFVdkRHuFLxfI
sYzi/MtXNZO8GHOJlIcicl48Z3TztRzXjn+8esl4ZiGaqROkQA0CrfWMlXCPD8A6
oH92Pd5suqG/MEh09eQWtzdCoMP700Ihn0n2T7UQx/DNapSNRy9lmpOjFcM+X243
pQKZqo/kF24Irqo1KI77CWdowtK3ULoWd5p1GTG+8/cJCNiDOLZZL00VV1YbMJjv
a9cYVCmq8iOXhI0ywZm9frFLvl2yKH2d7sFMK5xd5qJ6K5aDh2QUALtRAqiPspZK
EHPd1JBPGZQQkNJRljcPOML3Vtfz27xWZ5LVEy0K6uoUtmv9FFysZ44R85GajfHj
u97GxAjo1HtrUtQPMkhqNmt+3Cm8leozza7M8ICXBZGk2Z5a1bqVK4wE5N2rhi9f
rGwheUBSZOYJtODMIyHVY0UinV3WfZglbjAFv8fo8usUH5D18waolDaLASauyxKl
7DtgDR8CAMQPHSsgbOmBQ9BvFqAtpaaakA737IzC7WYe1I5C7rOoOt1pNJuV0TSE
aWGgiPcW16qs9n4dgM3ta+pxQk9949cnf6+tvy0leaSG3DxwjJOW85iPOpVQhSi2
i1Pth9CVxMt9caT1v0IOhsBah40VibdGZrmLTSSmXXYbsyPdgEXnumc/xUaB8/BV
yuiciDUFEtbAL1cvNc3thxcs192SOi02vWb9ssirBHZ4/V4/Mv0oR61B8o9i8tU1
AZy5dG05hQoJA8hpdNWZjkJ9f73bURgKXUHSipVnIrpxef9BUhweY/nqINW5trud
BFdw3BAretUd92c8DHANblPNKUTXf8JhXGtbzY1TNhHJUEGwSjt/kpX+p8FQuyV3
GDRadLQ1v6+Ln3BPEordvUiX3gO1dEaGUCECwC3K0iquo4ZWroiPi9xEV0RVq94h
BvcCFCA9JeqVutkAWcnHC7LlwB61uvSoq4H+dpn7jwIqzGQaJbC1po5c5etZjrrY
cwq6N5a23iTPfWpNiYO9hJ5RggKwMznv7zP8tLm+FR0Fb5EIeZTWmfJhmBRCpfsD
yAQWeOqttCs48EDyV+xVcZJ4eUhhLjuchbBDooiME5J7JQ5X21IRMR105huWVXPE
pHG7gvvwuqo91ABwV9a/kEi05EH8a0sKzWkq94pWmSOmD7AOdV84iOL8WBqCx6iR
bZsblgU7hpG5m3KkvKtrMdZmob+iNy97HNvtKxwb8SQs5p5+MdLtn0bvnAzckMEm
6decZiUKK11Bozi8b5KB6kYCZVA2dXCL6VSPD1/uUS1jmMml0abM4WOcGYdNDGkn
NdLjBF18gI9r5TNhKb0T6CSgHy/wu0NxanUmqcrZMBwkpdOIr6Q2DQOu7zNCFl2I
u4lO6STC5uZWwdat7ZZmpdvtsylxe8Gampm8dFD4B1WNasggwpLq2NLx0FlTMjwW
dhanwyqYHn6kCkHild7Td5hAlT6gT6iZCXaTn1XtyR9IrtL97DBwZtBF8eRpgkq3
f1gh3XEoFxnK9wyirbpAX7jV3PUzyc8DdHEB+7Zqk8xFUSdR6kM62Cy+ereitvlT
sDjoqF0bgelrSudvMVRfOo37LHsFnvZSfsoRDKkd7UCWSoPwtcFMs0Dmpdah1PCF
s0wOgVKcWcnGRunQ2H5ROqmBN63cK3mITwd+Dy2ygdAV9WQUH4LFn2U8OjkjVVBN
WXpxpyDRrQ+GRFYYPeqUVDa314E+AAcBjLfw6LNQlOQZ17iDukgYzVZkJ6R1uHg/
muxLwKVPe/xQOIVyiDrx8ek+gg07q8RpnQ/E2ZKeibnYp5oyECi5GuwgO07ta6yk
IWJ5g04UxZPIOflykykBoa00J9lVL/4Nm0hyAGPZOLWFbgeS98CUhbHqj1nRCtpl
UqJXfK7qYgxad3oyH6Ix/Ogxsb5kBB/t13P8EwkwcPgdbMt68aJZYzwP6k/JerkS
N4XuDU744SoWdnKgzg90rltsO9nXwaXnLr/nBeVCMvXB+S9yIh+WFhwT1jPFXRJG
5qSacUwQjE/3GgyVE62HWzv5D4ux77sjzSZknOBQT8NzOW2IK/dTla0AItiuKydh
1w0Iqm3ksIRcLTi/w2vg2xGP4+3aoO4U8P1vznuajoETDnpO5JbKpchbjsHOv4rQ
bmKCVW+DKCyoeLJYiSEsUFsyFz/Bb8vY8Wst0r8ZPe1cthTEe/lKiMW+mZKqSNN6
j4nw375KDvYzjNMfRlZ7cfdU/RMTlMlYPe4ETJ8IBR0k6gfOpDGnY/+DOB4lT8jV
BjdjDuPOEVrtSPmf8WWwWK/4Gb9f95aEDKM4g41/xT6/0DiQjzhd2wz8p82yg50e
0rxj9f0LzAmlGMHuTKggRnONXg2T0Ld/gX8oMrKDQCIEknLtF0RdVZew7lX9zYan
WYZMY59RaQP82vB0YlUncvxT/+u7XwXWxkBY1QofS1SiPfzG7owfKKzGflGck+k0
zzQPjXIzi8XsR6UITAWjFPTKzDg8uUNQ5pGaRmjk4SI7mC8ky8buodl9WMk8VOVq
uUvQHxQJhT2+ATR4USmutzL/w5NHaaVSsmJe4pHGaZRkQ8ubopPFykT3fQtnnNKy
HGRlsbrcJujzvKYY828oBAgrFtk5VkUOndunJr+I4srgvcrKH8tqoltBPcEHJozb
qzUxf9GgAXA/0aKr61d5RXr7iQzcw9Kdaf9RbeZGDrz2rsLlrESBes1e4E4/i2F0
6PI7oeQQFQ+0F4DQdaAi1LXwNpNqNBX6r8owUUSdY8lavohtt8Kc3kQ8rAb+uuV8
XbVDwACK0nNtSxzJNRzeP8GrSTJ0O+4JGTy67j71kZryFe9ffIE2TESchvFDJh/3
NfmBHoB4P6/eSCIqJaN4PdFuqLiDSRnBlCc+x2I7hKd5BpGq7Ja9Cq9DGlUtv12M
3xNc0/fNaQm9ZwqNKeZqHSfmXndTOIwRAt7faizIZh/f98pwHvA90w32Zm/nXbHM
xoxSJNFJxv4hMQMQvl5hCY2P63QNzCiBgJg5oDpxqzvT6FxQlumW7pbOYQStwMzj
azBk1s68SGoVrY8gpHx8M1eKipFyDNXVm94rNeRltUkMeWT/T/wAB/2RqAFmB9RU
pTYDBeliz04tWl0R4F9CehV1q1DTOCBuVQTmZhGxJN/S++Ogk/kdw/4kIlUqFETF
/wN5QNuey3qRbpuH6XkIAdgJp4mwKXk+/GfRC3QCl/RwCvx7VOv6JfKLvknR5K/u
NgpQutRnJy7TyhRRlrDxDbRn71d5XjeSY2QrhSQ00mZNsX+yequ1LB9QZ204Xx50
N7u1QLV0zgdVfTBtrPota71qw3wziZYMmRvXLNlB6ILUGOxceyPk4Z18KfyXPEnc
/IuM3zENZUVNv2L6ZS4z1u3GwDnQBjA5xdUwCkoc/dg/POr3QBZ/7dzYOwm+P80t
BmaGMyBdAq78f/kYJ5hstOC8GpEshviENn+QMV6PMQBbVOPNxDLXxo58ZItwP/Ox
ZGKofFVpgnNEIXNKqe+D5uk8bLIgtBuQVjqs01QmWXFw9udBujAAre7FG3SUDKx5
Ta3TqySG3mEDlhxDn/f7qAk92I3lh/IFvOOFsnJI7ApKMCIPTZDOqIG5etYLnL91
/fr/+aJoJ0SKYPcvTbffh50Rg+rbQD3CEF+um63eLxvaC/C0IzFExUnb/09ogpIS
/zveqlpfgwdbLE38KyebKZIvjgdCdUaPNaenIGTJU6BpuWGbzsFTwBkR5hlvALi+
Ii+v6uhJ68jj8JM98ts2Em3oTCKxF0sqhIZraR9PVOEyF92334TpH0BWX1/+CM4L
ciYspGn6fff/D/z5z1Ipy9gmEdkN3HI1Yld6uyuQn8wUdmo2itukoRhhaPKqDtwh
HxW1hLwDFeB62m4/y0t35m5t/P6n7tCeBpaDE4ZBzlv8u/w/pfD/oU6vo9iXURMF
tkLukjpqE6DKBuO5Rzi8urR+djrUwZTZ6x8b70uQJJtgq5Eq0/hiY1lL5e68qsJy
hCgw5MG0jxkPSvc/CS9EhS/krKop94oW6QVpnsjh+tQvThAsiWVk/gGY015gp+oU
7vOhJfiMKEgMCpK9sj2AhB2Zc9TsnkaZgVEyt/jxyA1M4Cm1G6HtCCjTBOX1Robb
Qi756jSbJGVz7UcN34SpTJBzB2QfT4l/eqlABKzf67EAHcyW6jchxSXY/qb6IqAP
9JxZqWuAgoKcoW5atvcM+LgSt4bgUcvW+vyjhIt8TfH+c4CWFm7bSO5Ch6+V9aeC
MWqYlBzuIvE9t167w6ULHMB3xN6pawiWFpUzTkEQLQE+yyIZoZFwQgKMZfWwQ9Ao
9l6kTpMpIZVeGrSvvGbrqaLpGNT1GIzuUwCMMxtol/+t1wS8t+oxtB2UTPJ5VWCm
so5C5WpmzgA2ZsH0xS8eERUvXbnfvU30AJ/cUWKnZ5vUaphFhCYOg6YpkZtPP7r7
wZrRLLdS/eZUl6RDaD0YF2JaX8gQXfuA94UI6RWqOOGbQHElDhPHDJb9K5dzvtgE
Cw4HcSODlM4JKLMeKKayTUW+kETpl7/H3V0mgLpa43BO5wKuZExQ2gTzMtfADqDO
oP2EAVY6zVYC9R9JhhX2XJNbwQma6COp/HlVuoHTt3c4a2/GZqkdIbSIaxY7kI2b
PGnbz4lXDLEMgGGZHWsqHswhxlCyQl5nkWT39JUARgbwJ2Bn2EjE0LqpJHqjugV2
sAob9SFoddCfMRdnB3anakDla2LufjP+9HC70lcD0Cpg+hcLaPq2rb4mm8AFemGo
mbMp1eEIOYu736Fv9uM6WGIz+l6KhIjIS824KdWAIDnRvrn3cEnIerGTtLJoW5A+
e46pSHPiXso13swzwco3WlsWJuEZebhCIF9GIg7nhBVhsC/h6fvnxn91AVLHl/jM
nJU7hy6adRTTIF5mCuVaJzaU7LiDyJQ6RjHj3iLEjuFZQ3VodcEKblvOotCtUHEh
967diHfOJHkTLvRBwNRGHf6LfAQ8PSIrXf8HGbIKRL42iYFLuUCnFFVnTcZLNPE9
0CIoAKFlyxHpgI7tWueO3z+xhjCdIO0T0ksq5WD07JLTrgZQk5VrhY1+Aake85ps
pfIWqpdNn2Hpv3C2fxIitTH/BI+Umb2dRf6F0DmlM5tM8n07YryfLMrDh2a+M8a3
tQQbs+s/5psVyimIjyw7T7iK9CLdEECTaqo5xF0FQeUs1kbk5/M7kP6GSRMV2a3q
47EemKhawjC/9dp4EF47/f9ckX2yb8naLzmYhwYFYhtgPnKgWKVzkgNTyUjgl55+
w9N4shc6GQy9mZh79W7X3la04Mxl+tQkHK+gcdnXgk7qfYkGvefXpCgF/CBeDtoE
MWLS3YJjQ9dIy4u4ia9Lo4eG+MsKR+hxc1CsuvKgtb5pnx5POywRDh2Eld51mhfM
CAZ0AqnObo0JHhbKZWEu25t9AV3HN4jBwB7b9B19wvZznj/fB5RKzDEJyFRViWbV
uFNCRIkdMuYRpzc0+GDNnOGghS3EHcn6x/bUbjZRxxUGvu+wGKkjxGGLyvJ5cByG
fOiJii0lYy7ZasnszcG1+yskww3NhwVBbAfBiIU8TgdFgbhDJIzrm6RfEaUBsAUz
mjSUMcZQiEjWzGeHetzIJ+pCjKamwR4ZaNAUReMey+sGbFXlyPndyHyG+Ykh8aAP
dlHrmZoto6cp1HIGiPUcAMdPi1OjCyV5r4JegznpSyig22V5D1XYmp/j6784v88X
r2NKimg4iug2vZQCoE4hFeXUN5iNGSHsOyPaVfIjcPOaR4Vgv7LgGUvEQIzV1qBD
q8oKda9nC8zcAd/3Isf51xXIQqV5BEL1ZceLnAclj9ljS8uj9Ed1BjLsVqdGEyf8
T10ECWJjX+iXQHZ8nwpWftX/+SebhVIofeRNvMiNUDZ+LCH93hMShiK30o0Adm3g
GRBjfJl7ugKKUP7V8052jnebztDdxSIlt3+XpytvpQY8TQVjSgMSs2fn6v1J5spQ
uHrt1DzJsHK4mR5Kej6ioh7BgeV5rUBk9hWWFRDrjTVhH22jHV9tTpc3JyC/OIrf
gkBZmSNhqDEg11/MFZTEvfq08j9/yjwDaelUg7oZyJkS3mD0YA55VOVUFcjP6pg1
9+WmxwvOSqksmDMOwBebbYmio+iiYM/J/uRqIzKo4jRTFalMKKgjd5kBGqPbF/sb
O+YA+FhhE5u5MGtKNNj8hfKrt+FOpF0Nv7wSSps+cipa0UQ4uJNs+u+8Z3x9lO5k
boKqnb1+YR+C7cIsGC2MHAf7gI1pl3amjTDuCVvGdq+4aoa56xM1uUEK+6fTmOGC
CBptK+Qnhi9YG2+8NW1XHW/XKZnqft5MGS+4GvCSSKen++98WaPbROsAXB9hCWR+
///IM+fnUxocGNeTeAbbQLVIZY0gKhAQI9ZF+Qph1r0nZaoSoMYo3OTeGRCamCt5
Q1VRj3mPIgD1UfPi64/QJqOJ6aPoLLlI2HXBMzWQAdt37KJdAliVkvDRM7MxS5Zc
5KwitlcrS7PAd5Qd6IBb2psZTjs9wxcCp9A8guN4Wx/4neJZaIY1xIZlsDgwJqST
/ywVJRgEqKWtBglnuQ6/hDez20hOUqf2h8AupiffWdiokKUh37GoylQJPklhk+YQ
KkFiwG/CnF3+VJlqKhKY8/lOTaEK2fRE1WfKAgqfEzSL36VQu6K8fAEs+5oFR8wK
AxzWstCBaISexneGV4Uz2oSYQIswlhXjTbQdu2mUep6GsaeOzQn9gusNt9wdePvt
yBbCog3A4YJQkWyxqMB9n5Iq225pQGLpP29v2rUJDkC/x/5VR2LcBSVJSpnyPDR8
tpTHRSVjH9W+BJ0DDBIbenPxkeCvacSMDb5135HwiLfLZ7wiYEzT6qJjpY17tsZy
lCfRWLRm8+L9WBOTViGSiO2cnFCmYM1ny+80oZmpTsHccKXmvVD0lCnv2v+/0krE
TXhUSLrqbzYeXC69r5RTp4ZIJEE+yUAxfnCgEqU2EBcl5qYeW5KZ6q69cWcWX0yG
b+mb3X6vbenP60WrsgjBRwa07Kdcy/NsYUygssUncE9lDajv5XRQo+V9XFG/s6bj
0nG3Q0JUwVI05LiRpMjcEGzT7azhYRAfgPKSdhN75+IzA8Dygder0MMtArFtSx2f
j7uiR81Ak99bshzV+tUcgYg+7A3a8vU5BdRWJB/OeDUpJdsSM6mbyp74ni44cLjM
enO4t1TDFhTnseaNBWD4uTeIWh5mLimDo9cebG3dzhgh68yG7/uFOaJVVfGELISd
AjMR59wsw3lDuNbp0hU7+RKvr+6UT3p+9OG++K2p+tstvFvhoPoVIHX9w6yxvkEo
BtocRLpqmxMl0chJmvVQIBctfpjxgZlPNvW7Wd55OgzEg/U/71wHfmjp7o0gfKzC
lE9VzlT89JzaAIxcCnvbgzq8SwqAToJpblZ4RPm/HJS0ym+avToN8Yo1Heim+an7
7JmHj094rad8nE9s9N8eNevZHFcfZkVZPpXe6mDd4Q7V/kcuBdg16TuQd1FBRSP4
IeMP5O8pmVM4xwVN+ek3FaB+sHTSJnfTCT9Qax2UEKVqSlSeefk///AmbpMgF1jk
nV+g7wfshztaDf98/hGAr9mJ1llcDUwdlaLnIZrNjMKgmxxEkIYYE2Ii+y8oy4Rq
zG4ymbnT9cuPwAvf2Mcxl9rimTL+Otb7XO3Y9UE4/2GOajjGWCbqu74MSb3EqZn1
2Z5qUad+eVBidQBL3dhwrLvZTO0MQs/uP0niGXlWoJekHZQLHj4xdVv1vi8xgtuN
mDHTQ7MaPz6+MmCR7AIwJqsewHhTk3CO7YaLxyxlYHZqw50/knLZKfJ239yKoXll
qS+qBh6R+eDLxY0+VSh8bradYyuTrLUueWLt/EykGHbvM9y6DDexy33W0mWtiTbJ
rdHd+1uCsBSOSzhg6ZKyUQxU4KOEM4w78jyZ6Q/w3KewKA60B494W/km8Y68JtrL
dzQYRjzt+9atRNcS91tsM0C19cP33n/QaU15uJ+ClTgvSrrJLx5+q+ti4EvOCvqd
L45CjzkQbgKUjuisI5Dy2hcTD/sGfy34xO3yhC2a7GutWN0Zgob3HHJIg4aEh4Pu
PXOkLLSFAV5ru5m+NybSYMpwYGn/OnFSGRAAp53ubfnDcu7uZMZ1sAX2/R4ivjje
Zxt7vMZmowFOmjeCSECzbGCahDpUNWx4/LaV3RIN0UByJe7G1J0gcHdpWY/G1BDx
KQILggAFfDRLOfSIfwDLoztT83L9Mb+DHaU3AnBsDhfYnnyJmj0sMamiAU8r8JRI
N+GbZO4tMcmU6bFrc1KVTnr//M0d9SlCn99w0GmjglN+dbHEuDsSIxkkaFqDXrqd
DTCo5feUutJNj98bb1kUmp2NAszuMO03mxQLlMa5NOTrIjArZQOLF1e7ZhbhTqHl
ECsveudxKwyfeSdEIaLROHVJPI38hawlJZtC2kTzJYf+YANCryl93WOCn8hSb8a7
YHEmcSLnlpI2M4pyFoLYudWNFmNDdEUXENhz0+IUPCHzcwLigj6d8/K2tMEJ8ASF
HRa1UoKBYsuw/DzkQ9PzndOEFG0R7Fpae846v2C+WDT6djJAoM5zO0V1GDpGY/Dk
FA34Ypx5/2GR8tO0dQGztWfhCaJaGFAWsy4ufDdBHuenp4Yulknc5MP6Nv5xeBqk
X3VnGCdgMJAtu2Dm+i1/7ZzkArA5mr+XtbOQpR5zk2pNT98QRxsxjs9Z+sW8VBcq
rxJi2M2ZGNNoQCYqvNNGHJQaj9AB/maNg9Aw7He+13UnglRm8YUVoywqnpU4Y3pC
6R1Wvq6lvz82ezX28QBEfboP+29wZqrlFKl4iseNDmukjbBvOLJf2trWbzx803Co
rUh+j7gBH7VHDgEkXCqy7QxGVrvVIq8kNpoNUb50meG+CXfGeBFErTOapNp47lAB
t9rvYA5yXQnjTdv0kzftTsnTzMriwYHCfYcTF1UPbZUElGk7GP5GqfeWyOC1mfqF
FADNA6vhn/5+ZVM6wkByuT84vLir3dfkSb8cHnlVvPMrzCmcBguqw2B6Rdsc9YzY
kEiAs5/LoY3gbhNFZM6vvEAZGk2B86kl7gA1KA3NEys5OsrdhM7WJ5Zk5UjEHbFr
fKSfz4rlmAtqyUTsFfJE/qBaTvciv+90jXoY35b9noirnTLUizbSC+bugftlpQKP
AQ1jS0IOvgQevDT/9jts/IJpGl28DBawAzPqJFYKTGfHLkdvYslpytSTD4U/NBg5
AGqfmAePmoEMQk4QPS/vGNCSfg2mXhhMRU95VrZZlA4Cci7m7NNp9Wo/phMS6O71
ML1W8S79vMkUOqNJeHLpdk2+rf2efUV3/MVwrpxqbgdQsgx+xFBKjkwORqW7LpXy
YFMX4pqfJEmfdkPThvdl6xP7Lkf0FJiKRqpcTfBYjFOVTfTHuTCfwJKozu1pMeyU
uvaaIFlzqndMuYlumQBEQ9EmzS0fwOfkncIF8vRy6cxBMFgGPplEvHHn7wYcLQFb
NxlQw4oCgk/PegM7dT5nGunVMh57vstZQ+L4CnlSzBW+Fr5vTaLiSStX/mrN9Q/J
EybwgOeZyvAvKufKy1nf+X9pnQOefmOD1C+OgZ58vRxiA4Zya5IuYf/PzVGX2JPF
OesTQ734Siubc99pr2Doxgc1ohumAzZlRZsBh5ajacD9Yp5Bp33iyBjS310w0UAE
64MtBtMKnuUdvuMbgUgZ2VLQ8GdGGlashL0wtyyZd2Kh6N+jaJAPp5MtD/bpRzbe
C2S2v2JjndGi9VWy03EMCgIhd7+Y7guB+uldK2ThakYg2jbyPx0kLooSafsIt2SL
83Su5P8c681DDR9Vk1xZ+T6jjj4JzdqBYFYwwtF3T/lI9FygkycSIShmUjkP7tUH
kugwlN7xMDjDOrjLDKGnkL47AyX/7CvJPIRLtbImfBkIEqysIcfwjC2TDvJWCnjq
auBUJEFkFHL/UTql5zFsF5RcK6kR2WZFWmZEK0sWPUoyjCVGXBDJHI5nK0j50aZ4
nasK5X9HoO5FqgGh9nt1v/Zj5gg8nROMoro3yvfd2qHSxpYazC7/mkkNo1DwTWQK
LtzL88MISbNKQGi0WwBUsV13EU714p/kBpfUSKYvIuhv1C2drD7sN/91kZE4hmtq
cYAIEDnR+9hHrSIsvi9itQPYSPpNfw6N73ij2g0ixYXw7i5DKc582RCTdU/Df0Wx
ImZPO15XxjoMUD3yj9dQwaxLR+WQh9T71Y+0hDpTWsuXhLXK56gyuUZi+drNN4Qp
eDXvyQDdxcj1Ul6OrNjR11hGkGxXPPdenDpEEXEyecNNhn01vIT0vhqT6oQ6f4W4
jMh9ZqVNYLv4vscSqRiMGjhrBkUIuodbLBq+FqeJTaHn98yRXDr1LuMIavJDyKoC
6gGknwGFBCL3+FM7jmUEKkztj3q+LxeKTe3s+QA51NPkhWFBmcksz4HfgGodw4CR
6Qugy+iCvyWxcbEHNA58BOpqXapqgJFyEGpfCWlU8rij04jqhFqJKFg3t6qODzwg
1ZPke1Br+WzFCYjV7OJT4FNB3N78m5re6x/O91fvzuMdILFOx+a36w5eOCWcBK9Y
EHElOeeoih9GpazN1ZKVmxnJojpp+cxsz3r2eDSXvfhsdQK2QqkslECdZ5UfqD8F
0p2Lg5NvDi/rHPoi7/+/SOuR9GFO2mhKzgArMp01q0h0XRhvZgm3PT2tbhGCR0lH
wxNXSom2Q6+QcjzeMAXct+CND3DDwsIb0EXfUNp7qdvAzdjo4QXXNKg8Ege1XM8i
KxCm0+MqLyochSS6zXuWcA+pXpLa42VgQ6hDe5J+iDSl/1uNPRLLR58x4HrsF0Pu
M70gwqBEukyu0kGP8QNs8BEfdsEoLt39i4wtW2JJyfgwcsQnhE36ypiNCoQTofuc
8MALRmIXi7OhW6JqkQ4PTT8D1tvlff/fjEfS/9CF995z2wo2KoAW8KBZpuHoln59
MBSVKNhHnfvBeOi6LuvWjHysS6rZJUtG/Dnp+RfUDSNFWc+f9YEBbvTWxqlY/et9
89o3d1RHW2S0AUqNnXKcyalWGueROyggml80pgAvbaE12s50dk7yAXtrrH4gjtlA
K57ycQ0OwD4LpPthpI5tSd20bcuIrjgyUYBAPCJUjGQEVqj2+0OQnTDbcl+ZMm+o
02R77qFRTK+Gp36scVKymIFJe4VaPtjSwcHwTU4hbOu3qxReQ8xyTcCAFuWzFylD
VWDCKE8wkvrgYZTmT54UOmqWy8qHNO43B40er24NH4cLz7P91DOyHwfJOc8tH8p+
JU+xtNYUGBFbEEeazutr94YgPMbXIr99X9QTtrDL+hlGcYyaaZXKf16XhExwy1ki
alw/cEF0fFxl+EL8vww9i4An0o0iWOnAoEMdJu4QmxtGCZEHq6JwxbN07JoHaz5A
xWE+442eaRehX2OfUBcMkQW13Yw9n7LZUoELd5JFYT9UqDpQd+av3sMZ5bwSEf0P
iIsuztTTtOcWkBOf5qJ4sApJtSZfTZAfZEbNp8cDRad+sHWrUf/p1b41uCKYS5Cu
aNfwve+uVt8a2vj2EOvl2bCyv3+hPhS2cfJlwvrUyVEGlK8IWKkQYg50s5dKVOko
qR5UVEGS2zsqRQMSy66SGhrnqMoQ12EBnBcTC3F0+h541LUpZE4IEGfjSYOxZmi1
325vn8EkZXSEyK934Q2XEm1hatJ0WeDcnh8Nt5Gu8/pjikw40qpPKbqBZwYFbbSM
P7t1a9xXnMIJLKVUmTUfDwOXcbdzCwNA0K2e743bDiAwY0am7IRFmdC6eqoIwfNn
M9JK3+3YoXnQF3+LEnZo4nZox0mcAyJu8AypXVkbTuxytMwzMyEgSVlul8XXcalh
zdKiybdIdsyMmMzzdgEUCDHB+psTIstCQeFNRtGX/lMt4XZNDM9NlX8RHOHRld6z
eVx+coj+LVnc6vIgo9lIozj1yKuhUFMLTpdiZNkF1YHy4CRE0W1AvDxPaJYerdvv
xfPWb1o79JIr/hWW9yuhACh42QttMaj/ZeyP1dzrjLXFc0CMrc6SM8iCToqM9njO
ljIna2SesTRY+GjzNBJv3X4BPb8/mCswAFWtdztFuyDuK7ZJeknw4u/1vksjtNxS
FPYMCs9f/UrEE1nSWoeZJhLsRuXSXxTdDIL/0C3J3Xc+ljt5s4m6RAcAWP8xrmUD
Dht2aWojxiO1G35pyIeDPq7i+3zvHv2AdrRSMj+fwW8AP+M/Qj8tF/3IyKJfGCp3
/WTXk3DdghYdfpBAW3PA2XLs51Q9Te44KWwWfp/pP2S6oj0CMQFJc26xExj9uKeH
/ySjeSy39ofOeIt2amUtIHVyBfj3YO3IdlDAExyo1p0J+eYKw/9jAhFLC50kqoyF
C5FFL+ysmWy8nuNfbaoBzy7rG5tR57dYaAKq3xMftxTXBZswpzDA/PIZ2lBBEQyn
sYJpUD7xbB5h4ItwkveH51uAB2o1+v5FP4PBKa0rGfiV1PYN5Ob0RIhNUxWv6STl
GZwuoBzck3E0AWQdBeTPS9fa2Kxoqk6xSU86Og84XAd+Che64bYbfBq5bxhnu0hg
9mQmxUB/LlvCEO01TOlcvo7oMaYCHeSaZiPL4lelrY6CWDKrriu73L6juFo7DMs2
k9hJ5ZODQ+RWt5E1M4etLhU4pV6JJlH/A0e8qTd4Zb3AfYNKM+8LJ94gmAEYk6ZV
9mGSvCWYATwcme7VcJgYRLPY4ziUALpp+3kdDrr5iEaKqRbw/oM9uxEAFUIH0roC
E7ztvDUBu0Mb/1BNof1AzUxp7QGswAWLpjmZb9Wb5533hYtZfLMPJCCxxUZC6z9Q
eZhal+5RgEeXgp+rWuorNFdAuyC5MNv2nX/5GKMad1aLFvDe7mmZcfHo2gSWGmXb
Bqa3RSXFPDSnAQ2Gbu76kyk3+ZrdcGibGBscq02h2kUSSMDua6rMKol4pEfWMTYJ
eIUf9iXfEpvsTY0NX+6ejzJEkkNg/X+pjcAJ51j+iRYu0sFXcHmp2iEf2bulZjUu
PrasUNY6LGum9/7IvYNqInV1U8mwfQR1kHXurR0SaSREVdcD37qu9Y9ZIyx/UcPN
FUKbJShnw1ukXnPHAOlGMa5iJsrlHGSrQ3AJhSZ/5ret6dntgx/KvElyxp6LnWwD
CPESCuEwhLimJOH6QaN69WuZjtEG8PJxGIPTsybLCUuVv4GDaD97I/OIJUoB8wcJ
1BN2s/1FB+RK+p8x/zgWCS+dSb46G8YJkttxBxBEFw0wZSr8+htXyyHoCKUgGTXP
c095gX63+Qnm7cXsBHMCB0PyaNN31IF5fngHvyCLdPS8ohs4IdK105yuzzksVviV
49/4eV4u08/n5YNU+Acd40RScKTcy8J55Ka2IcxzFZjC9riUHipZfxfp1RzeoAGF
OAYmG7u5VtrRn06nehT9dDRPIvtbl647qbkIIZJgD+3PdvAJ2MJTw5q+r7+A51ZW
x+jIY7c4V+5OoierDsr/Q28Px3+YMbU8dlEie0S/XDTn+U3GZDs2ZHckq2isyNJ0
WTwr/HnUru80aIh/WJqK78lG/tITr6ItJLkNB+f4hF5TVOSKjZ3Co5NAmcXN35H6
BJXE5d4ZEwpI19HFkwDopOUbmhL/57KgBmhj8pGplcKo6kZweyc4hkOcZiX/bFz+
2MHuIt5RH6jvxCSH84QtP659uE0QX8NzVbQFmurdN1uWCSu/Lu/LSRb1Yc2wcWUi
jUhyAeFW8mLFf7/b2igbynC/Ae6Sd3nPs5M7J+MjNkmPGIADPqVFunL3Akty89Ce
4MO0qs+Dx3/cHgiBCt7jYzX6DZdFUpR2nsDwwTw7Olft9Cue4zwMO7uBM5gQ6/xf
eylgelbIpkDzCwfAUG80q9fg8wLBFb5DMMRTzmw3nC/p+bqd/gcnzJcVmbgoec/E
y9yOOl7JFfMRHPyNKMl4s2YPF0V9VmlCCQxwtJWUfoldpV6GVhQO3gEFGxSNFljv
3wYbFOppSA/33moW6vDyOahLBZcLWYtiAeIqjO7GKPPOqTNGW4KY95I+m5bq5qYh
abhXAe7IpeagflAn8TnHpWlas1uSMxzMDC9vxyBy7NOTv8JER2MLMhCrCEuwCj40
dNQ50mTmUx7ZDiHcNYbw+5nh0hkFBmJXbfOwRDZb1bbe7PszosHjvgN1eaOyrH+h
igGGGjRPoXj/1PvTheIEAm3UITqI2p2Mp9HlAE91rnahdUrVMPWJc0RHVhAFNzVT
l09OSCICSK/xKe5fGUhE4g86t/MLktfKg4SAPNi6oAftVDiX2cQnbXNTRah4eruX
NlOKaVlo8ZfTaL/xhsDxK12zMkw+OJT6Be3vpedDV7sEuA2JF61RCzMygNOmVL8C
/VBzxWz9NR2E0jlQsj8EMnt4JxCN6noCcNrML9yb97u0p4NyuZ08RuddkyGGZOx5
RiXvK5TPZiokpuJihj8jns9ajYjz3pWuWwGsDCiZBGXCOHOrOjQBpZPIL0Rby/Wv
yk6XFa2LlbNP43AVkjg3WmZ4jQ9jhwGxjApHu54w4Cf4BWKeXLPuSK6JRh6OLK2c
l4iz/yvaMvW+eGmEvI/hFju3Jy8KsRtBxLyjCWQJ5tTk9kKFLIxF+M4nn37EWsUP
H6/P6ibQAntE6YKfMwo6LxJg/m4FyH3gIoWz9/YUkEgXbr/FqDLU1Vi/SwBqZrq0
/R/DS7HGFIuMqTA7FDaaUgc+kZ9wfPG9BfSwu6lDA0nY90nVe5LdHo7zCYjNgyfO
/RgT81RGliXBYs0FazVN/aMxT3Tnb6rLDzxm/wPKIntt78obKtVTh8D1nzcB2L3e
NpCSdggvefACll9nkQxKUr4jks4nu3IHdqkPuHI7OraS1PeeGDgbXDwSkb1wRbzs
HLGSAcx0EWrvEgXNsmrlnST+zu7nPfnzGSLiQwvD3eP1XXi9tRVMq8V5jejOUmcs
Bbx9RL6qW8KPe0ntjd/HTvYfk3Ijp2J/Q3pByx1kK8ix11vcsPlfExM52sJgkBs5
QZmi3JBWqhWXyKddeHWGZ1P/iu/WVEy5zXY0UpYaHN6u4EEu49I38waWgh6B4LO2
W3v9s/dXgOXJKhQJFxN40cB2j3Gp5KQ5UL7IDuDlziiUH1+4lgTjk5uRAZmsH2fF
rdnkwFKQu3UASx9Rl9UQ7wJyuPBk3wZMT+l+bHlQkw6d3S2fQupMRJxaZp7qvlC7
N2QHxz/Ufa1ZbMw0PN2daTKedyDbl4lCMtFH50lQD7c5wTl/J544MBz6wqgV72MN
N+B8Fez4TLE2DqVXC7HSvAP5e5lw9FzmdkuEI0iagaoRvYwvVkPPLT1dfyVi3cgC
h/VpEIaCwQ7dwlPd//OptGzcqQJYvsGn5XnIYRSSt9qqiq8qA1TvC9E7wHQddtbV
ssiDFsjp7tSl/ByNjY2KoLTKjaOACvkRDPPXq4Ks0tNwSGOdUIQmAdnvV4WRONsR
WiLT0Q/orRQ56PK1+4f8/LCqpYJ6IkWKWIYoD8mhjiNK55OzGD2r4vqkUDnHdP+Z
Y8eyL2poGW/7a8114cJcnV6veQRaQyKFI4vy0B8m3TqGQinkX+W3W1PBWs84ik/m
hTnI8hECemIxmIaiYoFHNQb2aP0SII7C0YQLLfHNmC6CyEzRPjP1w0jfC8XMdtpp
MH4bhl0wBE0yzbAOvn/Mseyh1iukVRIA4twTBrl9qG0kruey0JmL6aipkosqA9cd
+gQHAfcEsC6Z3TFIwvXdk642jgvYdUhVZudTiLHx8c+LSYxGyKNWH+7/AxQLfu2T
k14AWoSAKbmZQ4kDSyuIWhxMnb3NBwQe4eiflx+O8a2atvTTc/WpAg80EnFS4FJR
unKR/J+CwPLgtJJBtEB/UjRxMqfOpOgN86azKiMJRudCn7dDPY1FfslJ8WjmaI6D
vEfpICZ6OSpZd5Cd8+DGFTEWuvHqCsj0bUzDvCOFLpBGFS7IN66ODGIjhVgXmrCC
hXzs5+a1hqf0jVvlSZSjtQOq8ZV865su4M/BgutXRNgkxkwWW1aZ0EKRzwo+J/66
M0do37q+8B25oNpc1M7cY0VKcN2FDuB/C2Xv5NU4O40t7Gn91XzNLZnNBVplCgD6
FvjEeSWTtB9d2fzUROcnHYRE96ARttQ51MkkZQP3XvfH7febDbYj76bIBcGuDZn1
SWuswvqSQXHkHsvF0rXIDsPzjHSxOMnvfXt/fglvsbsFz0sG6788pLEWoeC8TQrB
g4E6A9suOMLj0QCFfd+tuVZ4M0ch/Riw2mWtWT3qC0idHEDSpYP+WFmKX4c/T6E3
KNgTsqMwiA5YDSeKsan80zhpaXvCc9L0NrseAs035c6CkXJJhne+oOYAscF4q8pE
lyGBUyj6zabgz7e/m4g6SA+Iv9UkU+7Zc9SgSmOY46iqP5y1tDqA+8p3JveyihPb
teaZwczZaoMPR0MW9VJZIVoDrfKmDxaJ0J2NszStJTq1kpG1PSdaqOfUWMTPacMK
XgrLJ/lrxVrgGyaYIo03dN+9/IqZkbh9Z4dIRYxFGaZz1CK/l8OVxHURJHbF4tY+
1dhHGHJDQgLogXtnfCzuCb/jb8+L2fqerYVdMOm89p3U0rYBsKH9eNHTC6fYUm7c
aXAEEhiX2TprHk88Uecm43iRWmvCfl/DqaS1bTfNySBCAyH7MFdC5+TngD68UOLO
BhJYj6sEpsSx2VQndu5oQ9ExLwS47rqEx2h2gRlYmw1M0eVcApLMIvYC5tzgKUra
XZhD83qbKTLknl8wjdlQTszY3uqnXujwMGK1VYF/Z6quiFyPUJemuJ9aVHggDD1H
n9R309DCwIuB10rBzOLM0/hay+uYKs45xrKTcKMV9kuasiOQvhvkQB7s8wPTE3+D
GvhMogfh9mQZ+/KFdF1t6ykb/9ac2sXSafWZLPVV5o6C9AV0HF5bv6tSOgGkft6r
AaxfvGOEMQiEQnOKvR8/3lYDXkyFUQodoep8Oc/6MUcIbjOB1g5+ouThijaUuFKy
Ez+72bi50aVrHNUUBag6IU1RjWk5SSW3UOYFCz0kdnhHYUVYfJgtKLpws3m3Z6Xq
5pPdgGzbWwRPHaxC5GuztzTfE7+G0UFlhoJVmT4otNFCKtfbQxSiqXEtDQnFLMfI
Q/uqllHoMOYLznPHrinqb5+2GDwiVQqcHAj/143vfHrA2ocoQTKg+7y1t9OsIOwC
IWFqqTNCzoSqq5epowtf3EV1uR2JV968awb04MttEbQcJijHHCcAIwSMtVjPq+Vu
2oxrnNDpZg09qL1JzYAXQ3ceOukfrz+3GQ/+sy+H0NfKkUO8h0a55s/EbjZ7/6dE
k0lpjjZ5nL2L1RS0OsDFHsv2M5yZkIV0Ekpwp1Zt/82kCB187AtYxE5jKTydZFor
dZrt3nlT41p0nArhccBi3DNh3L8gLPUwy8CQRq6sINIfrT02Xg7mYwGAnrIMeQ47
FsvKVwVt4vGeWngiG0HEUF+ImPcs5Jkyi1SKJiTLM0tI6X8TVtWY32a8Gqk39aOH
rWzM+CHiqBj7kiUDEJMcnTt0Smi4ErhdtuaYZJrTxHiXO931NW24f3issjXqm4uD
2ukxi8g48cK7S4zsDNu7fMuKWP3kHT0dIOzP3x/o7yOJqq30QjZOYsOuxuLXn0c6
OEhQWL2LblpvqwgOTe7fCqHxqLJICy02x04C6+OmfKZ7e4Z4jpy34gFJdKzFDXOt
XbmxbWU93GQTP6pEY+52TTweDkb0z943WYQwxHnwyxdYBY8wgU7f3pukPA7MZ5Qe
OqXcNfRmE0TRg5dI01a49EOBaBS1zPKHTR69BxehX7mtXNvZis1Ns/T24KWMcO2W
CMR5IQD4WHAmqYjnXFfsHUR+khX5fodb/pjs+1XuPvB/vhVMuntW94BLnfyvpzvv
IgnEEXlIGnub3ff0cNJvW4RFCAQIb3JgRZgI/ZxFlsHmUPnYSrqtYAa7y9atLgie
N5bgdTgVo41vCmynqDpZrgJ6jIfLo5cHJsFxkvLwnpEGzNmH7VVgPvG5M6YETsn1
RXGKOUF4LwopvSvQrks2dxc3hRRnTadpjCvUSxUNJ6e3kGRQH7+cPI86q4mH+zos
ei90SCXQzXfIKLaY1zlTGpmmZRNkG8s2psfbcUtsAW6iU773NG6Ieayq/Padmuwl
kXJLGu7MAkBo6O5sO2VC4pz1dIbfeJTTNqbXGDylRZ/5o9kDUo7MqwlqvgvVovWi
nwV6x8/1ze+xykBYjeJalp4fm5M7a04V6VEHb+cdF8vND37+ujlo1amaPEWFvJAS
pKVPD/P2TMqq0tnZZcgFl2lIawI95tBvI9XQsmioP/2eWLrmI1x96xm+7H83Ow6h
2t32teopq0EIKcLQLZQvrBwts6Zzezf/LMxJ0Op2kNWj9jMqTNtVWxrsc8JRfllC
aS4sfE2f6vfE14etDWqejdQzkdSDXwWdWtJJ0uJ2VK5rwxoUX8G33NIw2g3o799f
C/4W+SO2k7PDQmSQDicQLxZKqaFqf/FWxQPMP/DAd+7fzipjhU4nUZr98Y19gvMd
nRFkmx5wL7X7WTJcCo8kQeCiWtC1zcEJGoPwIWDmAiPmYQ5FLgnMjg4P31wNPNHz
rB6Y/Ddx/ph21eC48ciWU1cS3ot677okZ2dXwXAcIhsQ/HeZQZjg+FT2Mj1wKw3h
tk52XH9tQ4evv/DVnfWFRbhwyiALRKIVWVKSHrKB/2pYpLGlXe6Ob2lF6pRzdET2
7wCx99edRwUMu8/MjJ3UwuB/LIJiQz7V+wOPExIkISKTYrXVcv5m698NmyM2JkfZ
iG14G+aCqvJYWDW3+Wsh0R0jxjx2npMaeosmx201rz8lr4U/9iChYaYENPTT6E8V
4GbdSOgI591u1fS7KRei2mvRU+FsXpmk7oYW2KgmqnHsw+ZOWc/BkIzrBsIDScGR
ZU7wEBEQmkKb0wDHiR5urzoTHbjndCqPRSkl6V4TgH6AcBOPJeAYaYwWB3V2UnRA
nMMuGCWNwhX7IB8/FhhYdpL9bU1OBTV4CCaszB8fTuQ2P2Z43wmt1HQm7unTVkKm
JlDMI+8CEuZsQXpQiIEskolg9W2edMP4UXOMmzqAx7Qndg9ONSgJwl/i+Coj3daS
JSk7uR5B6nAY2YFXkg7xOq+8192+8QWHFiKD8fmoIDDNMaO5v0kyA7tQemeHsalL
hErAYWAvwfM4szfBVU/aYRVEC1hfmWMflsp85HhKCLIZXwR2io3xqGUm33D9uq82
vTMNtlb3xYDQ2vI39WnNAi1rUCVoN3HD/6ft7FBW2jyKakQnwA4AVDWHn2XKvQbT
iyM6ypktpIIVGQ+y/qfdZjJ6NXdtUjXt6+3Eaw53jXh4D/Nu/k8svgKU3hLGUzkN
J4bThiRWQ1/bwECPkwigkA0/d0VId71J5+aY2JJ+fXtEi12W7Afz0VUD+fJlEVei
SsRiUbcKWRdmv8PpN11w6brn6qxcJIZCLdNsGjU8aw90nhSAWJzHREitfHUmX3P0
eptmeKpldxyMdAQwvOU0j47bj3qzqmqpsZ9qSz11Rljv5SnWEZn8JTDfzyrnRQAk
We/lBS5ScJZZ0UW6jNnz5ueuu+jxBpvyMAqc6pg2iT/wpD7EZvoIp4+JbImDwJgL
Kqh7067zAoBYaSxduC3uemAi+8vkkl/24iB5B1Mhzy5TmBK/gp/IWRTv3Wxa1c1i
pSdmJOV2dfG6i0ahHTw66VO3hJqRIFfgw8eDxAvXDhRm/UHFPr5JYXMnx5bmsgB+
GM+9tWrs1um/XTnSdhCdixeZa6nFJ6S77QQoMNloeaVY1D9ouW+/MjGv1hCxE3zM
k4cVbVbPJNSLzxn9gn3eKAChqX2X8g/W7rPg4eptCJ6Dra0lRON8xQgakTY4M9/W
78SpJxgesHZaVCguZbDoTVohAKRnXb5c1P/bktHsm24apCegaKFtX+LwuA4qis3t
RI64zH32TRHggeYVTgscGOH/DmmIEA8+v0iVBZrPKSFVvDGxeL6OwI9dyitC659q
blAa+jT7ZeVEpi9NQMJiqqovp8FSdTECW9gKIfzRC0ZbWQGkx/cPLEsSn4tmBwGJ
xXbebZkGRwtdinf3SbU5Zm3axlAFfhJM7QRGYqkUEwOxsSrTPgh5DlBYGFbD9rMW
Bt9umhFFrErMUeFXtrzGXbJJvr4nG8cNcdrPDmEx2/mAWO6LmL+wPEotRBRWNhEQ
KJP9K6xfh0cs55a5wklFzuKv1Gxvs1GGKWq9AhpwMCmKcxXyxRj5RW8BJ1i9Dxh2
DJykEsK0g5RvNhKWCLZsFv+bJgLMrQTjWr3wSdLExvu1jNi/k7J2iAuqosuBaJvQ
GbNj5AQ60HvsO2qqv1TIOA5/8RAdGIfZcTTnFnKoCJi25KVxz5p4yCZe564EeBAR
BpCQLrIaUlYfjGAqNOCaEreUMyJUoQ0blSiRV2MmwU2QRR0n5Jboxl/H8mZ2kyyV
SEeiJgt10dxu4Irc10wMLMXn6mCUHE1rRvsBBx40fOO++39FJVviiOEOCcYW4dQS
cyA1uVTWlsH2QL2eKQQ9Ag0Y3SrmeqB88IFhAeDHKlX0gre9CyS2F/x7jtSGqk81
ThMzCltvNqrTDpAQpQvVvwJQdEiNUTkuiGBTlHkTNNJfWPsGByxIgzb8DO678AKC
mTE+nGBRfWTrArSxG0+LzxzvoLBRWu4rBVCuzmjSu80clJ+FvmDkuoKkQk9Cvg5E
OxftmGntxfyzVlCheX+3SKhU+Kb8UDXYYlik8sAf+HGPelvxEBt/Tkz1P5To2Pym
6TLfZSBvTbcysZ5kpucJpDdJ2YPkWHPGeycm0yhbx8uKRG2csXoYsLiNMtmrl2hf
MEw3nfgXjFT7pJsmzDRR6hFPWzuRYcYxI+HuHYL9XTLe8F1yDBnblRzqnVHDmVCC
tP8TuTzxCD5A32d967keJQX6flrlanhJ0bwpF5x8l+1obFfXxw1n6Fepn5gJ7Gyb
s76GQxDiwnw3WLVSrIIJZt84CyLIsEA+dNBSg/iP6VRK/UVz9Of87InaI2mQc58s
G3Sn6kOKsPpLbK/TAxY70af4cO47dS4c36n65uf1tnM/VI3Vx0F12q/Lj54HwuGJ
9qYIaOElGwjO0Mz4BjG0tfZx1aXIvSz3Pceb5c7FzWonJZf645w0xu7GmihXFcvp
jJaZj3Znu7cPU3H/ojrGOlM5B0WzHYRALGmBMUbhvnkUIBbmVYDzxfz/aHyIZVD7
qD9ao0v5HSpdcSUR9t7si90sBe/C0TvTKra4yrEpk8tbJDPQaUgEQQmsINb0lM2K
HyqIWuanwV1vhJw57K+bTE7YsPzfnvJIcidoMp+bmktWICBHLfc0/xGBXyOhHMfM
x9EibaxZdo0gjEr/SMh9l/O+0pA7CfWr6AKFpxKxcBqQBO1y5sXVRZstJdjqiRQN
NRYvY7jjC2u149E+Sl1ddsu3fRl69m2HW8vEtGeKopHLH2+3NIPRB55u7my6+pFv
K4p2LH9fBZ0MXJouGVVAgKjsIjyAGpgin9Q2KvW9mMgCEbrNeACaiq/Y0nZ1czGH
Skuv18/H4Ys3nrMrHQWrnpTBl/cnzIvk5IXtkH8Hj84ncQ+RjGWSfflN/GZDTXc7
ViHxf1syuIHy1K/yRjIQPxrerfLj/kmUbGI4nntjKvyvmd+93KEnaE6pZ3NCoGK1
Ok83hd75WA7c9ENjznuWrcLC4UlZDp+Lcz2rX4fr72vnw2U7yL0oZ+EUw/0ibR/v
p+Fd1PhwICY5nc12v/jETrrOtzlQwF8gjxyWpQibE1NXxOVfEdhF+g5QytEWJo7/
O4Ky8mqoPwr74e8gvwyfKec8ipwyqoQtOX+s766NTORAMMQ+NrHzzesGTmsqNmth
/aShPFXbpADe1Fz9FpXFyu8glcXARwnm1TKRg1GtAzXcNelNFYH3kTHHb3cOvBeE
7lQJUJiPGv1KE5Q2bEiz0Toos8PseV0R/AwGePyvZ5xBSvBfBK6hTrtJQfwz0VKL
7hsNzAJKHO8psBjRZN3QQ35btf2SF5RXILWrSY5ulwwSdDji5ZCM2KqrU38t4UVJ
SmPlc+kC/SUNBvLKJdguLzIfRjrg0DqjmqK9/GNy7OfNU1rlhCZhqks8XJ700fbD
C7Q56LOSm5QAgw+tZ7cn/tyAoLDsQDtPOG4FTkjY3ldGqwwZWljG5GgO4lQ+LVyw
4SNtg0k5Qix22lJ9yPBGCGBizyuqpchJe/tSQqRGwO9Z5rbcSyvm8WhkxbIfGDhw
LC+xe45LMs0WBpcVcEuf+vqY667PeRWuFjd40oUZuLDOcwcbGEtpq1IUSdAt9b+O
1tSWt7uBKEtLefrFQUlY8AtXtcdkrRhMqP/ZhkVISxVQXjTSy8N1xwJp0mlUUuah
Vj9wzGpa32kdjH/ADJE26AnqtcB2J2Q9ypW4bGT1cy4tK5gh+HfpNZioE3PK8l3Q
jM7b+m5nmAGAyQlYRSHVRIMRhd5V6XctPFqzHdZDL1aqGJd6bElT+ALzpwUWykG5
LDaeZv2IOC/ZwtMeF97FS0uJjmgAkp/dz8gqVXrnw31/SaT4fbdRU8LW4MvTfddD
V9XWZTFXbm2M1GlXY3aDbPNaG/xBNIVepLUHcFpfJLtXPPIwhSOiSHPCt4OuTAQF
ViaSg/BFJlT7Pq4NuiqpGJWXVUAFepBMPIhbLsd3akAiy+3qrDzK6zRwkK0y8tSv
p1/RcMPVFr2AjVdXIEvtJoRziHqhLes5xDWMXMLR0rMd0+tRYfD2mk7oASr/bFYJ
4R9guhAE90QKIQPUhx52PU6vH1nF2Gb57An1Z3WVhEA9pIaVxQDENGu1qttFoesX
Q106ahC3twBXOVt/UewtjchzOiFjmnVzXIPE6NmFyiFrPmP5BtEVsM5DIXOd0pzM
3dEVWljcwF4l0JDLT1eKiyfvM6XavWz4HgoK4FiTmUySwR0Bx2NMwvBPzXqByVVX
6rVlSFMqSHAyGQxTl6aiJLoSee0wKtU7qtS6x/xCC6TLy07t0SYQfB1iWb5A6cm/
cO75VwZTvZaAlGyQ8SGgcdctzCWooAmqdKhmwi2y6gEg2H4uClC3B49p9DWAMQpf
1CqT1qXEoxM0ogRBe6SGt1Eq/UhjO/turQsTZZxJlc3bwRpXzOn9HjRBR9TIfLz1
ADPbqKaDMgbEk7XItRVXOWRZCQRDLzSxNQCRJ7jGcvDksW1OHEP9sqyHmw0OBjro
mNMq9ianmTdNQK98HP9BNcLJOgB7MaYNRZDjn05rUk/UhcFvrWP2Jy96mWZRVJjn
JxYSfs58MClvMcJ9yOPAQ/L2wd8adnjGNO36NFDXtZ42oeYYvIbwP+yNdwr2Rut5
BM1oCNqIiM51UYaCgL9iiGn6KrmVOZB5j99EWX1j1lOtx3qFGc9ln7KYSwZY818z
95E+P9nYnAb+zYh87RxR99mSEPPNcBsGDSqYTYPyN3ERcgmeo7Mqq2oAlZc06LFw
xe97QhsBXY/b5u+DaM85XJ71KauWq8GYdRfHtJx4GtnzWsUi+bJiU/pTpTCUSKJi
TL59Fr5IvYUOBjFIYadTgSZP2L72InPg1o17jE7EWrM7AY7UR+2Su/6HoYKf79fE
czkgqiV63RO9ktRHrfsnKCfLgZ6JIvf6SZr69lli7VO1tPfBmkl3r5HauvNabwM7
kHU040DYYqWcPy6f9GxAUKzOpQyKdzmpxyOkL+jCYckFvOSarID0fvHac3izrNYv
tEiA7Oew7z4c8mCjzy/MlyhNjDPzg17RvB1g1I2eOjvw8cMazy1MF8eyiq5cl1iU
6orqx/WOGCRcGOUFcSQmnaYs3JVyeBIpQegT5JhbhW8PJFTln3htNswYl7V7ALIS
o02/iJLJbn/Yzk5NyPpgLtqQik1lyhkIIyab+KspAsePECVGF6NT9Tt6gh7FTDlj
41YA8EWl9L0XoOACCityjDCE2Mne/3AuXZ5US7LnR7fwUrtpYnkbCZG2kVvJuE1e
+epdmyDTw35jK2aaPLDW5SSk+79R4H4CgiiUgB3ywx6U85U0PV8Bi9jYfQAj4ptq
QO7Gx5KOGBkSJfl6/SMRN4irPA0Lj55BkX/h6u0JDA1Dczk5lgKLAEqVLAakU2Ma
JmQTKNe/p5i7UNWIdWa7RuCXrImpMeqtWUewWTzMeADIGGFiH4yiQgN81+W5U4V9
lMX8rJX2sozM9Q8sbeZCKks5+wtCyjhvG/T0JDA4JOUndpg4kHz4nQkXodQjDhfE
8+PDe/hFDzECbuhKaJGjNll2X6BMIhlI72M+1EkTIf/ejM5yr6wtamJfqJqZDdWw
/iET2UQ5tdxEtxsUqKsJvBK/w1czTS1CYkh2E6or/vwPcA7G5vBuZhiv4+nK7z/b
zGzPeZCus/uDtHWEJf7QWoabOdIpguT88AIYCbS8f+S8Db9UxzJZFloZQ+itBoZj
KEv1KEmorNhaKN39jWh9F8Rwwo/kH/YfUcA9cW3JRk09gsNp0aVLl/7JnncHFKUK
4xyYih+PAcEjb4mfYGSIwwBRBZZsKtUkCSeR8Lk8xuer34ag+s0s21yXYpzxbxU+
jurIbj5I6SDZbZ7e8m52u+O5pe2S1QlVcDxaLNS7ZhVtUgaRa1f+kx7buowEKU4a
9EqI8UpNjtvT3yaaWniBvkrbHc949D5trr8g6lVfe65852r7OuaXya1JkJz+/4SX
+J6Z8swlEKGwmtf3TwTmjKK/KLFJky9aA+ZEWgVXCzIoRXE3nbKh+XIuN3gUDTPG
GttfUCZgd04OkTUjnfgICnw82OpaQMddAmuUCTBwlxVQCg8PFUp+BxtD/YfR5GtC
vZdqG/WB+nR6Saa6TY90uxO9+s0tsmqzNyNkokEEbnCHGXWrpGMZGyK36efO78C1
IEDr3nGEyiE2lWo+9TP1P25FUbCl0da2Uv6nfHgd78F9bea/v2RcFoSg9gNihlKi
dTK882imLbDrGadGNf57vlpEsJ8K+Pkma5tK1WlyQ76fezUbQOML8K8rbf2VqixY
mr+ClxTTGx5u6fKSOHZih9oWTdUpeLB4Q0RYawU4Fl3M3yYVLCFSg5AeP+lpKp4C
BRmTqEA1WuUCM0X25qEGDjKMyNdeagVwP2k1bs68HdGENAuKp2vcxA2kw/Z9RWmW
ZMxgY3eSjqskIdym/FevMD3Nt+jYDED8KQajVZ8a1MqwPeIQACkROv1LAtC/0EJv
cFFqqfKzn3K5zwTdtcpqilAfr9Vq4+TeipCPZVmWhHjr+F48lsJyaaAtw6weWnL1
G1bAisPTDVpl/y6HqZtt04oxnk7fdLXxyBHTnLddHP7ravFx69yyvmeG30ke7aBj
aXRhLvidlzD7YeRsuQD7RSBtZjRSmrzoVCK19PPQeJnc7EfxFpGgtD6W4zn6hsQk
jlscGvil2ha/fiq3EwMg2Q803959EKMowRmBKqzYpOwkx3eqyF7DpJttiqYYef/d
98GolCHFrQ6Z5fbN2WOw+k2sebIEqoljr3Lj6cnpPQi8oxmtfeTVGx5t+Ly9qhUn
ncYyGz7z1KCdiczh3R78ZFU7RelZQb6UgZ0n+bvdlg9gACM2IFp1AOaq721QyX9k
pCPYHm9YJzMICPDe1tcvGri8SYR8MOMKODTyMlxdaRuaoYYV6YthxGkiyFGY9ivB
h90idoYeDvyQeqDSRT5vHf3nuTOmJTzAtg39mkaiin4P+YRQOwSdJLIvK3biHXDV
jYdEaU1K5+VnNMed5ro0HmjhTa161tGuYOAbn0gJfq33RL2IzZv4ymubFsNW8WZe
3Z0sPMDYnf0Fh+TTXAekc/QTWkg8qNv2IQ951IZeC4BbV24x6Hvp0G5UeN93Hx/5
V0ocvnTxbDzMZaHUIU+VlTZooJBnAMgxY7K4ALKrF4erLdlGZQkj0SNHmdc2ih3N
YnyUYPg9Cjbmjm3lZbsJYqiEbJyHTxBskuStLeHXrfjrkYnkGc7nbBjc7g8BZBMX
RuGYV1v2wC56cadDatIaXTyh6eD/yPOffEl8J8JI8yLsOog01xJLRyKzrzBSOAHW
diO2VRzRYFlVLmv875ObrSmXFA2ShyZ3JCrgWbTv2AqiiBDAiNOv44KCPDrDuXCU
u8hkZLBUzNlK9tyfn15yACVMXqQDVsC9WtGpKU0ORxqUZZa1I8TYfgFh5cVUp+N+
rR9Eqpoy332oTK5wBfrO7MaPDaZmN2KYshC3itSM/czOTCI8IrT2/dujSE3lPDN+
2QcLbjl44n6BCXZWGJStdSzwWzuBlnIZ/Rb3h93wlSAPwSdvcnlC+wyn+nquefak
LOYMBMuZubMrXNrWZBYSZFn8FYTGp4XIn9+XeZgq92o0a9efyxT9HpFD72hN+Clv
ldng0+sP3g1usBSzaIaGIhs1IgYa9riOGPaA5kOV/Z8F/zwkmg6s+WbMBlUFJtQ/
9ItMaNI5wfGXSeUnTZxwfY6+5/VFAh/eygJfmyVZ8WTfRUBcpjzNHZxy1EchX1eN
75KRK6y1+n1eKN7qArCbXRASIGrzuKsJ5PhNqsnnWF4hIhnloj+KHQSgHT+S9Ajn
RJdYIKaSIwEFq2xfSB5S3UOoyZS29Xw9iu7f1WvYZFr/c/fM7qIXv7s3VOUzTfMS
K//2Zaifhg/KGCc7HnfVDwqlTt6H3Wx5gPK9WehLVSovoEqNGo4eBi8wpeQ2kR3Q
ub3chDaB7BxJ8EIhIMeNzOUy+43NUdrZR8+9zYCrRauJnKTaDh3iONx7ap+V+JUN
vfZqtH/5eL0u9EpNKLKaWIYY1No5cgbTF/wAzGIWdrMk6WZakyNCwJE6ie6s+qIA
e0zFEeVZrTNOOh52OofSHAkS8MW9FKz52Mv313VtmSxwIZaxRuN2TRCmatPujHvO
Sg+Jde8xDxCoudwkaBR0vRDye6ouK6vTHJ9iF9jZ1pAUEw86JcKDInt3jAM5o9VR
uI1W5NKNmIupSiWusX7sYx8fiLimoB0yuj/JY2YE2rcExL+VMLJ9aoQwv4mj2wqN
YewZ/AVLNuMfk6NjPWjdlEkgjZiVfPEbi3N6Z4CcSmjKFySTtAUR3SHHVOyicdBK
Q0ez1l0v5mrwCOXPsomH8p0b7+/md8YqC1/vqhQe/t6MJANide9uNKH9B1lk3gy4
2w+FPKaXkZMLNaXNFMmYfWocbfl1NN7uBcJxaap7IxnU1hkO/rYj88H1JtWlrltS
x3dT2fKKuh5YSCyGtQ6Va3gLcFcRGGg9mvhgKdObTZkI1Knyf7vijQxVp7d6rzOt
4QTG/OHSBzIVSjOXcL2tWlYT4YNtgtYGQJ0J0NAaahxMHAsp2x+Txe4pZpEIi8U+
SvL+rcHzBAb4XJX/+BuHoBkDTsG9BQoBsoqQMg3Dcb6eskOaH49s0AsaNzSz+S2A
6+QZPVKKp4xL0asLz+ipHaK5Z0wyDY6RR+r/ln+6bXDBNVfZ0TzwkNQGhDlrUm/v
VJbuHvoD2k5r3dKeckvB20rwDeHm9cHIyDAPQejK8dLbw2PlT7hgTUcWYefaTipl
oZJ4bfQ4eqxJo68IypeSI1AxL7F2XgCp6IxxdFnnD87i7atY3HNZmsmfXjGPXk+W
ZwsP4X3/aacrqoU0UVpOHtgr45si/qrBj5wu0fHqEeCNir/kWVSzSaWxVQCEGLPk
FeQId4BaLu8Jf2GDSqFuJJ/XTEk6NPo30pZrRozBdRojxbnpL0xqOn7HbDdlT1Xv
i+CkH9mkWmpQHrWgjupl4pHkzBtzyNUkZusiBOBYgF2+VPbdg1aznzW0AWQO2kpi
dq35cCRFwPzlw5/2B14/cAJtd3TJwHqq7yhg6F2KxR1L3ycthlq3PQzS0dVzsqLH
7nXIVsR0HJkgvA6fb74y33QGuh6Y2K4GwBq/BRTeihtb0Z4e1ZLKh+HSxhF8eE4I
80Rdhkl+MHCjW6dysKna317TXbSLV6fSG1IddvZQ4/iDM2aQzgKPY7/e7FmKbNn3
RJ/Fs1X+f7LDdsFMp3vb/iym+VI44tCN7g1SfRDOSTZg9HnCF4MMEhojEYg/cm+k
b5cB1S/IB01b5TEI8itL99PeNLZlWJ2jrWwMgtJqK0i6u5+1Mm4Q4cL+vo6k3vsN
NlJTztGAx7vEqc0144laokzjlPgNt/ApF454HdxPeOYvNDTxmnuyH5ZTSs6J/PFn
FogYXLgxr2QelSzvaiyzj/mf1wkARLl4ZiqXx/+97bQb1kV5j+kxiT+Fo2ltO1o6
gPGytGT9XeAold6FUNORdbRaTffPTBAqeEnCb+WPE0ka0AGnaJkmznmyz2xdZ+Ln
g9BmabuankIIMAFfvjHs8romvrQvN94htU3gDp2Y7KLE+pZolBQeLJxwsFBJGuKY
qG3135D9Tnx4+x4epOiJL+IdoidE7NWf8zW7D6NCOV+AaHyK8A2+wdX4CtliiYQE
gdW0JOFeBWshXoGywoDfJr8b5e/fd6S6W1JVzo3MCU3Yw4BUImqeda5AUmDw5+hH
GAfhAajfHv3JhbCxAVDzK25Z89b8PzATZXQoJ8R8otnZVKQQilz9is/GucT4GjXh
YB6sy4+tSeIodqlRRnHuHDjlpImLo3AYPf1CNSfY/D4IDPsjhzdtu+GWn4GItZNF
qaX+Oy7I7Iv71PBWa51YVqjA3XWR5wxJYKb7p6VZT2ojtlaO5ie+zcfsY4zHXzJF
3cLaQe0AuCnU6P6Scrjv5+qHIRSWSZD11sXgmpfW4gPUTaRNrNcDbIUFwpy4Yoxf
gZ3AnXqdnKpKG+ykKIz3MJjWsdAetTKKOh17LKL0iHhmbL0Ny/JBqX6JwmAgr5Vo
/5di7wF7wTM99z9mVkMd0rvkdqKccePYDfQdzMuahNPLrLSphgCpEA8/C7Euw4GP
pKgvAIp6Lzjb40RBZsTixRUdr+6epFP31bY5ZOlMD+lYY8cV/pgdkkO+Qvin4LQF
auwcqtJuOty9j++7YeUY76gjZWRYrihUCxgE/8xmy6qTXscZ19nIjMouyaMVkKzT
m6LjVqMBGB0oL1gZxytxmlQnHJ35qTpd9wQr80Wri8IzoMG5RHTkAueEJPpf6os6
rximtxePqQpOMqYhuOyzibdrMrhZfmc9Z8JfM+xgyTTWMhhhosadqvVpWiG8JD4b
0OlnUMY3z64JSUAiGsAeB+5NlQ9bf/m3obFn/jl0Fv4TV/6/d8FtdVYmBmSoouRb
jUMYFwCFc6ukQ/Zz1XBheQQ4cKaaQFx9kMfIc0+bWewIKH3XNO4M6mvxOeTEmXiV
phagA7uNYz599vv4mjajO81GRTfJdr5leCi1FXqvdAODl49aDeSs9jbhUakP5SgB
/5VGzLf5LbENSTiag8ldyiWig1T46lLzssyG8/q31KUzcq+jofbW8CMxVPy7Hi5i
dNE9Tig57tuIUcU2lzUc6ACTMLPKfwdHODTNAmswOE5SN+KKull2haaSh0ZI5XgP
4jysdJY6LZVikH+STDQYkC2PG/LmfT0Ke+zAUBU0dFvFhITGpyUiu9D4ILRilXEF
mf6CStt6NhkX8gYoHAPzhf8dIER/+vhhljdc3vmAxX7o50IMNke/h4zt/+54Yj0Y
n+9GLQJmeO7CjZeU2CgdO3p2zZHxqnOzyF695UI/pSPcC/7F3AjiKAUr9Z2I6kCa
DK7q3uNJ770RqFdaOoeeT1aH5UcCfjKAnkohy4yGgxje34/GQz7lTHJCEJmMaQiE
4uM/M8mMAyH/22CUA9yxyPmqFDV+D7cf8205RA17gRYdXfu3+2VeKFVPl3H+4gjz
1HAXWv5kf3N4sVMwq9cdx9GVHGRT+SmNK0nMD4ZKdEpzA4jXoALvqLZS8eym5rVi
9raGNkEcXGtAX/kgMK0NHVRnkfK8IY2X/AfNsvOQX5dhgiW9qD39/EYIcDAd4zwN
Kre5HJ0JJkogIVb/X6PlO6506k4L6jm5ivMsowB78uGelDqe2j9LQ8HpobQlaNQp
rOrQvEHp1GCkOsMrWSjwhHoOzR+l7NHwr1i6A9uDPd3wZYKj409vkwqZLu5Kz+nq
b76dY89a+u7hm2j7yt47Og+x7lGKBWNbqadilGLbA9gSF9MZP4sshIgMIsnoxT6N
acxrTEdc1cqFVXUSAMPP7qi9GfrJYdET5EBVf1VUOcPCSoHrEDbN7tc1m7DK0cpv
8J6ZTZ4M2gZk3uVjIlHJYNdKa2IdrKIf//MNoBVA+jMDSR2OTZadctNK3DG7ZFGB
1Pa8iPzVHYra24LRnYNhg/oxyAlYpAaKX8/EwymU+8RFHzmd+9/Eo+opXi+w+ugV
xTTryamPMRv8oSm670Et+Xfil4nWVgbe4dI0Tqrua+/ioCAIXuBAozzVOuS+Wqam
TZI91hPFrJBfoV8wxDAui2EC2bg2QURFcQ4CGkgkiADmOSEbUAFVjQeV8vi5k5x4
L1GNqnkR/Qn5Bm+mWC+R/b+mTMOqLzvsS+j/BtWFnySrtCZbOZaYJ4wyEQQFCCdY
ysXC3RZjnI8lSehdwESeQo73vrYSzC/k4vO+AX0WwGLCBm7P/fd8+9jTmp0oiC9O
mt5H0RaJbSnwOBBulqbOjR15hy3N6wVAvodmraXB3vd6PQAMSJqvRu+aEEYrGxad
VsWZLkgCeauDPblwOLjwR14ed39o0/RzjNhMdLw3+1/Rf7kA+FlD7BYTcYXlsefV
dbD6Oz5gWJuuaub4bXrlDr+adgxmzeluJLjAFRfTvgvF8vacRtshTaNsL2t49CD+
X4hsWk8q00hE3z4bhC79ULrfUogoyTZ613wf+NTNjEFg5vnTGhnCGCVUXxNPBRtX
TmlinmFPnl9KsCJn71UUMrJVyndW3vIY2+tQEGxr8oRxTGgHIv3xu7NzD/hymAZ1
zdFswRhOsi2TGkg+g++hKgGBZ/y2smQjSaMVgKB5jUDT10MXTquz56sEOy2mjbMv
pIPUhVCziX4KtR3jrilyBdkg18pOYHB4VaJ48W+pju3u7+OHgyxzcmbq0OSQ5lnQ
gd76FKF0/5RIXA1ihOpB6o8h+nhS8v2SLd2MSB88tLmSCodaXKhB8IJ6b/x1LHbp
MKmgG8n21LKZuCSmaWMp2vTq2vFuF4vWEd+xiQTeyKa9Ysyq0r8RJT3bfHeuWKeJ
trbM+CDRyOGoUTp2Y8vxP1pLfy7TTrlDe/0WegYeaFygBW/D+MQEMMTJ3z76Ih52
tWZfo6WqC4WEAUiYihNHXCuO5M2JN5tKtG+C6x18TogR8DtuEgUB42z2xB+UQcqv
6N1z4tjAfXfbeZtMWWniMMeWNdOXyX7YHbtZAIjFs6TEXLZ3kskt+ul2tgFdPEci
SzcnAgeIQo+WrJlVHruEKPgtB0xYZsvYfKxy75s/dTKIq7/ACboUH2eH23sSz3qr
SXL9vICkr9twzsCIw0x9heGrjueB0ZH3Zmd66nY92Cpn99sQ8SzaIOjcbPfNfjjF
uhMT6pqVoMJ3CA23/twawJGsfLs0+a6GqUWvgwM8Ozms1hXL0VkWzCyI5ioC//Nj
qPjwmUOxwT6NGcxzCucCE6vezhG8b2klqgz5oI+BQoJpvK4Mvpc3yA82EPLUhDjp
FvuQ3L1/eV2CHhv1Hp62J2pLf5q5eLWctndOe/MN7c422lZG0DFXXugETpf9J8z2
bXNS6wrYWwi5ZaApUeKSl0wcvj/Vj7M7oYrD7AtQmaLZq86Mea9UT/LsaOo5mBPR
JFK/SBJFRho5I7poog43ipV7X/onY6fIOYGrByINq8v7DVKP3ASw+oN4+ctpzQSP
fK99GXrEB85pKXhGXAUSXYjA4TG4o64P9UbCi9+uLf7I0YJ0zUw1T/MT78Afkvtu
qhkDbkhoi3/+54uVRMTyazkimnwCCuY++5br9L/tm4+W6SnuT5qJIGoERj3Q0/Xd
4mMOXog3y4AtsSsnUR4GxItwjBWcNxznF/D5Y2odATmZaQhJ9kdAeKZVOSMCUdP8
/QI7C0L9cnp2JtSovo5OBMk34a11E0BHdL0Up1Ueo+4uwVcwgn3PelPfUNV78MRf
97q8KacSZzxqwoc7fonLKTAw8LsYas9RDdL799LH6lrHHBjseHZiidjhXElx+HeD
KfdxCZkCyPvOTdiqE9CrA5ZpWhM+HlIMcO7IqML4PFKHSWKxMmIicCbUGZtRPoq0
5oUUaNuWdP6R5rm4ymHeH3n1ZIUcQC2vnz2zEtsx4Zxn4Gts8ABdw8LcSfVWyDZW
J9+2fD48wL/rBY1NmkkFfMmwtEM1oXFlQrBjfZxtR8vqmIzM+gdkKWCKxfLkhJF5
Na8eeJuGw1tP7ylePXWy5JzIhabNtfV7CerTvhiIGrE0Q5ypAnJM48tLOvhdK4/G
55YBqoDapDJp/MMDacUkoxHF7mI3+1U865pigkd3uKG8tRsbQp7UsvLuZ0CjOGgL
UxISBbUOcvMzOEDWQlEVdVHR3uNAbUCWSd2Po2xM+5OOIeiJ961vzUtAwDPPvnp5
ttw3fihpcHvitNEwkNjquG8LI6C9SsiOBZEJpySkll8Xh0QA/HYjuOD9CuPVVguJ
IZ4+MBxhQF4/QeiyYloqoWosxCv9GMZ0ThISmvm339YOBAzjSztUlACJgrnMXneI
1DOf7c9SU9Jo1LADe9vK3LQ1sAODcBZKckBrHOCt/hW0xUUmN7E3ttDhrdjlWs4x
RaD+kZSF7/yDTE7yNMdar2XRHr4XD2hcOF24s3WqbV15n0sR8eiTCHsPc33lXlwO
jr9t+GFhGFvJfJyisIWHnYx00hcGDGI74pgFRyG4+tap+ur7o5YT6+gu4VUxlNjL
9hSBygprbiYVaAAHQvlQjxC1u4U6UvnSv1ZTuQA+/whNOhTbB+cF+ZIbiYcC0TKv
0eMLIxNVcVVsgL6IP4KtQbBvuDn7yrEbapbQLvDKRQHCn4UFc0CkXtFgTUyNs8nD
n33CHBulcf3tyQgZJoq/wznx8CUZCHwhBivM9ONZILMykOHM3RFuPkB1IhZgZHMQ
uXZSRpfYue51ktQsY9SjohcYuuQi/WVjinVyW6xTd7mmCOCqI9K5m+yL5r4kJY9h
eUDC1JqnWq3pDCH0h6oZOcU8ggu3baqzl2GBXqRCkzzwfhK58Ly4RaIp9TvPmkIx
XgGh73bmaZ4J13S1Zf330yePgVRPQoveWyfMMVa2Lawb8Ma/DSDBZbIvzwZoZiEo
sesyaZfTaJ5hb2KQu77j+dGmGH44lPMOtNayyoQmigt7GOSo+VcHntWwbkEcDsnH
bW6JPTx06FkH/dXOPh2g1Awdx/mCPvglMdVVY9zU6z4zD03MCx8v9GNTkO36oxWK
OMaw+IRrFo2mo0cj28luo6DsxVPhAPEnBeS+mm4Q3+Zd9qxBV30u/2ZnMM1Y4qun
gFYDbVFiSrTG7/X8b5kD179CDl8LVc/kIlAl4yANJnUdJwPfcenSms0/Tn3jUuau
E69mJ1GK1Z8GOWmCJfRtxGGyXYAno2UZxstcaWz9iVyF1HFpcW71ihCJJwRfTOrW
wUAdd/zshRVk0ZA+cNn+6/CFbkxqRSUa9KOwUcQcG+wkF0sHRrqB4bDy7o8n50du
nI8deO11BOeTIFsnsCuwulZC6fozXdN7Btm90Ipzmvh/F7xGrLF7CCBdaofznodT
M9QXmfuWMMa6i2fISDaO9VA+wf0texmBo2JoMcrqHqLyoziU8FwjSE4Ib8yERFSL
1t0Y9x3XVEDKtQK9ivwAZJIDmnn/ytgoD8c/GySYVFdMGMkkqRe3ydzZQPNiZz+h
s6I5qSKH0J6asUVAZeT58tyxERfd6uqkWkoVMmUS2HCUZdF0hP9EWOySpgGMRQDT
QnhwewylgHZRvFCxqVhIx+v/srTy+aquFNJOUmj7ra4gYUtNrmA56e8NLrS1oh8d
tsUdkipW+Ba5Nq0N+fVD0Ic1U99mvM9of8+t0Ml6QDGj7Lv/xBxYSNeyuwDRHnaC
i5q2U1CyRuuyHTsvjkIjBf9kk91S7QqwWT3Lm3YYoopDlekc9IgQUOPizYI0olV6
QCFkKj1aosgFTe/tak5JTc4BDki/xhLnGn9Y+pyMK67pd96r3ioU3N0kSPmTZgB7
dfvmLhx8rv4yONwXzNfa5s0vU/AdgB3GTzYIGYVrosQtrxvybJc9dozbi1bNzDLP
GKPNalcxkSzhschdsNgWRAsakNStGvzv6GHE4Kzxojq/gA9/sp8ZrKOGdOIxPIXu
z5rzU7WejwWVUhEi/OklXIXdwaxFzIGhx1bxuqHxdsiYw/0N9l7yyXDxlovHLHt3
EaZUA/1Bnt31pIbvuXKhOP7yStzbh5krpHxfeFRjOHTJhhLX08WD3hN0wdC+TP2V
UdlM4IA0861SQCSXKieGGuJIG8/3OQ9Je0usvki+u51jyyCKd8F5QWmuIc3sTebx
Kz9peVROZSBpnFW83tD+vyViPpEh2tQIUaY75vXb0r8Ydjn4OXAeSWPIFK+Sy0sQ
r1GlTIr6tXNfs5CLCuJFFw5NvDSW0qsSzPL5y9wEFkUHpQSGxtVIyV7MOQS5sDrN
IZWvnxEoXvXLMKV5R614kM1uTnPbUAUz1ioNwTj9oap/rXvkukp1I1A2coRZC/Ou
WZcXSdPvlB/ddEKUckSTlExYLd+w6407dBzv7o+FIDA+DawU98VEkmI6Fae7A4BW
SP7a61a1hFTGl9jLgPHdScnISiRz46MU1YzPa0BYREcQl70JqNp7UzE1+IzeJzyH
5o20bmeYUw8ii2ecBX3rWhxqVgiAtTyu8czqlpoxJZpGmCev197ph3optrUDj8sW
EUJdf758Rgw5+sfg52njPSE/FXZdtFry1NX3VSBb5TIpzmJVHwQiYpYHU3VMIbEm
LsTGiryc2ki6nnMSXOudC+uJa7XgeVEbv+DlrTYG/ji6G8dA+GDgVB7ICbA256hi
hzrr23lQNdEzLEXT3Zmt4rYjPTIhM59Kfr1rFl2HR45u1m7ji5ngUZgNueEsFVtK
gm2m4KjvFwj9DtjIVtcTB758uJriyXWhWe9VBU7PgY1+IRjvAcdMv/Cr11J10W06
VkGl13PH/rC5lfNaZK4v7zBS51j7XItL1IM+g/PJ/hrHltfb/kqT19lbbRWn2IQt
XLXNgbUb24iNLlbErXaDyfcrms8XASx+J3BqZsTgdEMJYt96bFBslvGE13w1eVW/
Yj+drRl0IY/mff614EgaejQgUtur2DDN3qO8vzlr039FYOPaOb+OBXXkUc7XKpe7
zzuwgPGXQ2sGHqVobySIW/BW0W+gMj9D1zoorZ4RUwPBv96hvNzi2W2RDW3RPL7h
mDVIcJdzPWyokhu9g/sRrBHBR756wykt7xyrC9sb5JkPWS3kaTTvtGJ9uFBAAzl6
Sm+OtXzRVjvYpwgV91KGUzKyrGzkfWv1RhNzjHB21yO5m/9wavVxeRAMuKlolgx1
XGGH8962gSGnEPnwhCwRBhysBKhl2WooKeWFTGZiVFaF3xGJJrsM+bV8Nr3Vu0bE
TcwVAWswvZ8gfItP9pRQ+HbrB51nRi/MKhF82q9rZ76sdv7QciE4gkfkSbEctsdb
WoI1YWuDHPcIgjddNdK5ZGPZkuc7IGRmx5kygc8qvTQriLNqz0pmzl3vxUgTv01+
hdWVE3JkMUMs8ebviPWYoJEPhpRbA12Eqk2BMOQkJlY7bWe0YCJgSCYLltKNjcir
2JlJYUkrbjqI9JPh5N78FYqv3Rwa/3YkzuukyGbqHMpKHhVjfAjlkAlVVymdqQkC
0ksrOIwE1Mn1zsDHhCmybIAx7tHhXFMyJ3cie4UHuVFMPet9r2Ew4TcBJ++oNMW2
bnuQihsSGuVMBe8YhbB+IgwwScCHIMyfpUwNCFVaKvH+WePkJ2tnH0wOynfF422q
MMP5piK3pjLTF/QghVKywKpKUZK+08JO75LBdBRTJ6TexHTswti6w4GXGpemzshp
kgm/fG6Hc1vYg2+TvwknrlGhEd8G/nVodP9uoqGhSTfbQpnhUoeDh+P0KG9Y7PoG
FEkP3m5QB89R5yoNp20Uf7HCOJl5i3ba65ztS4dEp/RfSjrcbzpDcIatE8ldPrlu
j0Rx0nwf7gCkqKXAeU5I3lf0eEhcAcuSOGaqHRMpuvByzVeNOiYXm/HOW81iNX2L
XxmtvytG83PV6sZ1hLp0QajiTOmpC4U4seG0CtnPhrIEGyEDeb5UJYg07xQ7m+Ie
rO8Vn9UmyY5FACGeNJKjO1gfoLioYHEk9SljVFwF/MaE1aAZDHFQdbtY14Uk/VKj
VhYGuPjgXUCkBms2brh2A9HfwhFk4N9LiAzup7pFczol+Uo2bpI6Ax0H4T4i98EC
oY7Bc3LzyQ9xTdOmZAs21RWqC+S26CHd34UkdlFAuzbjTCeqXjsxEfXnoRG+9b5o
L5QyWYcsA1GT/Q3WZZL6gjR3Mty200Bc19iXqf+xRS21ZAyjLs+XwtSj8mr7EPZI
Ol7FqSF0WcqAyOnQtx0Oo0zORZQqTHDlzal3jWE1OKntPsDj1/LDK1RIzqXWiISU
Xc08RvqtEI+oCUrymwR9QxoBMKXzfUiKsWTaqGzaZeDfXk8TdCqxcS1L+lyLyqR0
AZihkp9vFF23dNy5zPZcLBFlYYI3/eD/GDfpvd2kQ+322JqXvku7yVt7dS+tpVBD
93Qukzj4I50jBXwr6S+ZYDZ2fMvF6FWlSE0xF0M3iRnph9HPl1HwguC1nfGKGQzg
/eyVcNSY+3KGeohvuHhjn+BTkmZCQCSZ6HElfqh36hBIkrY8/FHa2qAwTPBKg5Xv
lkxzTomtl39VIMhX+DpzGMG3hReZ7hv/SkJN11tzUHGyr4Zti25jOq8nX/cBflmx
+lhy3lcps4h539IpCDbQj4POyFWpS3vHyxaA3bvVZsk3GxE1m6NAWLGhMDBbOPsu
LgA6UNEiQ7zNAl61BhOtfBYrM4Sy9AfbaBAYEOvF5JsY8dpGpELkYPM1Mvv2Orgh
B5JQJdaaBHKwhSHqeDBmYOGs+WTdTZq2E6Oz5usVYL8lXtItHdRc43ZabpWJshZG
k6GeBtcydL86Qpfck4XIAOBEAXcysVsLfoirdbQsXbojUJIInVDbcsyeFamfwuUt
bZBvqDqT9oaRt8wc0yeCgc00zOVRGMTOz3dsc4fa5yPdF/T8kYCVt2IpvHFPkvoF
yzzw1GlSqj9ltFyJI3uUSfGP7edqNHFLWRUQy3+L/JZv5GeQXZXVTpQBGS6u2Snc
tiTiieoPmzZbAufm8Gppv7+engA9lNfgcKxYPG74HJGFIOvwB/CC58baI9mmUKwF
BT2hMnlB2LfjdXLlSd4BmSY1uaQgYnHmtLbH/h6iDc4wJHwbfeKw40+7sx2NcE4n
xXr/T9AO/j3Qk0x9E6IS4p45u6B7n035qX433WD4qfhH34YJWsTDc7Ll2XTIz+xT
eNaAXptdf+jP79Cysd1lkMoby7DOvurCIc2CILB9ILEAkbHM3cL88+sayNbncgUZ
q+RC37reAF/M0SYyL9u7I7rwW6ibG600z5XXZhFaoWW0hTu6aMDAMMBrMdhNWPm6
DWEp4nVOSn1HulHYjsxoNpuqY8Iv9tEQONdoNy/mKr11Kro9gmbeMZ4GZX04lUll
TdH3lBJPr2WHgeXUEQ0W6bhNFJV4rOTXi/6AMqC0pSGCY3hTdzJUIpNPFuMDgNz9
hfpD4vm57lW8uPo+UsEEb1qpXRESZhJnj/Vqi7hDWT8nNvTRDMnzXKX0cvTCgCOM
+L8sT4Wld/IzhErAQuyLEHaldM/mKn6kjFP5xG0Og52jcecv84KWyP8chKhv42PE
rLA6OoopyAO239lLxOiLJPS3oDurXCrVI+93+s5UESO7a7gzy5652RZfbOZuTFRC
3yHF4YWpYtXpLAYtiT4qGAPZLH00IMP/pc+QHHhqlzVkKoCHmCztseNwo+enRv6I
Sdk2EmtPSSCOnkSjymu5/SIPrrA8DOlQ1qburgrrRdN5K8WHSt1EpoA4aSIJSWia
ple12e1NVLEXqIcfyB/C82dceHKuNNYLIdP5TdPCJGYpK1OGxkmUO5dIKP3hSMV/
pzNQqKAquIAEyVt8NuyH8md6fN1KolAMbjjqCTDHWdroztK05XU8n6Qpp3HYED47
4Y42Kq7KgbfpObsNAcJmTvJJ9/QLgb8FZ3PKuDAt6lN/uzh2XMEx/pr1QSnrZ0yq
EpqxuXlaLDu05XearcqXGMjC5jC+arB4KSRphMa/k0rYPuSHo1H+JCOyEHgakXov
+3/Vk20NcNyZbgcqg6UVt5dvVOC+iI1qzPlvF5WOZ0MCJYdV0Eqxj2xs3QBl6Ij0
dyfW72Y6bLxbb2TkWMkf/pRQUzeL1tBiZC8l/2votvUsY7/ih5nD8yAMmjDtlAs7
uWybwhk+OOrNvOzw5/40bWMBVwYV0R3LRMLX/aDEm6eNZquC4XWTY5i562Vlw120
IIln20C/KE0JoNbUanJxvkSZpiM1tPJvbWyFtmW6vKlkobKB8CnjjMbjnzZ9ck24
GX+pXKtlZqWmYefhHUivUfaY5nDsmIyrKritOO90ISt0/v54/QRwLjgai7Y9q82v
lImEXft6ocm0pSlHLc4Q2KWRzcRq6eZChZMoHpIw+YCeJR80NQ2kYotmoYYYBxSk
nKUms1KktLPdWFw5gZDix9mT8esu8NzcN2JP/cC5OoCc5sWYOSrRQ2MvgP+a7juh
gT7Ru29VWpwbrYd1g+hJFPdkrah4sYFe8BsSv/ttZbrVJxU8pd1PcscngYbhWUXq
oFY7P7Tj/BL7qPIc1uBhEv9NaO0+o7HfJQFCPmvpw/6Q6Y9+1GwYE8JYHcme7AOV
8KUuXcnrQ3ILGs+PXciH8Z2igJ5wUENI90N8jWjKfVA7ddqy6SX4KbxdCe6YCPbN
geH/xYfObO2IwPL6tmQxgkXYrGYj7q8lUFEFSRBMCZeMKtB+SOokWCnimpkzth2y
5CU43YhbEMQGCPsGesmmmvzi8U4Tfbdc2Wv6E0uAS4cjgpnkqMLvDLywA+Q/3JPM
`protect end_protected