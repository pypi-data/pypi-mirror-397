`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQMy0Nic0oPYTT1PeBRgvHfGgzllV7bXuEaGrj1yWjvma
ZkcszlwH7PEfOxhPWGxO/rNwDasdjkuQx0SlC8+cuS+ZQdMeSqldu8PD3Y/mM3/F
mUHqM1ma7FxMw/lb+voP2aI528qpnGGd8Vnm4bOM2BbRPW+MOO0O1IwJv/5GkDK5
gUINj4FYUn/gug3lfqKC6aBMGALp02lFDEJqb3oJSuG7br2wS6XtGjKqWGA6U8hq
rswJ5VyQ04v9Kq6MlyLB6a/7OKbNy9rmJAX/Sc8e2JIfk2NtCKbhB9ZcNdkMzTUl
lQI7D67yCUALN72x9ZDJ9XPfBdi05/9MO6I2wdaxhYne1E4mLWIOkSz0+2tVVbY1
SD9QiwnLLz4CLALV2Azi52roqfhzFJEhnQE7aIuk4yVMtoN0PSjVQ6CoPXgLQ5Lk
r29N8CXqmI6Rb/QWHNVfdmAUhZBT34KiZlrmjCaVKXnsOPMXXDGnKe76ZZdYac1s
NbzS5wV9HRsNms7cvrJOfrmREcxc6HmmLOLLrv1rHddJSypag/GfrvePWu83R1ci
R3dFcBcwQNJWIutEZ0EwDdVnKKUdtdQb+0fcKpWGwl3GI8OndNEWev8zCqdFfppQ
XUhX368DdkTlSFeH6RYqYbJtF/bd28+vIjLdhsnGW8vM1xgqFaKIVNdEGIXYc8KM
zGanmsthHqAh7Lexi5Kb36SdSeKf/09kpQ/2g5BA65aJ6SnAQOINNQkNGgPOx0aC
h2DFrSQ2oK7frMptSYcFmptHFPnmQXb71h6U25qRUJDrW74TqXw+3vLx86KJqh5J
Njvhj7jUuWbFzxUTnJRftybPAwtkVkYrkCtj35+QRGjnTPwelLN4t5vuOyQ82Xss
GyzaifzQe6MdvD/ZOPwFYDNRi4cZdgvZ8mSBBhKU+NvqrB9wVszJyHDTyENV2gJl
W2cxgm9AhcC+6JfrgyiH26wLnCWTs+xcxkN/uKWiaTlrKzlTdS0jHFcTos+GaqpN
SnWsPy6IA82OMRhjkLrIM3Gb41JscRekE5BXb0xsie6aP4T7DnJM7X19/rVOoJWR
nmzt1LpZzov26DksT+NIQULSglDY9nuxNhLsz3qDhNz+rSNP0/ys4hciRwbYELZ+
bTB9HYrMlfS10Rn5W7rHEdKvxhbI9fbqxc2QC3NTTH2N4Noc5xDcOXkJom4wrA+a
xTPy5kybH7WZaQI1pf0gxQVYiQUaCvbvoKVjl5GevSkHwCSRk0J3gGJN9VGDOtRc
xgckGBjezHWBAXHB8P6YByRZTCSsraorm3eGNkuT4xCxhR84owozV1tnWP8Iqlg+
hN8vip7tb2kZfkVf55wiRHhaHOUQW+eCzU+l6lr4j6lT8y8bnLM0Pz46sBxf3ls3
BMD2H5tCMsVYRblcIVbuk2RCWdXo+weIIwNpWfYwvIBN4qh6NB7yZ/x16NUy9BJ2
df9Hw9UsKUgRJ3M+Rf/piW/Ev3M2KEd5CuvA/+qUCkHbSaxcGtQsNxHTRAFSCb5J
+TOiQs4OP4F9fiBAnp/ZaDcl5/OUa3dLJjdnhtA46MAWOaIQrz9brhwQeZUzgoBj
iW3qs0mHOl7cr2C5CXeOXgJdUPde0orz1nhxDIDI0WYIjqhdTf/Epo7L9ON1YwcZ
wUyHOdbfjWexedGi8vExCjlUrKw7OIPuP6nGbq6MMA+u9wdo4S1CHZYN7NXOJeKv
9wdCNdObkT6L1Q0J5XvVTIjlr0b0XITxtXEsNRCoBj77Vm18Gkr5MYa9sstIU8SF
0YWpHHyS87697IkJj6C0lEScdFMLOXL3aSPp75zfW+divO6UkwTsrqpiGWB+QaMO
a12gCTo73daWxAw7Tzqtuu44iU0sBnr4RxiBdw2/C+7B+D3qLAH/MvLXnuRXqfle
s642jJ7lE4FGIx0YkoGfJCR7pPgSmzRTusiHe54VkQttj/pXOdGH2eUDHq/Dwite
8bHEPvj3ueTGhWOdXKzszVB/HsJvlgRoZkBM8TiCJMCE377wqx9AE/B75tkE6m5G
0mwpH9a1uz7zVrKm3dlSn9sVuiDXtDo2eYxXiOuCo9sx3YHv2mN91D76mo3smSRd
goOqBDBM4kNRONf6trL4WMH/o9XJA+eOKftTLGIyYqJZhp/FV9Vc7X6r//IcAkvP
tHR6H3R+12g8ogzSWsIDKRjRS8izJdnZMyzqeej8xEhPpKXGx4zwRgzEyAUjWoOo
fHQsxcvXB2hF3MXMZhOXd1rTltn1WPxNcJgMYPTZ2QNS/Iu73DtbG+S+70SoNkwH
uTd+2DdYe8Z44sAHkANrHuHfPcZqYa9WmD0p1focEqzi0xoCnKocwH9r9DHfciGh
AN+BiVIgPcOSLqZyW/KxvPiYVqEN7JxsFhtf2TpHOhS482JvOWSSn267EMfb9PAg
4StobUKHbnMqmF+/evuAGmAiwHmex3xPReFMtDARXkJvVYYsIewvVhruRS/p/a4q
PzdWXp8BFUc3A+OAuabI2jUcBsQq+mgQqSCZtRwxGKtl0EBCKjpUySrlXkMR5iPg
/NRCu/yp881xMQ3XxbQ/YZYGC/EnIYULVLTIL51lhjeWiJ0kwmzErhNlvYEeWFbj
At2pIMI6DM53F8WcJIG2YmSXB0hYKLKrVcGRYYo4uTtdzsqlDgElwhvlw0oJSYPx
b5f0ON8kTem/HlbeWmf/B3ypWSX9MD+Um0wr+jcGUR/DvAfJQwuMs/xCYJIKAO8A
rB8rjW0sOYpbEE1Qk8rvVfsmb/XWtkXfm0YyulpRHTHn+7HJ2TAt+6Auc5RagYK6
+gFHOWj0TSCiGveUY+O2oz7eelnKtllj8i9JcjE4Tbb92g0qs3uPn9vdw5MDhsfg
pUpy/C1Q3PnqqIzlRMCDpfTDZiRUMha33j5NOMZr5zbjFCbzr1J7iap0AsOH+iXJ
27ZUInvf7guyYFonhzmc2tRAf7Xjow32aJOcKN5XPSr/glExQUIJetdbxAGJuePd
zYXxairbLESpy2o7CHa8Ep+SN1uXIL+Q+rmjFFQNowhYKzU2AplnydNeILiy2yRY
xPUuhjT4eUv+FiaNuWL7xqlK7hpnOvXVTjfk0Gh23RBdO9yA9/4i1aklQ8y4pArq
CdNrXP6SZgb3XgiAdOhUJ0DycC0gvzHyG9mYV5WiSnLS5wRK+bVH2CqxyLwd0IJ2
40JBjkZQ7jBRdvUkxAZ0BaCuhn3MTqwNOl2yivyue0r48o62bpi47lLg3QZ6Rk8v
+93F0fvmqR1RScXvPca0mcAG31icM78AvjTQIe95Tk4xMz2uVtSuAT0oRBp9APA6
IMm6q4qzVBBf4JDJ6T2nyiys+FLNHFD5YVhzD1Fkm/iN7uq8mE3X3OnC8Xo5Rf/I
VE7+qORbpS2CQXd4rFKhB+brMY5Wvsx8NAj3gK3z8Ft41P0q9pVgJfqTOUFs5K7O
lZ9B9YTBIFyrLgUyp/YrHwfOSVXO06IfDzBCpQK+bR//s7MmHWNXzSZK7xv/eRA3
YAb8vBM+APFu+KBASP1Yc8Ps9Jpk2jUNTqTNO010LSgM587I7gxXPgI6jxSPIc7n
bQtNqIWbxkXptcVts01a7jovt1pE5u4SkTcdFACBdEPOk/7scWPFkvagWT5p/MGh
ii4t6j7IoDBuvi4z3Vvoe0Rn6Iaob/tRa7DVlQkBznJyGaiF3dP8rTui7NoFnc0H
CbRPE0wAxkpvIydyrCXUhqXBwE81rUZbwIWj/QVgQLPYCl/hq/Z1F3LYbXRTB5JU
yzChI91bb4mXK0Ec3SD4ZjqaT8dswbFGXzDmO1AxfZqA4eKoaLHOMowzuHcem0wN
gsKhhKRi2op/Qa71nlu1NWu74f8teJBKrArZ8MGRPi9cUgbbbbLPENc9Jif+1akv
c/zSD5yNUk9lyEHoLSNRyNwB7KYfRMl5t1ZvRTnIPjj2LQy2GP21DBLpdLEKN2N+
f2hpDKpMoWjv1YNg1KZVr75pSc6hegF1tsUpZ4/RNIEGeLsrt9P2JKmZCB3Az+GT
V7e2baUG/htSw7p7n5hIMlkvSwD5sU4/8x86IbwJ/a6mibcbtZ5F2Pf29zke2DnB
rSfEiO/vawvb/mS/h/p8NylId2DQH+oXB27QuIuDqzxoNmumdYo6vdSNXHxNbYEB
ijmuBRSqqhuBpoaXDmro5W7OOXL5dlmXTZg+vD8H/N8kF5QmlIXzLaj+iJXKUm94
t0guO8aMuGYCRiIevq4NXFKHc0QHT70UcymBi53NVes6C3d+CpzkxCsrdzYdJPnh
+OwGreOuHgm9SC0kW1jQUqurG8nraYAMtGkSp+8Frxm32229VPi7T7fwomUWk56t
8YECzRsUNR1TTMebAGyYiVyu+Sv5AQEed2QEhVxa7DlQtIRLGkBzGsV6vALxLJ+l
M0JaW0qSDi/MWViQMW5He34VfCEwve+5NcW7mAFvvaVk7qWd4wkMd3Fm11lLCE6H
7bBaBnwyylEq4JJ5WUR1we57SgxBLQmOpW8NRxt1v5S2OPxepPC+PPo5V6coz7WV
DKMHCNl8X0Uqh1QCUCa7nOae4bAsx+dsovuj1W37odwsmWIoJTeWmcj8lZmuLGRJ
45q1AUlSFgshNeXFh/AJrgXX5pzsvTKMFM6kvRMtu1LfuKqcVknEGvNx/cV6wThd
FYmgCHO6QRJYbWzRVMIcLdkXZY3YrrhH9GFJU21mnpEt0nNtjYPlmi7LxflK/zT3
FpfkKH7rGnzzjzZDtrxyLfaqGQtYiY17FRAwagHqJFs2IjQId8Gdhh8o3RuN9wkq
moHi9SM/Qaj205LVsALct96zb8rq6aHT71lmLYHuoAoyyx60cGSm8V/wsbSxhp5e
qHkQsI8ShegLY7+ybyA2vn0UiEPVTzG4mzOBWmL8+TZmltzSY3HWn2dF2UBfT2EM
7mP2JUEti8u3zXYT4p9X99eyFOpSbDUZ4oN6BKzDDaNLKxGt1uXszk9ZrgiiPANI
xHxwQ4sWzzUhtDxJt2vweA9d/Z2vEDYb0l6ZVLqOQVEN+jELnw9mXM5j5qTFvNuK
nf18OuAZsTSwO57UjI3XQVN3ZXPy41XBBUKt72SgyvqlpDv5lprSQflNsN3V72eu
fF3ZdSKB2PO+P/jZ6uYef1O7AHqoa/aXX3Ijf+VPFzNZbrAFtcvis4BrMbDWB8dl
de88a48U6OGdrHHirImfKKNo8JvRZjs2cScgVtP568qOU3BxmnC0A3wbDpcjIzHI
Zgw/0fSKmFuRGtcii7l6SoLXHdJen76GtqMFW9qcpKjpsdWbgrJzcDSmj0VJZLvp
I3LL8lRa0MTISitsTECzRdupq44WW8zO3k3UP+4yqmttILBv5TTcu77mgEev5ksI
0qGKHURFySnKoE9hrL68BSh59bxPgBRuCz6w6avCozHFaUZkzVsk7gmbnvkIJ705
p4IQZo5/wpEDR/Ehn0coAIwlexZlmQu9og6lnLjxZR0cDpqRHQo2x0dFjSDGL2Mg
2TjJLb3lH3UmW/JiXnDpZwADTfyfrzE1eybo63nKKUW983ISaPRUOK1M657w011e
7QkeXPU82mhD9ua58sCqWei6aR07mcRHR6B7jnL8gorwiuOmKBecXF+t9vMtIeng
4weXCiKLJwpQyItppm3SiOYnOprTO9KTlOpenruKecneMuDrig83cV340YiCC8Vn
Wv41aL8WMUSM6fL+K59EJtHdvuPT4VrMU3Up5Ip2sPxP5PYWVZQ29w/uSi4ta408
NR7mSm1svTKio9wVuAFganbVlH/KI47tasdulX782CSGXGQNdG5R/aZZOqLgfzKn
r46Dkxn46+l9+IXM6oHQ077ovNeM3BHAIhxAbiXVgBHO6lPDOfx9yhK21PItlY9v
U5lXNmtAUKoaMpUGgNVn0duaLiTxKyvc2SzxlXFuu/QNcbxflDbGqaxiKLmCxnes
tTQ6MCq6yE69lu8Qi8RAr0G8qXENgscbcU+iV7J1W8fRz3ZjBFMf/wLm4xzwLRaE
NKOoyWTQ8iFMCdzVT5DgKUAJhgNyyMGvb5L+6FLnmbWophegJgtTXU5A6iI2bEG1
XDm+Fnu+U2OoB1I2geEKThlpvwBm12j7YUxgBtbQiiR3b3lPg8gMdZM1sljCaV/N
tnHZlOWq/BVLkrvhOgjvbCvHVObNZkGpds/djdrBkWsuWKea2P8U5I0AxEQ6NRbm
XREeV/oxPAGjMMf0pVkXS5xFK7J0/aB2qeQAPJZTzhgayG5d51SK3mYr9uh0TFEv
HB/qvsBSsiYVWXA0Al7gvohCS3hsRJlkEnwnoUPf2yoXpt9uVEmpFmHKIuFyKoeG
TDI9zmRIsvqTyAbFBDu4iiOxD1kg9bmzhVO4h0THGJWzRrVM5nOUyTxuUhrnev/Y
z8LWrfX1rzX/uA7kiRgXcr1yxd6mz8B90FQAWbnVANnbTbU3B/KLQ5MXqZ3NxDXF
TnGNzosjy2DVpQoqyvDVteMaCx7HCd8E1256LvrpqG5p2GHsRmLwRWT9+rGU8gc2
Pt7Go0rdLhRrdwPO5GwrtyOGZpaa2S45uZz3hciIWoVmsYDrfQ4sttqxr3nPdu1P
GeqbuXJP83gDFd3xMSwVlg5J72ucJXOcmnH5ofyMN5W0a1+KWuePE+sJunAXkuwe
OM2g3E1TOMglz5kANRi/Xi2qRz/39BSqtGFbFkUyRqW3rI2QPUf4NJwtZEFPuRwg
1XgIqRFucPDiDVT8R18Ql9Cqg/mHHNx8AKM8XwdlMAlLIuaKyitfVat/Bv6K7szx
VgvNmwUflNitOofsOuFjSlCwJaYfTUAjwZ6ruAJ0ySSe8iCCYNYNaBOggrrcZHKU
6EOThOcES8z4F1GcxTkYFpfeLNePvktSlkiGyLTncXgeTnEaF1ihD0sVkJXwcZJ9
UkabwmVPx/ZAc5+1TJM3zY4Q9wvUkYlbbAoEuzT9/iC/UyMC/U8W6kRQGYxgeBYS
G3nDKxA+t5Lf+/sItcZUEpzhdXp1R8wOlXjHZljUmqGpMRC7KeiBNJE4wXQe5Cni
QMXUADBzgr3QUVZM6OFpaQ3cViQ6IwQjaKc1MhbjTARvdvv6yzVCakNmjG5ka4GC
yHxz/hmENMIVVx68x7DpBwJSr51pDRjPg3LfJCEEbRHFuKuT7YDxSeG/XWhcyowF
deCkKSNeSnG8ZaxEuhRdTp7lDGkMB1Ha+0CdpCXryH63KlJa7Z7cDpqGBKaZ9BjD
1TTW0UQNws6kW1GpzKvbYDO84DE2LfVrF4hHFS4fK0KVI0s017vYlaq3bDKKWL/c
RPAeN/qTg95+tLKfjqGdyhpz1GeEF7ihw7CvL770IOyM794vHWhieyet0x08Gq2F
H/djdIN5458GKe7r1jWPQdjt1qOd7d8uhq4xJXCeWzfPsro4zWyQ07vM7Z4I/e+D
02V/T7zXHP+iF3165DBZgMGUnNV7+sNjUuhy7AhFQmgs3dku25Z9BBI4+E94aPWA
V+xs2boxrm3jyvi0N18uy4Tn4MoUvuIrJyrWU3SjdweinoperHQYMEh3d4SFCM0B
ZJOmi3f6/TurRQoZ/PP3g9IiXtDBvPIT+1rIdRULhhDzp9Ujkfbp5EetKuBRY5vq
4YRKQyN8fcLkDUxCmPLnxMDZ7O1CYbt58INWXhK6f4HXyAWK3azeHHFjCYXqqatY
sGMgYWywQIJC0HyOA0m0UMk1mT3ALRVZyEDLjA+to+WD+rlW1hkCYKXBmdGbLGnW
VBfewr0BQt20VnNlGDZa0FLGsCcVmjReyqolYLGcMthLfTZVadhHA3JX2MM0afeq
rrU2xlI78Q5TZLS+9HU336Xe1rX8g0TSfQBlaV/2Qr/5PXucUC0/eToLmrn+jcRM
yC4IiBcizTBkiYZre8TYiydLu/BtZSvfeeofA0CtURQeA6Dd51AMsl5X00d8ONxB
A9BEw/1Uq1wEH8tjFPP64m+RhH2XRzGSQ4tdbxSpVAxlzCWibTbXmABGAIHi/Brq
JKctC6TmfyFtaXu3xQ7MLL8pM/qq0HBB6V7X+SaYb7reAARY2L4YSqwquQOR9nz+
R+Q3hgN+9K6jMx6IVupFpx+xKjsafyF93Tfu42b6ntf/drus3MSgYqUn1Gn9WoD8
QsYiPYDHAKbe/65mDb2Hhxa4Gk/Y7mGwmM6ROq7KT1puR/LevblEOHRYaYaxpf0I
zUc0Drrv2lwzamnzmjUoBd6yJwq7IAqU/+KWQqrsIbXXL8jPGSvX73MyGxNLCFqk
ep15zTN1mpQI0N0KFgBcOZ30WCz5BxgPPY4E6M1gHd7UUc+SXGN1UQ6lUWENcV/Z
cBBLW+RpYOrbz7QuM9ql/AN75pVi+wXxDPAD7sRF4olDBzKnTeOkPJs3RCoWMLeX
7THt+RxcAGT7r3uCF9hSOnXm8cP7F6e58FqyPcZAEvcG1Z3AKrvfHVBHtNYAZhg0
kO7xuwDBQuuk1yCCDpL+JLICO2iUat989vwiULNz9iwNLQ6DrliK5MU+IxE6rib/
r03lPSv+/2dFm6K9L9S7SpXmja6XNybLyPTZa4IKjaPIkKBWkVtW6Py4tp8V05jW
4vWRnSbGZzkK+cFCvyW0DLS9DnpGLNX08X43MKKE09WFzGxbbqYnoA4gMUa/4QCs
ONlXvTImAJ8lu8cXZyV6WSorwlkSo7+T51UVV7SGpBD/6r7IORCgI3A5f2LcXvFQ
y4zeCdOf5sn/XrVFy2IvyT33zg7nN/is/Si3ejQIyINX8KEfQ+XWHZ745mAb29Jg
IX6hVCbDUwVLBd1pKh0FfcuO+hceIKnAXiqgGobq24xSG27SRss6OMTL5OY46yjU
vVdHluabjOBfzLW6WhU2f0u63T7pI/BDyzeeKnIpEgB8sCtopgg93wDzNCb5TEjD
VDOKo2oXr4rR17zoLNSmCk1FeSFEGrRvKltqx70OzaW4VRU4IJJ8ZrEV52VZ385J
Sn/ByzbsgWNdVP3gcFXbQMaq1I2VaKunvhRovm9K4aI/UdvdGrTQxVAy9P4NFA/T
TH4dItrwy66eQoE9129g4ADvo3/4b5mx0/HSR8WLFWf9lGHdTIt9xgl5AJCmkniG
eQC+GRqvUsarNl0YP51FlM6fZihsv8wJspoYtWDrBi5+6Y4fteNdFpFUMikeI9Sp
7PIBO89tTgdc1UvFbRVVwivjvCBuLogZWFQB2ojP9Re6+p4dvw7L5L6QCbCqcDli
06VU66i0feV+Vv+dcv/vFT8H/iPgmpAScfDkZBv0SKQ8EE5kahIJOTMyci8Rk0nk
OoHjUaPV9cQtJ/P/1vOnRFLJtqzQjG/ABkI1LIv77Wl6+4OKTaROyxiepLxEY6RU
4jqveZLRRGu3+1C1s6c1aiDUvALJO4vw5kcMVXapc6D7LiWjwPUhaZ1QKyqoB+1T
`protect end_protected