`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
zZSxD+gXg/oJR5jdsH5AQ2RSsBVI0tb8VxmTK88TCDQ4gf+irrfgkrDBjhYsa2ft
3hfVrMETSFt4yfgxXBjj7xunt2zekqpGcisa1h0mT1IefNiSiM6aFreSL9qdnbyJ
JRLXkgV+8Q2G0T36QzGfGGvxb5IIJTsF+CjbDRhZDzeKYdZidRQwJ12nvTZ4QG91
pgtxVsAKYBVQy0tx0NITLh2H7eDby7/FToVu1ZmklGUOTBykEHTzk3473iOcBWFC
E6brFOeHJ4rs/SYbqq/qaVc/Pt+UyOXMCuKtJhPppbDCZtfpJytFlkBILgplZFoV
ts6gcrEkVC+5+L0szv5C2vOQsdntQ+akx7GYOMOlPOUxlgk7nGxdadQIvi15gb9p
nddIgOAH+0/1NnYLe3Bix7H/UFueYt5mCQoP9m6HG/QPZGpjYuZTmy4PiQ76AepY
QQmDMMAIHHCdcRXHQAMGbYVXrQgPluPgw+uuCWy6eBTqLDo6fhS/oO7HT8rxYlao
xrkoL+eeuinPyp2KNAWcaQeSjGUxWaqrUAp9RqaCeQUVexCcrIvyg8nq5xyJ+J5C
HStDfFHQH96eXTaOCMZ1KznXJciHMYtLkUZxxYdwgaFnFDKLlY2mAI6bKK+3r3cL
5wfvKoutS3ITNPoB9uCxVDbZ+ttZ/Lf8eFH1Wgrk4QFUKGQQz4aORjfyZt68sU1N
WpWtF6adRa369wLsIU5JAc/zL3vK4pjIPnkWdp9xUsbBJfh86H7Jeqk3hRyFMjqK
qc98fvPOPElL1cZMRRNSSL2wNZOm19nSe8FIy2dNHA6G6hMU2X3qn24+tt6tVE3M
Oe5xMBG64bQalH/rKleZnAH12xyLxpxtZ4Zt0XiL+/zC41BF2Sf2yK2EvfvDz+ph
MqD0yMtBAbGwEH89B+hhgeWJa8oYdDvazbHHSeXN3ZlQn0NKYpkE7/LDHCsZuXGB
XecPww0ovfEW4fQSuYHe6Xo3TwVd5QxKaHNe3e+qgVQIFlG4JUgkKTOzGRlPwV6i
qTQafGgRxYuPgVhxeJHRbBW7Iwog9Dwvmlrx+zTtE+uguQuSfVtB6jT3HRqxkO7N
iRq9812H3TI9hJyDOe878CLl7/5j6mXXb01nM1BVTXendGkUpMGRMbQdBdroiLSL
DVahwQKpNl5yzJri7s2cTAS302+rDFIOx4Q290OuzGJqGYOw4xCzBWwayhYBbE53
yxH8OSp69iV3+wj86Q6TZ+RK5Z7WrH3Ay07FXXZ1wxq7u40aOiX9pdhKspQTfDRn
0d3uyUEhgG8qPiRSHtGqzXf3jiElWTaQQ5bSNctOuwCtIm/MFfYESudvLn9f8DFP
ToRnCNGPTq47ZjuW4T8axMweaAidaRHAslogmhs//VxM/gDRJX/EscC4Mc+30Ee7
/6KENBRAcmzEKZ5s9yM30YVWCb2Bzborh2rVGtvG/jUbba1MQgD/e9wDFcuSfqD6
/Epg6OiAGG7jNVsotjsEfAdDL+0ZfWOPLmX8E56BocRl65RKDHW5HNnClSXfFhOv
4TxJiUQGXNALPPcG5L6/nDdqpzu1RgED1qW9OEIoOOQpuvcRZQ8YgOn7KoFOoB1S
dbw6drxfAx0ZZ++uvN1o6rvL/gYJ+P4wX0ruuv8GnN+9IN6+vUF+QvLL+1vO9xSk
VbpNKN9Kcmv6W4ze8CgfB0KqvUMnFAJNVz3ZEkLOGC5t1bVKhocn5uAX8FC2uEp5
lY5c+A8c56Ak4l5sfo/zmj609MfkeGlE04b/TkB3afsV5nCJXpu4hr1mxwdL4x1t
zhV6lt9sq7xdef+57XIReLGyDXtEIpko/2kNm++KQXJJGBVLzx/kwJQsNwAi96Eg
XVt7YoqOo9PUpby3+IbmkaWjNnO6NiB/3Wudv5bvxuUQo/OH5ygUxt+Es6YGajnV
6W/WMl93pJf4x/6QEqrxQUwhOuNygp4JyyDvRasfd/9GdlmnSLWdGOc3bMs2vIWd
owMDCCwt9Ub+DeM9hURkrTlT2PfwZmfDR3xxb9dII4zNmE+MIYb5xy1fMdsEOoqn
SfYbpmpeSeS/z3i0kIwfT141pyMuopsrn9yn/C9ripD8cVlL14vbUhyXBg7KcOo0
PKbppVG99hHtpZzKlfwT0fUHZ5uTdAazMUn9dfII8UP9HcbgfRPG1epmlZ63fAdr
dPifea32ENpMHzT3/pgD47NarE6WCzGdfjiQoTyVOO4yWRt61HHnOwQh9rv20uYT
ejQRXFzxwTxHQkhy/JCgBeM17A07tBUiWa6QAS50iUwn6rBXXCg+fsUlABNvYsQm
LlknoryN6fYhu+Pr516xBDgMAmrXwSCrsamiA49FHE6JvxwsYQxyhgyDiXEJtAgk
4RvErt4rfR+px9Tkg/vVQ/OFrJt/MbDI/yGl5p0msFVwqfH1VX0WSrp5Z0U0hfTm
8Lx4dHAhtY4u37ovgdnXoiAqWdHyyz5KB4Kv57C2s+s+cpZ0vPwCuIjXhVLZkJu5
FY+orp7N0DG3jBvZ+6FVhh7ThtDrmYZphkZ6t3O9NalSdtEB/TnvJ25E302dZi6Z
R/hyQ/HyCuIC7uXfTiOcJTqxQdTsNlXtO+KXELsggjjoYrlVyJwhhbM3dyTxXxR7
4riA7OPK5dsISa5oWWtNWB4WgngzEPppKsCDs+dWJDx2qBcgICaQisUnELTaMMF4
qc5hVg9mdo1viZRpazJAjEbO7hT9pMUcAGzzx+rr14Qc/olEHjHzdhXBOFocflDq
M4D7/1S+QWwShtKYby7j/XSDX874Nu3NAjn87kG9LzN0mKDWu5W2HYEnJsApdGSv
kGMJpFP69o8pYYDbmAMzihsiijG6QRR48YtQFaV8Ctc9dYLayiN2oms15WuEEc9G
aqSus/RslsBpXgiH5sDWkV9VH4aSPKN8T7Gwf8KE3WQna57YYLVEsvnzqNgH7XD9
oNDWYp3Pi9N/AoytAhoMwF3tqdIssC2pyAxNHn1zBTkrLbdSqYs4xsrpwK1Lio3p
OgpzoDz1NicIIGiM9Mfn4acq3H8W+zIBgwOtkGG2qnAX/iZx/7Yk/LXadraxJe1S
JwfROctfNojtKR9CjYHtB3k/Sjim/OzDs5Xqo6/C6tB7LQqj9onW4pguyqIr0PYE
hJA8da2BZPZbmWa1KsCyEiCFGBHOzEqvMo5pKKq+F25ZU7Dc8J8KA+L/0jVJz5D7
RfhhY+hnSm9WYkvXUP1pfNbVMtF/AJF4Gd1fArSuuTbk0DaUO9dRxKQRJ957y065
pnyonxERfoqPBWE8YLPdZK4SNErFkNwoo2G5Y/aCucQfHB8dJ3zaZ2Y0eJ2SJd7Z
RejxO9RdBCNpJBVbcx17UMHSTes3BEyT0Mt1oAuHB1AT0yemmJPD/5/QkGPfM6WV
oDakF5JtUDS+B6X3uPG2Hrl+iQkz26+QmbVVLz/zWhJFi3WKiIvTrb080/PZimmq
/vUX0BcQq4RJIJsmbD2fyFLQybV2xdZeE+P/YOSUF0NNvajH8bZPI/cWyYrHwwyn
NVavrC7Wcnh8iFDwdRqZf1CwtFsjMTU/AQBnjaKq3+/OydS2tDYT0Y/tJux1mnKa
85DS52lg9gLSnYQwv9roN9qhf/gX1wYisot7kEwJtBMp8BxQZ7riCrkU4L7QfC0b
LhBzWz59y7H+jz+d6H6OcY894JHtFEQEQIL/1TYvTiatExTBWYqpXLo6bkQU7Uu4
bmox85UdFcmlj3MsvoqeBE34gwT25qX4tPY54jfW6VmjGJFh7ROn1E2NcfVZk3w1
puIqM5NzuuXL6fKiAPnKl5NbSZDa69FgLZmldaBL+t8jBt6OiEaq1WdM3n7ESYmE
mEaQ8r4YFUYLcLpUdXQvFFTqUeKR0uZzUeY5SPMDrhwnhNWjTeaoePgsWW6H80sw
GPtFDrErwdKNJlDR5i2bRyqvXaDuF3OFoFH23niNjjpkk2sOAmlbr/+pg0XEXQDa
wDBQ5UBtErOvJrs5IDEmL3uFKMQaN2s7VIIDBlO7HQcvomJFXE4UuHv2yVuYGCoW
MKh+GiYl+ibFEv72juZqAomAIomQsr4UocisQ9pZT/hlIDV2syqYKSjLYuQZ88eC
NkiSkhtUEF+CKfqn/hGcqxq+73hGuEFowSdfrll8X2fVyDuiTYwdgQeLJw3asmt9
eizei2g5y2J7lp2bkCsuYgEEkPM8BY6oma00Gio5/S3kBWF0b8ZPC6WnXOh/AEsz
gxgfjBOhgNzb+bXesfVuUE002Yf/Us5yo2Q8KHibLrZRuCaQVCIm6sWwMm8+2IoA
G0B9+RFJ7fI2XQk5xIBjFfLBjUkQtPnRkiU7MS5LKcNTTxEhDZC/ICSHdeEvMWoF
jA8O3KLmhO0+yml7TWmhfQZdae+aDuor+vlD1jG8/OfLrMnw1gOQIH86br3xI34V
cVaqK49zhZvpgmUJvdFRrcUawUI5CFb1j/mQdnYxOW3IWD8lMfbq1hs970KINjVr
bMIIwHgQpPx3QOd2w3x2ehiTb1mlQIySqOmVAZUJeC+s3aiXGl1Zff5DMnTtRbaU
VyN1CyrFTFiIsDt2yrJTGnRUYQ6e6QXh2AjYo+QvGkl2f7IPPxL7/fFlGbWzcprg
lLcTjGcOvWmbzc292NIyhnvIh0yMtw/6X3kWEGLbOCAnClTqk+mpoa1MGFxR+DTv
cBCvTO5YQOSgePNlZzx7xuMRSWJ03hV8N3j0GwBS+3V2aVdrChGv1E5PzmKAqUpk
kBtYBGH0b6+NkGSEZ+IHABUw69GnG7qPOKKR7HbYMgxU5Dw0Y+BEfw0LOFJqx0V7
CteZoJueYAKc6wQ/ml9GFpF6lI4fv/frFN15ZAazOw09m3PwbUIguZlwK57H6Kj7
3P8VGSlhfcmNt5S4UP/6/WF+TSH+OSYm5QmimhrbD72/CbblDgVJiFdxe+ajmmxf
S6dmT4iSu50tW1fcJ3bFXheZPzahPR+755/CRHQV6lNMbTGTO2/KHl+e/XAnIjJp
US6d+Q4VrkaWqB0XEzPHCDhilCjaxh7DKh7Qiw18m4VuzavsGZwVThzEAmyldcBp
UMZt1+smFe8SDi3UfAZ/iW4YXTBz8lc6VN+08WP+ikzKIXutIdp9VnKI4YtMF812
ee3VyfBpTR/pb+Kdb8OCrC56kF5O5g+xXUlGHaoPdVd6YYXGklWLbK7TtxH02SBE
JF1+jBj3LSSz6fUgsIjq81qBkcCo6iXEP3TR/wvkQIarrHh0r01J+vafnsDON8H1
0LT8CjBmSP3qTPf6T5vqqUeJzZ3CjHvber3AMtjYxVx0aJNWQ67le68YhwQc9ye2
9mKsf36OkNvfRNbBDl1BAlj5cKzLcfrsMhuan3hQonPjX4XkhZ+9+WyRLpLFNFwd
MhKv1e04TQmlGeivVb61cLXujHH2LUF27F07ORKhGXnmi+TJKLn8A6RFKif5u7Df
Im0ycnX9SVK+b0bL+XDUfhlnGZMouJoeP1SOr8EswvrI+cV4K3KU3DJO6gNABJ51
A1slk+/VOdeBxfmh45/PMVflB2Z7EEBZtt8qa+YRuwp2Q/He6qVFjsiDcNDrbIxS
GtDMXkRGtAx8psv9iHnKCz4BtkrqAIZe70tukcUYglD0dxTAnFByYIIOCP+Jv2ns
G3JJTFSGgx0SfLhw097DY3Jjs9ZoAOAWUr4FEaUx9U2Zw9d95D6dl+VLxcGDiDxZ
bn1EEUREYzG7jFGrT7GRn2vWV6EvEmgq+9ITPNm301vgdVAFQul95IaqsVDpfd7C
QmL8cnKj06fnQOpm4hcnD8+zexwCqzx644WONkMT9YKO6LrWtr28R8xdLit6QXLW
b0wA4kp/NTIegy+Tf6xBP+MUbaAQrNwAurRiumLa2WiTxu8rhkmtgi8voGLawVit
cQI8O0bP2Q2PXHayOvMvb8QGDTthDwS/xUUvy7CU2wNlPDtSBXI+PkOmkVPvI3Ug
F/QtC72OmY4OU1u9YdNhDqLx/BDfITuHC4RCh0mszYZasgIWiX5Cfw7QvPJDTYJu
JZjn6rVTr5PCFENXaquuoksVeeFr0lzHsJ+bcsFeF/lCUStHG7ZTV0HFGx+NtFff
Sq9X0BnDc6ZNCA7rZQ+sz1AXx+oZT7AHQSuxNIlO2mWO46fzk92Jq838DKMey+Ny
5sCYYu/1RKloJT6a8F9Z+CEXyUNa7/8nhQLsTwM2GbbK2L/0MqhbijSOe9SjgKNX
CeXfKHztHcoEpxFeIiUSYVbivWjAkyakNbfnGcN0LKdZPr+CT/y1jEOsSzRx+9vc
fI+yhNfxjTe8vYSZmXAKQYkVsO1XTZwbF4MznEmNiEByV7+npw9ElF2HwV+EQmxq
be+WgbatF2BlWjST8kn4ToHtcp9rV15HangampnAPzFUv34ohvFVkoIS90G79s9H
PTBjeOdSOShrHx5kUAPpnCJMQPmyc0Ct3Eh5Q1hCPQbvkQvRKbyujyHF5Ziym3/I
Hbob2Zq5gRmqkUnylZZgWVk9J8QMS88OrYzr8MDGlxNoji+0Lm4lBPghVEFixgaR
BYzzqQRjp0FsOqHhpacjky/Y/qGqmGIwKbc7n2nywvIJrFordltkcRM3sICZ7iZ1
9X7sjMHtwUxsPG2PoyetJPXcbush59SdXJTlGLjFffecZ4DWWsDHls1FUMPUmDUm
2p4ScEoof7PGnc5GBR26oLRHXhzVdlo7vaHLN9SYx7UwPJS+7qD/nnxArZAYPIF8
jAr22LOMCn1zx6b//dB8XS2vDygi0uHGxGvHUyQl17Ey6hkKc7iktmM0ZUIe4JeY
5B0NhRRGqpY0xlgzfoMqfTRjWeGkliCiGYZundKtFxrAvkMGbbtuIY9TEbrn1QFZ
q3R9rDv1epyU06lWJ4mYmhAg/TTOENythYonPKqw8YtW7WLD1pkqWVatijXfZ9Bf
vMOib32UyDNG1pQS3VbthKWd36aDWI85DMOUs96ojypx6c01EriDNczdV2yjuuXL
SGLVINB2iGGuWC1BhD/2LIjQ3jZvNZy7AlVYrbYvX88VLKYzKhRleq8SUlS7ThDN
UBTEll8r9zPt3Kr5ENvFtGeQJYZv2FEh4tLlP/r66SOtHmnBqaw3PAYUxhg2iPPb
MNiBt3ME13ZU9GeTibVBUNGu6UMPiit2eqWoS0klKCr0YdgjeVwBTjhz4wfwOE66
iFXTSgP0khiQZCoM7A5dHx09ju+RJy56oNG26r8t1pdCl/uvl5muJFO0Ans7KPzz
o0HNBVVTElmdCTBX/9VXY1i9BERcsjmN9Sqw2Us3U3zhIWWkJcvRrs/ZdOtLhwkZ
TMXJg0nP+XlQu9sOjtcKVF/edbgVhccxf4DqA2sRPTnMFqtBHE3/x/arU/TSBgUx
ISsGSLULC6dQvb5W4thq1TYW9/oH2OjmGpcUpxkX1aFl0yHtMus9vXVon1MEHl1n
EzNMq2/isKkUaEGZ/KDa+GxUp2hu0kH1Yn0INAwVdsVFUhX0fcapgpAV7SbR5+RL
O72GT+nvNnmUt0PuU0DxMslUDfYqzcOwhPYv8c1ZbWMKedVbMmPxJapmm5NReo9v
YJV/L9LkTiaw5Kp27H9ZHMtWHVkmwzK0vwswnjrdow7V6AtUJtMGPwQvAH/Q2coh
RM8VGARnkl3ew2IVY/igBsB0Iksqfd1RfxwKDfAzdxcKq3TfAyj83LZYKRF/1X9n
ZQ+jUnZZaEQdEuy+Jq+YU+zGDF/khhIdBV78Fk3hSp07Ut52vjy051HMcDUNL1x/
9nTypqZW6MEsCCH0LWgDrC/nRdRXickLOByv03N/q0ghfYUVXEAZCuE0hh1+K6SU
aYZdD54O88osVtnB9Fj8GrbEjV4Sqr9fr3lws5DnH94h7qKGSnkg58h4gvVK+rUk
8x5EomWL82hj6Yi3EdQzaBHOGOXm8//G+4hh2VVAz0sLwiJuvFnsqwvmLlZa7vzF
CMcJ/DysrKCdZXKwqdiFfuqvYYFodioXX4/xBIuz81YM+3ZcXJy8cs/psPwfF6H2
dOqpIoLPrgSh7tKNmB5LOw3c3rqaFJJkDUeHPpu+038S0DwrsO5nAp+CSlu8FyoN
Y5JPxjlPYUzOlBrZ2vOH2oa9SAB4IR8jr72h4AFZQq/n+cdwIM0p00+4RUnlVF7v
eeb2BfAac9U1fKCHGjUm2o29lhScl0f6YuwP41eVQFPNyoO8eu+NQOmc6cBcwEno
bBhgsz161YzzVefwjg4Pj3+RGuvihEjNiTP92RKfFdNnmh82UzkGrWl5uyxj0i9l
XwZhPCKhe5NHj4SgQQhcerX15rp3ty6sGp1xOvU8xZ/gkV/UWiRiKDLQDYEn+2gl
PejXcHIpiMqsm/qPgIdriYObvP+Ns/s0GW/GPlZZK2ewdSfojJE2L3fdI7QGaAcD
EdbCSI5cuFxrQraris93f4NeFJZr54jyPN9SvzzqTVRE9u9KAee+p55gtQxEX47/
2tjW1zxUX6/WrWBDoni3yBk/Oul2+u2rm2WBtFk5tq9VqEkVAGqUhQBVKWXUuPJU
N74NolvEnN7k4hMcYiIs68zcDrGiSyL3C1i8wWfx2S/KO7R9dEXRLp2yBHpx5Cvc
3wMimvGb9SPavKu0ezew4h9RFfEmKf7XrPvTPwGYyjLR4M/Qg/Xx5yHHmumreLBP
VT1h6fl42xRLzZbl+nCAEUftbDA7oS8BeIHqMdakUVt9fMtCGOzQed16iEac9rg9
PvecU9I6cj/HiWHNKar/tB9aM3K+gD/XKxqxXyuvfhivojjbL9HmcU8WG/ZFHZV1
Z92eDzESESHSFdrnc1TqQ2Iyc64vdFoVnqEFEik7cAccM1bOBii7pKaf7PbH1h04
A5Hs8R65QpY/qVLzgkdyhKJOTbtBqWQXxZ9RshwZO3+7MN2LiNMtrFjMVyy9dU0o
cwnVpv/qC03FBDp/u/dA5BPTlrpc8eSPYcSDyiSZ0//u1DaV03rchNLGRLNEwITB
874DHLjRMkHLm6Q9PlIh4hsGjel7GqKja2EvfgUL8A7zV0ndGK/yUnjRN7Yuouwu
OuiDeVJsAaWm8W5Ft459/ZJLTOFQwsiLNOThjmKN3M7QmXnBQbBFUlk8S6aac6DQ
c1HYDMyzz9GCe2tdMiLt4nguY/1MNaD10h4kh7M2iR6aAqWpakK8B6b7jfxRCN1T
1zpTY0zJkG2tKD//ohEAzDC0nEZBV3r/E33dwNoYmsPMewCm4ADNXRxA/F0BS2Xo
Jn4Pcc5WKyHyrNqYEvzadnfH+kDmPeJIaIoyVjJ6EVKLGeqt4R9JzsAtF2kuJJ2y
Men+9E/C08i0k7i3g+9iYih0zO5mMGFC0GjUKeCqu2Pt8jyn8WavrtilgQHSA3xo
+bonKEW0zhyGhuJKiT7Nmrk+RzpwEqvVmdd71pSeYd13iLoxCMJjzXG3Ot9ByuYr
+oVoErVjqI71XVahzlpVn8aTRX1Ncz4X07/qVVT9LOeSMIQvfA9wqGTmzwEI2+cE
gltm9ipPuVpZYZDEh9mZPEr7f08BBtWg70SK/wr4149a7Pz/7/xyVDQkZv47rmBB
la4+jY9bTec1vzBG/za5z+VcPm64LM+5ekKc3R07ZYJneor1OU5BoPJ9wvI9XsMz
tY2aBZe5PqxXSpfo5LO4G9EVFPc/G0BN1XNrqxn1fFBku/ofT1nSx1W8QuTq3/c+
XGUx1EM2HOHg7CGCuNozg5IeK2kbGOClpS9nDCku5BbiVsMVZtpko8ij/Ejt+hi5
SQiRJ0e33/P9kXfyj1XTYZCrBAHjDpptm/GuyzMz8Wi3/5YR2JTrTdVXtl4aujhd
yywDo0M8LzJ2j3Hz7Iik9ZfKQsHmWh9j6SGJb9F5wqSQFryI2kVM/7S2fAVA3vok
GAE43BKtKIT+FzxN42ECF3PYJD0GoIC7MM2mFHkpkEN/Kz/systSLifRNTDgdZvb
yYBne5r0fpVP1Pib3H/JUu/v0Fm3+RkLfgMzMnD6Wd49a541Y6WHen/ANVeUgAxB
gHSbnn9pRxAuxp4RoYBAlVbkwDpp6opJ1RQCr3BhU35ztVQVB+dkq0LfhL9B76Q+
DCeKnqG1gqbY5zpKGC/L6F5Af6ENYPdJ25sfYiFya+AaJLXaNBQ+yEQeFg7c4W+b
uqM5rRotgoPEckhfLtpPquiLQEdw95yhHfEfh56wS+KvOxVNIdV1NRH+a+ANJKxE
FyZTPcNCAse9ojE1QDslYdyEeUn3H6WfAN75xCt6IeZQOnki1mh7aEsvCXTBI4oD
NdnSbvqLlaaguYOqqBzFenVDzqawGoYHkSqFd4SXIfsQU56GJOfu2ko7EIgjkNL7
gWLVHXIN0w/Mvm+5Q5xGBD11DY51e13eXvchKF0WDzaHaGsR8TeNClQGgPWSOd+T
y2MbhzykMUFzXk4cIpNVfUEKX1JuGASY5WX2mWrsDrUHrWjspY+bV9SbpZ0NEDHO
s2AGJxRSYSvcP7YzUnGKSfsFLX4apIaPobLSpEsAnuwwfXrz5jePu+KPsYbwqtnk
QUWUi0+BqbWaElOPA3epS8h5HqkcHAUevZLzRV0C2lhaUOLcwgM8oe0drvJ9/AvA
6zEqcuHdbp482gkUbWI0pKD/9h1KbAh3gzoxu6JSmei1VlEJtZQyl/6+tfqPh9eX
lb/rZO51+IAtkC4q4ioSY0VMAOxXb1KmkU8gIyeExV6RPlU74DR3x+7D9CHyIOPY
nyfxRVrBnVJBjkvTHXYblfMLGuS+yKO71FsNAMcbQaR1gDnHFxQT/oClXDvWQac5
/OVF5zXZIAnZaNlWA3HDw+q2nC7bqSsv1wQ8Bxn0L5o8oWGPG2afiUg4ZAJqQsQ7
/rwIyQEPHUhS+y+oGMSgY2spEX+imvdT5Yf6TD+9pLV2WkPF7Hr4ESp1L9qOQtcz
MIntgQGQPB+0CwRHF0kQqwZCEgtazecfA/p5yTMDBmE6JWzxfHLauW65RvlNfp4o
XnumfB71ZuHN35bnzjehxtvPwuc4lYQuwg5GgHTnjxB7jcJkGYfCcpiq64yw1pM5
fNp3zZiA9lRHGyWtqLZmJFH+WQOlKCmL+On5CCjXauvaTdu27GYIXbu+HB6ZPu0G
bzJeTOMmKaQRmqdrocYWPVw3dip663AeTouYWAUf4Wg2knDZm1ScBPvgbW/yxkD1
HGUxP2ncAho51OR+iNE/oH+ixuDEoSqrLWNO2jJqGByVACSHkHb6gch+n9YJbbq2
0qlUTbWuRAR+z9SbB8utSiOUkCY4v7UbKu0oehY74mBZfQbQ8gTI45zNuZKztObh
kmXcypyATgrrJWBrwzemYVBCmGgqTHWb0XhWwbZeMLjol3VnAkdA3fMJU+DJyelQ
XXcKqgGEqlKP8CxC7G738yagaccedE6fWQqdbTQHbC+DIHSDQdcBPjwi7fmXfut8
Vp1Hwa0osG+3PBBRg66DoStoS9rvULFGPLK0NxlMRjPIoW/QYw8S/lAWqK5PNbex
0aBX7SCUA8Eorhir4yU9KzOPUNKz1EZKHjFimz7xKcsLyZC7UnqPcVnbeYTu2v7D
z7sFhI0Z0RAXUbOdbf0/Ez/JNqb5VszBgTy8fkDZhB8+QvFtua6j7VGISjasMU0K
MrI4LojRyK4haCb5ih0GBtEYI0z43IVxEVCiA/1Kl31GOZcw4p2VPlWhKHlfkBLo
gN8+rMKtDAJPH2qCpdMhF5K+JyjwJmSEaXvvln7i9w6i1cHhyhVRywezMegiyfos
zWSW5LS96zACdzSkqSmza2gyPKeydujW3qymYY86fvdMKYyf7SwJXBWZuD7n9p0m
bvb1rHItDJD2kNCzl3tJqmVr931R3RvFEsAdwiImafXKHS1lvksvvmlf2oqmu4iu
UAoCnbHxMkOJKKS2i0VlFUbp3O6b35uafF9WStpHScSBmk5PUj8sg5yS27mHzcTa
S0Y4CM/wFj+4Wuwqs5GxkShWOj8YgI3OdPa6oTxodxHx06NSHN9BcPKNb35Raeli
SPBIaLYb9QsRjA9uEYSeqJkj/6UDMLeZwoIS8fgxvF2UbaPx5Jz3U4xBsg7nQAhB
vf0BdmEAD9JtLoBSu1V1ym9YDsBmCYXmBr8cug0gvmICh3SW/bo6DAQP0PPv/+gK
h6bz3gZhIJngnYJzZakPST7nihHYYZRE8M/zil1wSihYlmSjTxpSFicpHrxFd7oc
D1ySSz6hz63W+xGbbnhiG5HiTr2g2X0mAlPE0gRdamGp8o+Eq1oSGK2wPXgCcjHM
tEH8/KGOy2tfEMx3IHgn83N0Pntzqn7EKoUmRWqCzlo7fIUkGSLwMAxVRUbifKUR
SbF95ryOnmkYfmzFGk971bi7m4Ue080Y5AUEaZipArtawDDsq7H5lYcAI2NB9Mck
sgHLSNedNC0MhgsW4WTxKs+XbZCg6DR2jZCA988KBEVbXE/adJJ11sIYkv55vAcM
wXR3CaHS+UkJGVUbtHEKf6knIuJBON9l4eyoukC8/XkKVeaeB4eL7mXsVG2XFYDL
WhTHCYyhu4DoPs9x8rWdAkU+5PGjIyOBYRVI2ULBJPnku0cM5QM6td459y9WVbZA
zq/VnLAgrkqI+mU7yEkAYAGYJfQ7/3yJGQyAiCAmS/k+HHOIOa5KzUw+oTux661s
fbT91tlqDPhhrPIeHBH0phn9pz7IFCPzlUsvSCT03mkyK9X/1I9AoJ9tB/Zwi2S0
PNShsPPahS5eAaPsF6K5TeQcL88PcaOTvzA+YR1yVhWZCkJdWvnrqmhXUG/OVTKR
OrjdRIvaqihl7376EqDpTsQSS5ABl8CiyD0uDeb/OwO14uiWe+bw9LK8nVS4ABiT
9teId6O01mF3xJdXVYeh4y1JWVXYmBCBT0qE3VsL7VwLSDUkVO3mJlu/tN9OikEO
Z0CD9IoITKHVkUyn/dwJkv2Awid+HroKzMvC/S9K2uwL0RDL7CTo7kbY16o4A+fm
3keOPyWZIXA5fn8CbdxGxeXTuSUMTK5duV/vYiavNz9+n/92QEZbw2slyHH9Ys4i
COY1sLZGeqNWTbbW1YgLpDJ2TJ2b6lJikDcLJpT/+50qx6mSEPqhpUMyfviebiKP
eH5/tDTJTTwUQFhI2fONz23gB7/pXV9WlTNW0lgKeljw4sRG+ZBDc8x4xb3mmeOq
1/u+rU+vu3UJVSJOEv40VFwxQPHNNI1ypVJ/Xm/hMVpL2cBjD4f5fBlEH0vIuHpp
Jn0X0BS6+RwTMcUaj6klKjP/9hOiGJyl+EgqmN9sn5Ak3cW6Ig3aYe0BuZfJqdBF
rrxUmB8Zh0KMZ/DNjI5wMM6eu3az/rL/5JpPblImnS6TYe+ZMMeJjGF+EiKfGs0Y
GP07HHz32gEPpnuQrYQlzxUwykVXFKBhQISxbmxcIcsWbrMLT8+86JVzN1Db2wbi
tgnLrqOJvE1lOjwNkwe36lbJlN+FNfd7LS84Hqf9EHEFMW8dcjoMnYJgxlOJFDXC
/SS51oejEf2MyJV7WYQXM7rKleEpxMZzE2lMXVvGw98MQ8MoWwHS1nY2Cjsr4RvN
yVwgdHgMW73ZFZF9hsrRKONDaa4ynhg/IEtuAOfgN2AP5cI9/tUceSk9XLLOntF9
+zkVvhcnWcpsZQw+WkWu9Aj7EfRprlDHHlUn3xxf1/7+1n2xpNKLgfvFRhc3NUCc
V217P6wlSxtRChaLJV4SI0L/PTBMrENMVieunlxR/XC4pqCXD3BbcqtzMhKsBXTH
l5kyQNB6QMDel2Q2h93MX45EYRcPirh131saERjquA/BN9ABq0gBAOq15PmjrP6H
Go1YO1hSnHHE3mRwcn55bGB6U2cmz69ohs47Wku2IhGzjTxefdLjUmXjWn43SbOM
5Bg9tkkMiGhGaskYYQC2e18WAnHdxQTocNJPegTFH83d/SZhdxRgnn1icF5zVsLI
UFWxFAoddBuf6AyHE3k0P3XwJWgtLjENQfNGQDSGDs16uINyb38umiaBWszpySJC
RThw8lqknMUT2fBm1HJCOHqjL8TkjPCYrSC4OR4uUeBXotiAnsxMXSGej0iw2tTQ
Lp1W9YlhcvexAYfdZIekm2RhGiMh79Er6TXOE6kLkBPyZKI48A9tvHJGb+ZkGEUZ
8Fn/tOL64g8+7fRoOvCb2yjPMiouh6ktGBPqzc8wYBLJ3o0Xn1bgD6PoAHgRXFzI
tVOq5DMMPrmqGZEca6ASqjGe/PqZ3khTeZAtVr0qfklPe4WS91Py5WjO6iy7WgWD
Hu/3bJMYM18ERGAJ/hFP4QmW07017wq8cqOjSlrDAIjDLEL8OOZW5QXCrwcm5wwP
HRplJXl6OC7bWBDvkO26P4LzlFgAcQSTNkj1x8hKAdOQf/d1AA3y2MG6svoHvffo
vGidpavhsJGPNjPTA4gkWkIkO1p8Atc3QXjeKYBD8LFnwqjO96q+2Cdqsy2Cl62v
QrElkzqTeaa/25duPy/mH6i6cHXQD6niyWVKuitbuIMNolx5YzZgmch7EP995bmk
zfEqWAqPPsJyI92bq6RuD82/HQWbVdHdKCvlZdvxzcj8IIv+aJbWc12IBEyf2Yjd
v3T+KhuD1x8N1qeb5DwrbEcfLHg46wEOHVxmIfdP4NeVpPtHg/MUfLMXEtWVEgDf
Gm7dlvkFWnDa0n7qEE87pQZXBg8GHdWUb5/r4pFkWE9h+dI+TxsjStcdPwk3k6lw
pYgNAuZNcoic6mmmMISUkiTyNo66WncJLLBzidsx/mUHgLZYq0R/aB0BWWMOTtQx
3nrF+u1Hj/Eki4diNBgQa7xDDTJjL75T81K1a3S5NIxkXcEZFHUXCekgSeH3t9nq
17GPn9SU1vIZv8uruxrAzfxXCCbzb1X8DPyjJM78SKAM4lEPSdbtzrhlhjNCJ/pZ
iMBnGfxGunY1EhXSSGfNmFzTMUG6QaWSWN7Ewhx7xPezkWFQH+VjZ5zdp3WyjGaE
F5IeiFrqZ1RUowReFY6olrFutq3mQJgyicD7A1FpJEuWOSMGIkR1iFQLfTXT0EXO
l5wRd84RzVoj9PiBSs8wTYzwxtAQ0Ix++Mo+ll5RULJpCvSIzAXgc2BSodf2xgNO
TjeqM85hEX36QQgZMieTFyc5fY/w4jWaavYFJvI+2NDmyo+OUEYVdxamORPr1neC
Kd/rh8tKAsMvILcoSrOoX186/YHw4Y1nKyyludXRorO5XMqmJyc2cigmTBk2sGZg
/ZMG2ZWaEtAOTvTsZf9t2W4n9p6DzajOEpTlMuSfpO+KgWjNyRkhLVCmmqjCmXL5
HM+X1rEXiknDQjW0ytt0OQrK7BsOfZtSbpnqSsIxmkwsGV6jCv3remKyFMxQK2mM
m2oQ0v632DTlQbzA0u8VyWKvtl9TOu0Mo0FHXq2Pm74TTlwcitkNe1q3iWui4cC/
Ry+4aU3kcRGnaRXtC49LblW3TVCnU8j2ODgrFCkIv9yqUJGCavFCyj8dh0ect00n
O/AZF7L+SnySeti9zZ6by8oxlRKsU0RIVF3hvqK8kTMq1UK3NwTyq0pihuz7VeSb
vTu8bwvrQx0MDCd/MVPxi91FlJt+qAoQd81kw+hvj2wcb6VcsqqW454aBEsNu5ai
PtzCzeHc8jjBK+ihS9ge57Pid97ax9JORhQwgRnzZS4BXYnsn8olIhWDJrVFQBSo
u1OVEPosDNJTlL/0OsL6kG1gBSFgta+I3tT5Mr/S6K3L2ZliDstI2ovCMwoJ00dS
M03xTQV/Px6A6WWARZz4affs0EOgtddXsdfTcA/y77lydL2SGbMDQtWFytPJ5weN
0ffl2FUlx0HIZpqkJziB4b9JYuVVLTz1/RV9bOKZax3WvJWItk3R/MtrNqBXLuhK
T7qpmXWk+rr0Fk3vpPrDdVvX1A5hayR+pjXFtw0PYkcBhYDHKqb9nvRTZnZMU5yO
vwAK1l5rexwWlY5AHpAXXF4vSDmguPVwJGcrpbXw+3bnZGV7Wy/mvuF12J+/IiRC
5RDIpWMuc3Zk2pZnbvyyKvSZ4eyTMOAENzya514cSITlEIRP5hQjvRA3GVD+VxPT
JhQ0jw0hZUTDRCJgr6fdZ00ZwkGZJsPVX4YKiY4y5uCITaoGv+blPXqtgoegvo4B
y9u8xpaeglaXHdHJp71qmec/ZIz7US6wriAWdVQG3dBps/FWHb2yJEDR0RB0dJMG
hqkhBlBTcpCqD5kIJYzDq3h9R0K7ig69/fsVe4umC7m7785MgfLlpIv/pbtg1WBl
aZn6Zr91tyeLiHpLqFsn4DEgyblOf0vJY4jEpmY5foDK2R4zowAbZWLaifjg/tPU
YY+I82/RJZ/EE636eFUtuWQ+uFue3PmE/kcESszAGnGNiFBQLYrOln/AKnb9MvwQ
BVVzIHyLY8AFWRz9BwHEpImJ70wUcUIX6PXLfpss+KsTW6pQVoXt6oJ6uOVuQvoT
zuTWx4tTQVsbCtesO581NT0qcGxwoiQDj//rW8fVClt0lYlDPh0mc6Z27V66VFkP
DdJ+i5XZvW6yWalCfWrFLIVAscBvkOr2T+lqvsAiwq6cgMW/fPiHxP6Ec/o8aMWa
Zob1B1glL8MrgodUgM2uSQLBudKac8VBEjZy5G9wVqdfz6BgpIqWyzuCWv+D1tlc
Cev9wNzpQJIzGrP9vXPi9E6TR2zj/zK8az1ZgwXjC7ftSNQmqTZgaWH67n1Lgf8G
UmL7nx4rNXCAkP+akmaKChbNmawIhVjDwWokMtaCMCO6slqYxIIGlqQqVkeb/MwZ
lgKFY9z+hRn83HgRjhDyPO0Bkr4pE1NHzutjctTVFzwHgcBFlErGbM8CXKXlPr1m
NlY5Egi0hLiPGRTBEm7XrbpZ6AbMMCknvdIaa0zCP1JWtHgCJx45j62L9uE6BWPv
yE5sMu9hflwyjQ1A6O5THyhZG7Vw64lLVCZXT+X96T8SXxm0F3pcA+zzSOPlNjOm
1j1dfwlWdz9fBT+y888iyA5v+HFlxjreGu+ssFJdrnggxW3xd6fqMEM7zQG9FqJt
RA0cNzjPRG4FViguQw2zhCFcYAsQARMQlc8fiiGxa6xBLQfW81GFBtirDqxid0G6
S/Svoqxic4K9Lb43OSYsDa90xNY0teVu3E3VkJQ3xzMrrT8oCIvghZr4aBX40Y+Y
om/YK9Pmz3TfUrEF1niA8TZ7BhAzianiiCFTkToJL4MKzYn6Qlo1/FXRKDpjOdbK
J0H0cPeDew1ZbSuWvSCfPgUBc+hGP7kAnx0XCUjW3RQY3y+/98ae5f4T1PMGKULd
xsk8JnAK9jvMGtCg1pCXYDRZ020maf3RXLIjpRzkO63T1887kohJ7WQ8wxALIevr
XmUc0QIabVhywWe/CrZWDJQnsVMkjL7kiRV3X49GAtrwlIvbnuNLShQI7Zr1tlrD
k77+agq1C0faQ4ThXt4aoMhB0OhSrDcE4lFBR6jq8TtB+yg1WQGn4k83fGdu81KW
mN6TJf9cYnr/PXQKrOo0fnMyG+m2yeuRtDvuACDiFwfFrT/C8iL+VRz45lMjOCQs
g1nunE2hBYrcB4aTrSd44JJsTugmCubQIlkY+WzEZhkOxWNMOa9vc5ipyWMm5+jM
5lvZomFT/l+3lTTTBaXMFE3mW7+5KKsNxBsHT51lng+ezpLIhtPPVUmwO2FblQY/
7S5TCsezpfKHMbAM9DqQK5yWPUwKjWDY2JqcD/BikoDyrjaFRQEVMgMmsbmCwnkk
qsIsBn/EF3QwbbZjlmW/JT+0GPkro0F9yd3n8sycCtEyS4SmqpFo5Ku4qifxK4jG
0RAmL2E4Ec/SGKDiHXEv1m3rQUuXC6ylTod4lHXbPbLdNd8fWU1/dNKLCaVo9ybq
bTlJKwTixN8eQDJzNA+La4cTV8nQjefAXUIsQFzkgLVAE3vToB98DIBCAwHl47ZV
1fA1HuPqZBhfFKIZjlAu8rEylQS6WMC+Rbj+T1zjHATJs70Oy2/Vap77qNytWhib
iUjU6SSTdAIRGEpjBdoRRQ1QpNOHE6/5T6+LsCKh5cJeqMw5LXdrUabic6p9mwWb
nhy3hi+ugo7AYZWIezUtm3sArltKv17wa6g6IWzdW5i23/orT2nCZ7usHW9sELYa
h4f6RNjou6XwjD6hDo684zvgKCwlyvkli2d0fLdOy7zuqbLSILGyQizdFWxc/QEu
M+Wo5ajATGVJ+TU7boTO/CZEq/wLMwX6oRzHruTceMcJ/cnYuYfma8ZJo3m4ZFTi
tHhKIaOVrsjffXu2o29wOQjTWAcXF+2cjzujhWKUVI/V9i6fEQiZDqBicRg8eHT7
otFngg2ICQoV8MtoaRRB+E8I12PnRtheBw/v2cefC9OrLDXaJHvHy7N7CEF2klfv
SvtDeyyl6i6zuRBdSNmYagrlVWW4GXjU7dXo6NbqjfvMG2TeyCkMoaKY5h2wtsje
cCamMzBClMp71GC6+jruCmOzo4Z/TK/iVz07c2h0aljYM2mn/OF+Eem7l0d5COwc
S2iqIoZG6rl1WmQJeCdeWkQ0TmWfgMVywtoGeWR++4SuqnKq7Lu0IH9bx+taX98y
N+ElFQudWzQ5aLcR7uiPYuH90rTZRi7iR3fJl6aS5K8QS5dCmMF9KZOS3HBSnjJW
drVXbKq9UlYsoJ0+7bB1jeavIh5dKH14ZNa2j95/Juf43mEZgtQF4rmMkXoZsCDf
bbMIlyt99qrPCBu/BMmpsjk7svJsgClKQQx5bNl8/eBlyaZIZFEc0Uw9oWvfggXB
wwopYpFkCtNaFJ/vmX64nBAEr1MYdo4xjd90pMRHmCKG2zJRKLj/Sqy+6H2vE+MA
kEJ8KXhBm3EltvXVtLKQ9K3j6fiMfeG2qR/HWDnMnqqF4MW7nZr+/rwZa0oATpsD
Ng53zt1ElJ219lFcRAHkmdqkaeQw/GT8FbkBRNRuiruAMsjBfq9ejON3WljxNi7W
kFXokPjuMkppUxoZFPoLaNksSXoKtWxC2cGf2v85eYIj+jEm0uZORx7ZnRtclNbc
a7vFUnrzqy/ax0BQK4n1u2z+4eqoQR9FO0VUPcCATaWJ9maC4+V16oGrkAH7Fki+
u8/9UU9ESazZNx1kYBwFZNZcmvlz/nNqluMzqZ2DPtr/++vRNhSHjuyDXzpC/Z8L
ahDIE6B8jYLHVase4pjr3O12Q3oVJN5dfwMaPRRMARdn2obdRsueccUQwHySU+W2
vVToqcyQ8fdzN/fYlPXl7XqGS7rH6ougIQKhlhi90OjWLUIJAl1dHmge92LcE2ZA
H8wLw4FiWgo6cvnfe9RQPPf4CfBs8hsOjqwRrUtCpukGYbKSNZ1SBpK7yMFWpm2B
Nroda0cqYDfzbfwqRqxkW2Cq18FkvZbDHPZguAooUbtk5fNIezctipbfQYUqlueA
/4pZN+YQaCnQ8b4zSIrFddxC5AIKqMyBnr4wgTl1IVzx+6blan4MKAiiCeK30/9G
dMTPoAuTnlBrXFIrvxyIE8zmTbMaAhKd+Saz4jHdc9c08PwpbeXj4UH3tLtQukgH
1SZ/VGCN16AM2dnL3XCPKnQVS/GRhsBk+s2JmlglWY1HX5LErJL9PPMdPtAomrH3
bitCuEXNMGWEFM/pDmui2f6hkYx2RWWXRxCoKJnrn+pDqPySoGaCXA08Qfg6D/Gr
p8ndIkBfmpEHqkZxUEAgUwqj1fFL3yCx9lwiMI2ucRu5I/rsEmdP3c8SeyOHyPVW
evSRGIHCm5B9N/rcRFOb4ofy7y9ELNMy1XzHjef3L4QzBomDvnteQhDuC7ZAMVxU
3QjgSOwb8fZmO35KnGVcOK38j4scoox7dacz1OQEkZzBkJ8HGBJoZoJ2tyZjmk99
MpZUI8A2pENckLpKa+AH5tY4DFpQZ9RvZYLaD6QuZCyV/r6clkUfYqFU0eBj8kwD
5YONR2GUEAgLAB1UqAmMz5XkrruycO68RYGzsSj+QebvLSVgcKgMSn0LzbZea5CH
XeyE5xexwnGuZQ9C7bqdKt3OOIMoXqwjDknz59bqsNyqasJjPYeWm+yJXhPJk7AX
LAgUbFeUKi/uUJAHU0VqpoWawV7Nnp71h72AFvvstlSWqZrOrkNzcxgye0ifqZn5
kn/+6NnkZD0yA317GP9YiKPnojERIB9F03zpYr1t+hiLw6jCdyD3NH9L4VNA3JMH
oMTo0j8ikWs1ZYDydI6vXCyFKNX4VQ6QxSEphRMUQej/8qkrKG8AJGzFiNQxw9K+
41Vxo/HZG8Cg1D1vGQOZhFHrYCEGiqLkpX2tv2ZHQy5GE+l1tlHzFh6eVU8T5HI6
tfpr51Io+5BjoAx5qdC02VBSDgxdI4N78N43zE5qsK2WyoZsEJfowVqeHm41OPYs
dFiyKEJ2P8ODbdC5IRfGqaDaMcrzXN+GauLQ9xYqqYgLB4pnBKZ5xY7Iyaba1Xij
1FDN6IiXKStxiBHUJPQifAY7Ts0ljhAjnjniSHS64fdTxfVe6BzvkagHHFg8DL/O
2RzHCGz7bpY68zVcTJh0mOlS5TQDIwBCXek8xD0mb2UvU1czslNUTGL5BdzJ1fKR
yxfgLmayZtys4BkECvlTvthm3wdiWcTapj5ua7L5kb7O/tzG5CRYvPlxXATw2Wce
+lXuxeN6Xfh7TnEeJb6P6wA88GonsL9oz6/fu9IvAYka0bfgbKT4cQOtX23gWmK1
AhEW5wiIVikNyJ+k0dQA875SysAINcwtu1w6NYV5ILW5yi+tq7sGfm0RdNqls9wT
Xyb3Cl7WV1OkoHtnYlffQi3ZnxuSxf8GO1UEpQpjcpAaqEbBJOF+yBnTKkd7CZqw
htFb1UABd7P0sS3FzlL2k8b/i30/UJ/SMU6qi00Du1CFj6U3jpxDE1mcfL6sBz6Q
3v6u0M8drYplKukBVkwxxNXWxyEHObXThLE9I2XiUUBnfBoMWIpqbH4qRQODYH3L
Vfk3aKi1Uu48Bsiwbp9gc2Wn2ggXHo4QHFLgN/EmCjLBszbK9Y8+XP/ZWpQq5dq4
tBfNaSVofo6AydpJf66+ZQTXgjMHQ0wR6hurRrKmlnNiMf46N+Hg+ZwnN4dNlGYY
sRKBNyS5OZufUsqoVZqZwhP2KD/eCK3TqUcOg1Pu00ciHvtraHZFA6SKr+F6obfR
De2RBNpO66iYEo/XQoPK2avtpOFYoExXVPOaYTJJCYt9+yxyPAw3bvchNnNuQcou
fkYeeZh5hDMfy8zVkliK2FJsTuEOib8esxGEs9vUcFmQXIquO+9CY/Wr1AcKQxNm
9G6xLP3Yp93avuzHMYOkcCr40SLtMMN+AsJzQqpLg5Ag0pm8K1JnbCvz75km+seB
JweymLfhyPcZqhMuNcUP9q8dzutenF99A3j44lO5lj5Dcn4yjpA+LTPisXVPsp6/
rMlknMqWiAx/laVAJ8Xy0iOl4tcH6Wea/zIgcvDCq5OMPpJKyTJxOGtxq9SvyFtN
LPmOchlolsQJviInffuhNcj7ej4GuHtsomTpedA3DYewkg5qEdfwRjWTGvMRv8ha
F4a9ARjloa8sC/jIkLtLBHR7LhZFqPnq3QZInYrF6/vyNQu3xNoRDWXGOI8Psj57
EZS9sXclrQbs5cCtCa4sP4N01zJtkMWmjRQ9WsVdzTX+fj4UgDjRt8OaNb+PT2wR
p4l8tFRBHEv4FzKrYTuKzJGWir/SOVXa4axyeEwTn55BRbB8XF4VNvUPkDh/wWBw
azFcCObhQTk+nH7wK3YA7acYpQ9vCPUfZA4V0iyc+n5OIK2H0zuodiFGU5JQM7av
2+leFySeN6KMo5o9DlA71lo8kBYEYSGdrg/AudCnjmyitIB9MLBxIpDJPTAf6WGw
sa6XdpSF2DCnDX6xYQlXeP+9rrdy5NnHrHYUBrYbu8SrREmfy6zI/LrvsOjBJ1Uq
xPM+wKHDNO/F/9HuaviTJZxdr1nDARH9MpdbcgA0QvRarkWVXmD5z+kCT21+5Kf1
o7m84EqyXWLQvLa4lNToZ7RZnPDJpEO8dQisbIm1Q6ypXt7GKJxO2IluHyCqQlvX
GYbvGX6jHpSVgfDEXqbcIprLyx1+PVGhY3otMjP9DUdERSFXIuJoTHy3cWo929gR
iaNpUhwasC5A+vb5r4tk36RnG7iTv8TR/knDB45QKwU88yLAh6UWe5yj4nCuzpzR
xIhxldyr9jlbM0KDJSta8AUhIMh5Wp6euD8ckaF8uokvWQHhonWKX5bOAib5m4bu
iXDj24eAj6hxsuOP7sZ2Gfol1WPbJXym7I+GFj4NV9rjqLYzSWACt3u2jRAIpVYi
JQDuY1kAJ1YHV+wFcaPWwQT/LApnDVkNzdhXqgFbHs0an5X5UodskPS2qH1S0ZHJ
oyf24uo1buO0WwWNnk13RcnexchezJ9Y5Oy0CKqb6GmxZ7mRSw7yfeIx/OqqxL52
+KvU0r/TnBu3uJkei9ze0U0yYy5TYqAq8j1JBOKAq1Fg0bZGPcek5ywTegSDGLZy
/SJmd4oz2EczIhNEEDQx9J2D03d1Fi2cVKNzo6rpWWUy3S6sblIfygVoA31HMr8E
kHTmOyKNRPyLIv1pOui1yQpguS+GTjE10hEmkIdzA+cT3lUbeqw4CM8sz34pPMBT
NBFG6YK/TFYFQRAMbbX48Mx6xTpDT3ctCxu/m1Pn7gnnOQYdDcn8KlO3VBYYfyvr
5PeM9l3fZsZFjYjvTt9WajA01lumquWM64VgRQnaTw4ot+zUX4cECN6mQbF2JyWL
qOMc2CHILhkSjPCSqlGcXD4GdqL71TKYXReL4Zq+LR3Mi/eu1/2ff8QYs/y/cADO
EBce7MoGlLMrJ8uwTNregnFlKnIGZHIDySO7uxVfUWatrWq5w9FKs8AGsHlP0o/p
ekKXJqHCVtW2Y0tBr49B8PwcQTkjvAy71A5JrfLBfGh1TqXMWzbgzj1v/ZxoD00A
xmTjiWCgg0hOU4XxF7pUeiiV46C8RIDhYCHhBm5MOxCAL1nwf/S4sJz7eJTK8S+H
JTMPZEtrgTddCQNXNbWel3UDi2hrxzRSL1x5PMJ9JnaUBJe0gH7UkS0594Qcwnmd
csiteCiluv+dLMX4o5lQIlCU8Z6fkaHq0qhwV35cO9tk++6Oc4IYQW7gloTyxfiR
PXPMDizk+GKWL9MGio4fw4SmO86psJYaImoVPNe+3psA2vO0cW28zZL8S1j9mhFe
X3kzOXm4IknEgKJ5RCIg5yJL2qBUJ79106pEaH6oAVWpG+XcnbHxwL343v2Initk
AyXXnJkshi/GV0I9QkNZ/LAi+CkoBhZmZKm60lxK6M2PTe7b1TnQ/+1wuR0jnw23
2u8K7M5phh9lP5d3vrUU7jZazWaSOsVR/Bb9dg14uetJQSMMeKwejnW+PJbz5mxB
Kfvby0V6iVshE+wYlGx8Uffe/JsyekRZCUG/CCfiKuG9vUv4MQQf1WnGx3BScCIN
aPKp96wAL/Ib0wrh8CbySmfwKfr7TK+NzbukVFljGPNRY0U/g5aoGLgglq6e+nrD
19nGfCFyxROOeu7iWkPazmqiIQzaDJxKMJAx8bQ9oToGRhT8EONd49qYMBWWW4OU
2mgIzeSVSv8fzXBs3XRV35jDOwIQDuS88Y6ac5m0O0+QVtJyfg4jvhWDwOvXKD/T
HNBmRgqxY9/XZ2L/genW/tddnU77BIe+9HSQ5gKF+nKx8ngCZEBepITQMgx+y7n4
vKmGQb+U30gyDQlDqsAmIBz10gFrOF0u+cFKWLp2tzQgXAQalM8jFp8tFXF5/fQl
8dZZuuH9vk0TJ9SdGZAvCdVv+f0rX1FVazDEj0Gc+p5dQEe1UZ3AEeNlVp5fEWYZ
Jt662aQ9cN7+4ubuEWdpR/AMPMWbTPnkXZXV4MENzRUHDi5o6dp24K/aKXuDdo10
EL1jbOkPCEmkZAeIrrm7jeuXilOkqrlkRKb1WKjnzfbdnCG6qymrIY+8QI6WvD0j
3obNGY9ZqhFl/ts3o2OL9EvGcl0SejAWHIGncwLHXzky/WtaKUdW/s2Gd8PiGKt3
f/hhMik+fDAnI25EHuaWc3uyAvEGAFOibmvOvi1K2CMitd+FF3Ivk+RQItMfVIvC
cbS9evz/d0vRI0KtvohaLIYFj0rYnEUFKqfh139moVi9av3FQMDWIG2MOpWVzqHL
8p7J1qh7GDf3+AAo678reTaWFfJ8WEq/FGErjt1hfN6J+W8QL8cBOW1523QUs2L2
bJ9o9/d/qsEUecCQ3KhhoMmMLnAr5TzdcZBX/ankGC6ivVHKYynzC+lcxKCR4LhP
sGS0NHxJ9Lff5brJGZkxi9CMbC0jM2cCDtlrqVDjC5PvWhpU3XxZjYy8MGG1GCG1
QHlJ5oxFAHOeBOY/fkeBKAXVcBnszmSrOe3FRnRd3p/T+73UbeNoEWavqiE1RDs9
g3v13N2+SkrdL8RCBXfZIRw2EJU71pZoRiMnSrhSsdf2Ul5gAHgMvQ7O5ixrIu2h
DItY6oFXEqxBoCkM4BeQXYhN52Bh3a7VYNDKWtXHSccUKbM3uSMNL3lS+pTrmnrZ
nuO2pCAzmssVsVoFfr7APb8kJkalrXjBVa3+fBidY9KBtFE15qvGvd4tD35TN7v/
MutGfybi2OhmwUot2qKmOIgkBC2zcTI8UgMOTVbuGCyaOga7Bmm3sZgmmbW634DV
hF9NWo4tD4vN1xcOPYpvw+HE8bZyv2aVT/HQfOzt81hW7N4fR4ryPwT34HE55MnO
owv3a6ji+7EnkorBO4E+FuBYKLL3ZnEFXUmuofpJSmcIHTnuBMoG5a8nUqvW8Nlv
ZjaV+VZdq65Nbdp18m878lj3WXIKK62zoDAVtgEvbzHrDWP8u08bBaY++hjzUTlv
+3VNQo1rbD6VqVd2G5Iy1bfQRPZdIBIGeikTAqOuYTch3/rCbfRUEHzXNGoAcFP7
JtRsMIBruKbujHZAuJ80rqrAHou/rBq7euOpv63N9ue5pEJ0PH9SJpMERFJcpfD8
Ocvs0AB8Gc/YFxl8CLdqFMGnGa2B6mhPXvsDhpCTv0enhbTL3LL9buGz2V0s6a0D
G9lDFXSiSoEHHdYxeoIMt0n4ObCNAcxcvs01J2Od6lfQM6P7WYwTqivRZzDMcatn
zK7l05jG5wc8VfDj4GI41/3t01acPWdCGZOPzgco3XV3dip6qj6lLfUu90ec3cz/
Amvn+ppYKwm/e0wl84dxIHKzVMYjRwCXK0VjjUVmuXBUyXCZs5HInvO/mhDk9ry/
hvD+jVo1oBBXMs9ctq/8KN/zbLXRee6eJXpKdqFgf+0rmYMI5bCgPY5w3p80s/1u
6HJtcKM5SPMwQDfyKS+BGCJ/yQ7CMncHgaGy1y2iD1jZ/yo1yhKRkI7N8tLLpFdD
wRzcbERAY1F4YxPr57IyZvChayjzdZx9sMy5wZtmXEwFZF7+OypGhWpu/M4PkQnp
CWtAtyNfPNyIl6q4Ibx3I0TMt/KrFcs6/0tKxqEZ9dCxYlKC0sW7oLTWCq9PIaK6
maPwRuS1yelygrDfNfJfl1LjpU7SXNE8A09NdU0JU3yfA0OfA+bZxTjhPh7bjE06
408haotgFwWPSRr9q3mXWTr/rs5Uq9bdLnCbWqoTKfhcdwaudPqilVcvMcZzx4yD
sn5Iku6ptwwl+KWnPzeEGi35NkvNKJlkYTVfOt59EuAhS4dNHArEArjBpXgbqjJW
oy9C7h20tlwTRIMBsfs6Jmmye96rHNXGdzK5QQDVmA603MQCNjB6P0j98lxKQQHo
09dftZtCLXPOWVu5kVxnI/dNqvDvPf6Q4w/3TQnOxTvpYGYpQQqxZpXgdl4lFf7F
zLggQVLuu7WptKPi1E9B9v5sn35ABdq6E1ZBayztuvgKbFxrNJTuZibHAdJpBbCv
YSY6dtsB6ohtyokRBH6WKDfrats1U1aMotIFfIm75LwuxF7Oks8ybSwIiYipiIMt
w9ORjco4AMM6A1EFJtE29dC4oQtTA3nLDS7w8s71ayt8N2/yApIGulp5qo/8+dAt
l9ZW904FjzDTySo9aTD1NiFk/QcPKbFX4jdILErhytdZMkOs1ePxk1uey7UdAZyx
nys0pkRU0Ibh+QNbQG6+ApEtTwYon8+IdDMdTdGt4F9d63f1tEsZiRTDvhvU/4ur
7W4ekSMzaYpDK37Oi5vLtBp5NMCdJTO9Cn5QOz3ZHleINMmAn3xtz7TsAOUNPrIA
vwt6z9O6Yg6R7w1Q3QbTQLNA8BBRAaoiM7bAtzmVUquBpVWsokCdu+LKaEnsfRPa
nsxQa/ym50Y3BQ7fBuwyCDG99Pjo3fQ4IcpY2Ue5X64UeCXVbycdifpJjO7/NfjO
BYH270cV2kzeU01U/4y81iUttTyWgLQ4fRckHVjjfMM8sUDVgiLaVqD22jMw8+4r
vrhztNEWqmyxG65FKLJqyMFYbVLJZt+I/SrXlMI/v5v0dKDKJ9dtNT3l9bkdtZVk
gC3pI5cw//xF1xtpqS2nDQDSrF9mgagmToHYakkvDU+5Uuu+AzEyZt+8TFT86WL3
29myKEA6HVp7kwBNkG1uqRK+i1qMaTEqRKy369wh0aiPThGdxXejzO/xN2Jjw3OH
F14vbtkCOGf8spm94854S4zx9yfP2N2wH1A9OZo021nkKK20Bh7H9mfOyp1UUoD4
xMflK3oSArMneAJk2oQ8rvII1Fnvs3j3S9jmE5qagthvu7k80g2vAp59OklxIKss
df80kBF5+qgOH7oLrI5+6fD7zV7d1r2IDxg7ZdHSgeNXcDhBDin1tiQ3zEyNN5/F
kEw80tBr8EsnH8pZB3O9Gt4ZDBygfKqu11zhDRExDfG/Tlp3NqFLJGrTMufEwrCL
7CNUp9bStoa7m7UZtCLarFTf/HqHhhTEJSm1+1Z8GbnfyjU0hspjWkFtVodvW5+X
dnDWCVC7J0jDonArYytB/5eKa6xNpKiiTIsFjDFjSTxeIrtli0Ntxj0QL9OT57ng
55TjNHmKyRM2uW/QRST+/G9F7ZiI902p1I1pZWxrQIYDWwby0s7ZZ3gQaR02ycis
3L3Qy2IORBaWQIzdX1RcMR80EW/xoqG3ekUGjp/84nrRhJ/iBp/lCF54rHbv7vlI
py46W431OBv85mgMfnI2ZGC7hiJzqBVxRgsp+IaVGOpZLVeQugPCgvwOFrO7gFcb
mTC+MHFAgxD7g2t2V3RGSd2OsVqPfdIINbFBSQifOx5t5yPxL3qDffWmEK8CaqJR
AHDm/PWlRe2IV5LIOWoXBQl75VZnMZhbNG7q8/gq7RU+ysCKPwenBA68XWVJnX7+
gar+zzdfQGQyrGFGdVfyUEFHc9709rzCHy8eW1KS0DKvEgIACzuTOFxSbEk2DU61
Z6TDnAv8ifGNrVdNlVV+t3Kzg4jVbQy6V3lOqbKdvrz0CAEaZwgxX9L9Jw5PRQ/n
jphXKf03/tLwS/9PrU1AOHoiTdFVidBA6zOgWO9BA5u5tQbFuj2o6E1xLj7OQECy
ergye1SFier/XE0ZrTmFZsDlpNx7BcWS65gNip6FbCkpRYbGFP+HNM/Y1u5AkSax
CvKw0Kjes23dFnT13gow+MpZLhrLuq/SR4ZRgjoaeirSQ148nKwjYTGqgv6ZSWId
ncIbyxdGSIEx7n5fPutI4HbjtfgI++ylmLO1+vNLZxe+SzD5LlEUz117vIjvVcd3
jEJco40Kw/0I54cCTgt6hcluX9rPS0gT8V9kMOdgVZpoEiov88lfBU4yEdfIA5Rr
WoShi0GRh9xYnD3zg0T3TmXR1xxzbfvp6JVUn352RvS/lc0QgwAI+HBbMkyJyj4d
/nIUDK2+rxEAOPFMsfK2QNdNGL9oR6sFW+nNds7ZUXAybxBZqSX69pc0d6bx3rd7
ujct4ftRgR3eCLZynsQOOOcvhwJ3OdDYezOeHVpo02vHYiruTbwXsW5UMtS+80zw
xRwh94g1ArWIJnzoiVZXmpMeQHrhnbazZnZ/WR5DK7nY/gd7RYQVT1k978aN9nKs
hyderFaes3iU29B+KIpomuiTVrvjSj3DCtboRiO8HwND+uX1YLzSHNC0tm56/CkA
fXi86k793xfpLck6639ubWRJ3nXBPmWXF+2DWkS/1hnruEBwSwbUr4ldAjzUEVff
Sp8xDJ3XbDj8LagguQAJQM+lBdH+TS2pdhC9mJBbYnyxZbC8KEflIeCZcGZ7LZQq
EB/xWvd6Z+xPsES9Fiy+pRt+4Mcdkv0m6o6zEZS0isCM0FfsXnf/n1h4CWVTlYmE
PRwZztf5vqamLDsMgMVexUj97FxQORk/JEji1d1Lb8qqtQhIn2wX28/ptIg3tG7W
frXVXuWPv22xyE6K7Kz7ytK4ncYZipuSOr14Qhf5SUEv+RSyOfM16j4bkiEaKhl3
Q0PI/l0i7sqnKGi++N4lAb4qIsqlpOs86nF0aWgMpkL94OPnGGZES30QtMG8J+r6
dtFou+kmL/kMuttethgmHs7+7BAGmk4bUEWAU+OcZMoruA0IIeXdRsq8uh1Yz8fq
jIBMkfzO7RZWiI87d3Dj6QNUxd6bHQ/W7fsEX2U9IdeAFR4luh7+Y5LmL25QY7FR
QnF5BRh7sBgJgg4hfLnBkObPvedzU3TNFMisllpzK9BhgQIo/WlAv1kiGeK0eGAG
1fmHIHYWN7j3rQOboDhqhxfrr0kaKNvyQg1J2CDiQanP1+wqeFXOLWd8mBhXlK3D
PsxkslWsD1Uj/Lu2AygnZjsUrfF2R5eJv0ej4HCTtUsnoAZjLZuBqr+Ct/ZTpFT/
DPjxpJH6Tpb9aN3uemyoTNmrIvK3vbpIa16GMkG9axmRBiE6KgivCRzVpAv5kGmf
P2yNOYw/gXE2L8ABNerG941w3m+9D1ViT0fcEg8K8WGjoW2wy2NBEvNUt346kpJE
cUXlsUgaBkGHhzFqRTEixLsLM96h41lhsvdOBgC74W7j106PFvxHjr+P7juaS6+Z
bCIWiVD82TCLF8jNGlyj+LI9oUy7EROyT2u2pCv8Ez8+FR09hkYzYecM9wthGeLy
B2VAJxPwpKxFSTVcrS5x1Z1KsQ7ZQWp4JS8ykcDZq8fjyWxM4aid7Bc7Q7LwudgI
SE+hUTxp7yvD7kY54qOyVDK2F6gurXM1cpsJPIEJSbHzxCa5Mre9JPGVWFTan/cM
gQD6LLq1Hib8qY181MtGhARFlZSls7jT6NY2Fih6znr0Lhhvg2vRCM0zuo8ayEdC
ZFvL05WqdPc8yjqvyeQRfdsVYhQqn9i8j/Ac2WYe01MqwstUEWreIVd7HW+m/uNC
SDSteKQoKUlzm2m2ydaYwxAdHUiarTLvQojo/TLXWSljJKnBgEMyDRao0zer7if2
R+yOKnanKqhHpRmuaz4FAVnA7FTw5tMB8B/MFtzhgcDF8lI831dSr792QXumqU9d
5z7bu5RD3FfN1CUkfOUF2oE6eJeHuL/oOcKVsnsKWtMaZimEfKxNOm7KQ13hFjbr
Q8tUOyliyvjiMy585po4DC201suS41oMhfcevDviH2JNbVkYFVyRf3/r14AJDix4
AhMel2jht2RPqjDlLtrBwx76qyeLK8KLTbrhxY7ZCT7FCcdu52jtbPXeIPEvhPey
9uLXiQZ+NhjrYCqj711yZKVn4jUSV/ykqJpLRnOPmekTk84GMkeJMPlKY5RPRJW5
wwc9Ao5cmwUwL6pur7HoqygNlAfH8FfVuP/fPj36H6rArtgr0Q2Iu99ZMcXkX+V/
V7a8hvxyzB+MBilEpKBIdbnhYJDqPfsHBGhKVSteR5jEi8EbCbZ0f6oxY+36Zshc
Q7l4GUS8S4wH95BH4wH+/6VZRik5uIzpvyW+uYOdfLWxK64kagR/H6dgCHk8orvP
v+mOM+aTge7HU4Emi8lB6vmb4DLO+caBWj9lObE8GuYNLZTnB2X1F8XnRrsWjE9l
blNyqKRJS8xPypK500wj6thtpLFvmYGMFhcx3B9CHIalLWMxaT1ec897TsKwqqSU
pK1LV7dv/vVbo/8Iqy1qu+4UBS9JVMI6QTqYCcJqViWnuGzELvevatimH4fjP5GT
H8S38E5rJvkzL5RwsAT62udPX2TPrBGNUBPMMfyGNRhYDMe5W0clpK8KG1vtXOa5
nyE/JLGZTjYcWcDFsHEZVSGaRbDfRhLImYRCdhW1FLSL95KqTo4piv0q5VCGrKjt
zQ1b0Xi+gCht1uhnpxskFS/arn2xM3uFgBN2RmCkGtIKnWOdSTOjV2GEUipTpO1A
ed/qd8i8aEdOFcAgliXiWo+cemejeSo5IeWhhV8fzRlYUzhk3sykLyz1S+7dtgQ1
7IbDnDlajlxEczhxIZanLV0O1jJHwhcpqquLXsW5oM7iFGURDYAS4x2EuKF3Q6Xz
8a4ovCyh57CPygrlULL2tPOZKjLsFWKLncoLOE8iQfF3F29QENIglURTsp0IhBiL
7lC2l1NOHUTQyua7spPbdjiIe/ggYcWpSBBRB7qDdE+G1yfizSmMe45vAz40FBef
WSi2c4tAt+BXzF8xqTBk3nGE/MDocGaztVlXHnvGb+tzp4VGpUfHx14H+/VGRrl/
3lrRq06mqrdHUVGDUelrpA+r0XDhZpa7UG9FMSvgetoRFFdiUnRXv1NqDxUsPAhA
ZYv1Zx/27bA1ZW6rywIDdM9S+qap+BeFiYe1wYg33Twlwm5RepSW0NWTE4NP/QH4
tVHs0NES/Jtv57YhmtCu8MyEMXX1XFkzvVIIVsRNQ5nyF6L+5OHaZnc+dqfd7oVx
EVgQbYN+3KukeyZwJ6NyY+YOEhlT3Y0SUEQHj2cNIa6e8w9g6Vqq2w8KQ1OW0PjM
jGvsb2Ge0ET5NlMG8pkRjUzsAZoebGzsqpjz6+NTsfRFrrAjyZFxqVnz6DMGYA6F
FZDBp1u2ABWc9E1n3mJ5hNaTaPxyFWgRk/U5FMYm3NAKYCH9RJY33Ra38IGCb92x
lq1BSJ35EMSD1VewdnX3HQVHD/2K65K+V42fsQozaQ8+X67os42WA6MUkZ8IwiIJ
vo3MY4bzrLUO4ISEPNDPSYu27iMt+w/6//QqAvbD0Nq4OD9x5560V/GqvlzdlpsA
HlKiW+5xVAuxiweOp7Hk0wA8Dqg/AjkwM8Qn46CpX7iKnXlBu1kVmyBxKDCTVOw1
xvWSP5dKLRL4suQRjjnbJJ5VdDE3zLW1gYhl+H0Sik4GgvnZflvvA/u2CxVOV3hz
r4iewprcjEQa/NoqQ1jZALx9MLN4kgruP7Q6F02KbIM7ux2NcGvpfquzsmzyU9NC
PwIcZf6SSpx55xQG3xSMKfyXl+NR8QnldtJmDdOWVwVN/ZaoIb3LpTCqX5qLSnV2
/KFaiv8LMnsAPUmF0K1Ks0tyZyn722C9qJsw4XoubNkRvdNKuSvSv3rv2Tw7IQTG
ieU7KwJw5tl7yWZxJWaP9GmZ+nkDRY33MGI7DTFfsFjwc5BjW2l6+URBJxnUtb2e
1YJRn6ffD+vawQTfpT1DwFM2HLbqERQ4U80dwvn+q56ov79rhGMQKWvAUx42XC2x
XaL+msu2sdw5fZm5kzXzYEAtfq2EouTNovrndD9maokV9whJht2ThvkbjOEXy9R3
xKC2i/NDHtJJbTU5/9O2nf5Ab+3s6/1Nn8/ocFJNMJGnhYE4tBXcN1gvP9jPNIdI
kOSaJHSPASFMyy/F+SLzv5Hkdn8SOXiAfg8Hb3J9vo9tv0vBTixm8NSc6QNcwWQB
NY0Cb2UfIsESJ9XtqiOtOPLy/91DpDfzQVcDicHkqqQhyWGOKRTRI1cdnnypAIsl
3rWZPZx43jJ6otrlMg6Oi7maoS1BhxPLwB6GHh4lQRjk7vsJg6GOH+Q6hOas0eiO
x6+VX+UEipyVIsh3dKHijs8lrd5PiAgNBUO9QNl7RejqnUnb04JBvsAZONECpyDh
JOYEcVlyhZVeb8ZgkjTZ3JeCGtiwtYKwBxhyBbDMi3WRtgXEl6UmKadN3lDWUoQR
dpvQ97bDznxKndiqwqfwx2SwFgEiT7BT+xNWjHWkOwGnKyufKplvS0ron8DtR5t4
5sTCbyxgsaVKJSgJVz0gKuRP0PfyJSsDRAK+prZqnUqXQtkfrPB80rD5VsBsfVvR
qjfuO4lpgyJmNcSWLfSeicjH6D+z9DNixD9MEoaGjhiod5hfL+EzME3G/BtGYV0D
9TCAxeA4HbBNO9BgevLNWm4KfcK1kLTxan67fUArNNH1hoDcxea+TGVE2YjRqgp9
QgTPRbSYelNrRLOxi/OwwqqzKhft/G2kEH7POkrW1T+DuxWP0Iqfub2CtCUq+xOS
eNRVAtTobeq8S5YaQLEWWYee/zndkQ475HwybA7imaNLsf8B2xObT5b5HAl69Gxu
lYmDOw3lon5HCLAPhvglHUrUUcAKen2lbWrsRWwcuNkLcpm4XPEqQrMuC5xnctuX
xh08MxRhcvMyGrUTl/bc0RJ2PTKalNhuTCxhz/YzHslq7/P9BXqwXsIEpUdSlceW
HFt71Q8LNFd1NGqdm11G5PV1qQLp7sS5h6QidVXUzngA3cDROSuvOSGFZMMY1XGU
gbzblgITgc57GhljgNCzbJiiwOc3sl2atIXj2nDR8jwi8l2IP9zn8d868/Smod3e
mMCVXEay0+XtJlxf51ZsWuYkTblnmAByfZbUhbVwPBlC6Yn0kBbaAn+51muOK2zg
rOZlRiOiJFlM/uNfmqOSNK2rNBRERyNAllig9A+B3dZGPrsgEnpDl6oI5T7vSIO1
IEtgHzGdPNl0v090HDu2ewHYeZ2/9/S/XnF8uVftDjS5Ufv+T74V5zA8ldMMRrTU
85BUyO8t1RnQ80JhuDh52FcqLg0j8LNHWy7bbMVcl2oxZ/MuIcpK4JRemAKMohgm
jfxYn9mVn04iXlJJnJHCubt650DQjH/vV1hUR4a5UWD5F6/NDcCsk6nck7+n9L8T
ZcvmLhSzmnjhtGyzvTeXgFMX4NWYI++VHcN2Iu8I9q1/u7/1hDNo81DQRlAYa7qd
z6lGJkuEhi8zYJksNYBEh7Ztnpqo+mF/61AoajmOQYbuld1CoxEJM0sEhGc/19Ff
aT+dvj2Sn7R60IxMErUap6kJ5fnMAbl6Y5Mq+sEjj2dUEjEv8Xy0w+S/I2OskFtk
KHnHTbHKDZhYpd3im600lThnAnYp0GZM+Pmj+EnioF2BXmnjW2SyLkRuFqu7mbBx
BUSI4zbWzvFD63nMz37LYhmSjUE+/RlikUYVATT3mytSF2ngaMqIbqCPGYj85W+l
GCioQ0QC0G69Z9tMfpreimcI4AAcirdRA3OGb5BifW4R/z1I/kYeZdQQeQPcaaSD
DIs8DupKXEKrI5mj2elnjvl+HLfSpnEUtaKFAeVou//a86C7RS/4H7EcHGP2vmVk
LTrMD1GYoOpDEu7xtBr/QUMmBRqO0TgqSSRNSiTH1M894/oT+kBhVB24x4w0rR08
MQNSGuTzd7+TxQjr2qqxpxJU2xIsqhUhiMeTgOPXrf91qgBTX1F4qAOpI4DPLab+
S+iYmh1tdFj4ZbC9lH7NSqojHDE2XK02mTgwxN0vz+7uykiAcINCI1T1mGQfXYPI
tm/PnA+4VczR0zToXhK7URklOXyov2moZtyT7/HlTompdOTlX+AWvo8vMxkThFik
Hp0/2+04QcRvg2eeGQRM4sPJoZ/IykyX1oT1v/EtbZGZOWOaUHcf4p1eT+3FAfzY
9q6tuKuTZaWt14je4BtW1XljL4Vn4wSlClLb5vhrfggiwt1ChGBod3g+ZAjPhxek
kLkIg8AwpYXgu8g/aH8lf1oUdxVNp9XbAWjUkkPflX+ap7WeEUY+Gu4957odsdA5
apqlKxRAsU7BuE6ci0vwM3fiEBtsWL+v7Mhu1PmM/4dtQYwBUsk54B9YGyImLAdk
6xsqBNKNrW93j5+GjYbqiMdpHlZl9uD7tYM6Zofe20dcCetqOXae6zBLEBPD0Wf5
3zoeIRaKFAUk1liNkn9CajbqmPStlf57FZstE5zi0wXMiajeoKYR5/p8Y1YUJZRn
yeHSwVeOg+y2LkwbqKbLEX+5gr14c9rojrAobj9Kcx2tV1IxLWdovJ34LfrWOkcK
QnJUL7ph7/eRj/p1NRBrxpApsptAiPYLuBBxBTMB483VMaECvEXECvL0GV5iamDl
ImbEPqyJ+/OxVd0GgyXvy1XthmA5ocZpqBq5ahmwLD1dKjRRsby2wVXtU9NfqRrQ
WGEFhQquQYX6UqF373sTGMXsECaij+3N+fTJJMbTgFXwKFFIYAPkOei9OxgR3ihm
ZP2vIMnUk6p3pzfLV3JSrw4MxqvqNOSuaVGj4EICNnxzn8HI1nV4zRn6aHp2I3GN
eagK6q5N3InUIkwpeBhrVED/PUIueKIgP63x4vQkuOrRen9lH/dskNDdlX74BMee
w0spGRtSfEHcYmV2aIpLmzH2woMqw6AheFT6eu8yfIhVmPDS9/8YwMMFWFnbIVr7
1bk0NVuLrra/5bWF2Z5aTkOdR7MWdQ+jgmKMZmQsOZkJbS4H13ICj41e4/0IJ6B6
1ztJjCjAq+6KDnTI87+A7Bmazcyp+Bjh3JaSgJvP0SNgI5v88zsB4FWanY55VMh/
Tgwsp9OCypNX0kmSSv5XJtiG9is4ULv66PI0oAn14yBX55DUPgEedUnzrJHiuiqB
B89qN+oiq1bFdps/EH3NyVcxF7eumfmLby8Qm8iQaCvXc7CmxNWrOEZC61evWwkC
eEgFcoapvjuvLRMrlvQG2MstXuoV67584vu/AnpDCis8dYvak9b7KYybJzbMtM/u
GDBKIB0VVYBW/ZMDzh1DlOTVhKuUnxpxfrJc1pWhlMsoWuNRQLoxR3K/2EtQ6b35
/MrabDWaixc7VyAvxChAMDq2KP5ewGMqy3ALy9aMZ2jVpRkuQ3qJ5f5t5vE1bXRT
KJ6n5E80UwhuZARvTzG2rT7SxU2fy9LOH0TtAR6tnXEC31quaX0NS9/ydmrsJDs9
X/f8OUbyoPc+VOryNMIpR7w32WRr1gqevPwxaoO5UIDNYnr6B2yrGwMGukAqIle7
KPQYHA6l2EA7wXJtxymmL5wStpza7O5F0FdyDGSHwyGwDSQo8ClDoIBjleVKDkr2
f0x4XUnGRxac75nmrDLtggW2zXIp0ur9y1PlCHII4NOwVRTJnNDIeezqumXtM3mx
wwc15BSVkxJhKOkT9/vy2srbYcxnUPS87LUAuSBDFQKg7ZRACX9c4OgVMBj8IWgP
pfou2+hIjSX1Te4v1U0KEUIhLFfxuhsgLkYaWHaZp7ba/BH7QyNIRWbZNo15ENPl
fJlkYu1tjrsNduS7AzeZf8UYNoufT4MSV3bG3Re+YQ2oT8ccy59nxvKmbrZTNBPI
U52jaHGKpq5xH5/bzecSDSGLdBYoJOGsASuV01sdp8rsVRC8ZGTfDG4zdoLVfRuQ
RqVJPYS6dPnNqGNOq1EYisz9byjTXKaPIZ1qKuZb0yLg+X/RTKMoL54YFX51LojM
8XERuein0Ac6Mj9kBWezS6SvF2osM4QlTM6URmaIypY2DvkvpiSWibk3HZrNyOSP
95lJg7rJ4W4ZQIthJe+Je83x15WE6xXhIJBicKXHYqbcctM1jJeS0doWrXyH6og1
YsFiOQAD7uTB3bdJUmDv/2g6zMiW3CGnvFbjR8/zkEtPExQRS2Ozi1Nq1Ln8K9yX
z/8TjzbhIfO+t5m+oiFyAqwa8LnG0Lca3LzGMK3/AKtRr5m4agqjrT+fNQWU9oDg
S1FRXTXwjY7M/TWYFKEgajPBSAXzCWxCvATHJdPX9R6T7oZerhEiMVUS+QztWYhV
ItXO8mdngjWzeZXegFkXeF/0DBQ0w9UPmlSEpG7PLlPD2rKhzqdw3MQegzNqockb
ROuysh5NQQffDHCrf3RmFzqkpMFiBm7IodyzEY2VOfPbnM2ropmMsMIfqHih9/En
cCkQk1HXsdPzzJOT0ZtX/91IVuKJe5rJeDUIto/XudGJ4bMj1sVLhQEdjQHPxptj
9FnWkrPr4dHnmwj/wETBEAtMrucu7+rsXFBM1W7MC71ItQ+v8i/4qOXukx77dRxC
3M9P8AjdxqtHVIyGYTYhyEDkukofZkHMPGbshozypXrRKwxUBxb6dc/btu8iVr0p
ddMAGUuj/VR1UBp7dMbk4N+bIaO3iyCeiGgJlPmXAN4hw5VFWn6r/c2vJdEajlG2
3EPnajuWPgm/dBxtkh/zHUwPAyAh4uw1WEpi4zFJW4dAwaN6lnhEpPw9LVLQIwMZ
KhPIqPX+Qn1AvfIOkp6DqcmY5a/Q1kG8hDVv0ntnN6Be6lTiahs5nqsEvznKk27J
Y07nmdfrTAsO49tYBTbGqhwyE+vBQ31eYdbN03LnfFW5F1iSR3/0+Flx5LBz2aD8
3kOqhnHa9i/3YX/Am8epCbEUnhJA5F4082djBfATJTgHYvGQWptytuLpHsdz0x/Q
S0LYnVeX9+st0KZUZsQcNtG5O1EEhMy4lUDI653569o7NtWLCrI/q5ibf1TLJwQi
hAOpdMsTb5WXvjdyrNufAgWJHVVHwlyQroTkjvjWp5mNV+zWKFRUzgO5ZQBrnZUS
i2IsPjwBWt+OL0mHCX+M9OPA+juLc1fSauJQPSbu35MZFivQzDkoBo16uX0fR7OV
3XiQL9fRMBZEBX6ALwFPMt7clzm3qb9lMPsxUrzDno8ju7qkZylfPfy0Q97m8cCw
rfMByT6mH+nKwFlqedJtyQ+LL52ErHWSBeFAG/kPoeUtOSMMgIe8Sbx+/Fbv87hK
XPy88Ilvnsl/oxXwZfj9iW6I/wEjRb8Aq+9l6vGZLewhidAjggL1hvWV425NJ2/8
98/lUHeNy7jaB/oOaBufHeNGO585HufIRBeg+ZV/4ZF+VeAkEVSeAWFbcXPDKTIu
GEwxtQX0N4CsEeTIhNATDJM8/Ru9QMsngAMpFDDM6i2NSC5BEG+ENymZnZgyxTl3
/y2vGLcyppX5PTkGC2/IPmhDG4nKbfGPTNsb2yMKA3V2t8EJqLpjAUwzO/QyiVLX
N8zorO2fD4F5opUgntmYwsPXYl0tIu/LhV+kiQyP4jxsLJbeJ2d3edqg15eiTwdV
V7/EJvSkMwe9hTfb9eykNRScG7D03vsTGXHEfx1eD8fdRirgtnRPEFA84+vj3squ
rR1XcQzG0Cn0XlZ9PZ1DxEJWmvCApWXwMQP78E9L+eKhPhKs9uwjCjiTDioiodQ/
gA2myWmA1TKWRF9c8p94e1R8himUVu789p3t7DEe3ASxOtqvjCBUTsSwZPump97b
RKHHPo3Hx+5bD4Ewgf087RPaKmrTaGGBjlos7zopAufCDC+NaRyGUzekcg81F8ku
JnZTQgvwTn+fXOn4rUEhEVVixW4yJTYcoVMIFeLeQxEehFEhoouFomzi9pUo2ypd
Tfiz9ctYaRYhu50t9SR4AyuVwjTBXlW5IgEvhZqshpWG27/Mtn+ANhQ+bSk2+Aw3
tK8dlpFZBxIO1KLnNOMzD5/VyGhWCP4xHGfoGV4B7aLDfITeSb71/Urr0njBB8tl
HcQKqcEPmejmU9g21JwjMgn9kUmTpugpeMMnHsziIBkokGkYEWG7VN+0zZeWeMY5
XvtkPQyRsARiJqBHGcFlRMXQJ9nUB0gGlUZa/4+288l/M5HmNW3essH8IN5PaqhJ
FO/A/TwUy5Ry+g6XXlbOtAYmjHrJEPgZkqmwBcmnb/QZUZ65/+qDUohDQxrjeOxm
wlJCggfytSIwjzEWRKeZsTIQyKGJbQcXvvmzZoEdn3Vy3m7dcbt73D61dA27G1Je
6xq74iSRpiYLvfu6DA8p66p7SG9g5dvW59v+nB0fOMcdsQXz5EvuVtN47i9P/pAz
u9zFvaGpdpz6CU99jrKi5sBDqcUDt/2sxkEDWU8RJ8kPtyd+kjjlLkuRunOKSdo/
OHtkECwk7uXRvyfVtTsmpmE/D6hiK1TS3thJ0Z4Bcz+6497W87chL6ge6I6VgFuU
ZHaAm2UCIoFGIhXEkzABvfhJZAwvS0ETPhZ1JO12QafyCjJ2FH87/78kMUUuzm+n
dlLYfDIOuylbBhK2/cpmxV99h7TjQdMMjrQ4CJTQtM2B1/MpnfOS+CrXPpD9ROvf
tm22LlvX+J9EqL0Hnuq2RC0v4WtZMV1thxljnWX4S1rubpiBTKNrU06l4xbj5tes
QIu+8cMTFuPz2fIti8JUCm3i5uHvji0wkhiK7xLIYVdoWx9UqMNQYG3Ps9yJIrBY
IA0sBKdIsuomNAPnkrp5ynXadw7t6SviSP5krHWrKH+uG5hcJcNI1eW3OrApWW0h
QLxYG9W1K8+2CUlIIxZ1nsQShgUzhJyofYDYu747wHsy6W91ie7LrZpByVu8mwUq
HcEIcRQbdPPdXAuIisVXWGqGe0dLn94EipRGNwnU9gLHHhMXCQO4pdPcpZ1esCR4
N7w4ETemyykSZapA10wXrPOjke7UAGoIoMZWcpeyTrfUIbBRUeTr9kHIftS2SJmF
1IjMdtDBZicglUpcFkAYc3wzoaVLkTVEBqEYi7vMVkX+WRwGFGWPsVSW6E+A429M
o2RspvxhHQTfmLtmYBaC9UihBZNQT0cXtCiRlV9vkKgjUA8Ko7xoBhAgV9C0AsBs
yZQ4cTtxoigFbbjyMvyDgnJ3fXIMkYd6hNM0tOqkBrw8DzzO9jJakynTmMHM8OKs
8HNKGsDvnToYkQUxhbT5dyPNHA+Y48WVQ/XcD0Nk4P6V+jIiKwNuMeHibcF6OvPA
lxxZMmYk6SbYV+5hF0NyuQM9sNS10lkgCvV2US/w3THYPyt1v0JkwF5nxnIVh08f
RbLuhRrPIKMnPfeRpWcRehNp4IT9XAu7/bJpS48tF2ILI+38IgkYCFdWxo/7JEi9
9X2rFpDTO5W0pJLxkzYwEktMJWwOU11oU4u6D7Es28LD8Y1y15AfqjTr5wer4eSn
xi4pHgdHw1+TfuC6OUzkkjv5dFk6hGtKlHvlqHr53ag4M0JOrqRTmZccFtUw4g9d
AUL4AgpqoJJzafGZ0NeA3ZHZzFDeQI6u8DT703ITJz6sImMl4h6eW+hHDlI8gW/G
cNMVop3yu8Ikv2qWYBMwCHhaa27lFD69le81Ze0foiLT923B2St55bIzFSGX60qv
7tAR+qX9qCVcZR8ZbqqHtxTad7FQkhVcTwCsCDB0ltv9FGQEx4vd+V3TlMOFkO2r
xVM4RIVdCManFyCBmw5yDxHJeJOzCPDT0o4wtvJcbD/TT9S+vGrFQUAGEFMqsAXq
lqGPUG/HN5xDexrffIjWXCRJPvKXYtJItwpptl0rq+3CC/so0uAC0GBkXOVToWGC
WweUz2SF71+5hHfWP6FRkldZkhhab/iaLq0uLkyIrj4xS2rh55CKlPoMGrQH4N89
NCG3Oe54p+Kdg9x/C50xjlIc/kuwXXhaMJYMFt1mZ/d0avxUh8EkF9oeFFGaOLOR
JzCWhtemRgkGScEc/K7sdc+uKeSpnGOrfHgVnm1qttjc0+E8uB7YDSedTlMcFVGT
+nHSuQbeePt8LX7MXTsa1yM2T6WpFeRDRcuWNIDOaXaafna6uuO45N66fFTxbJ9y
7pmtGyik48L+PuN8Nnq6NYOT9amZxodnRT4pzZu9KaFgSjaC7pacUdhdWPJV2yaN
kR9dVGKnvZuJZuExvAo/ZNhoZ8By91TGMdvmCGGJCLnjsILwaMN2g/OldcJ246vx
+rPkjDg50Et1nl3Gb+lx6QWeaCjxR2+02AY2euSuL+Wex3NIS1ZPBwwKmmY+lLKs
9lCgZ61uhgRi6wSFhPN59pIXkGQ4XwsbHnnMX0PkXSGgCfnlUp85OyaLTJ7W1kU9
RKhRrwXceNP/LTO1M5jQWwFsNcfLi9jBItoK9hdRbPfnlbwvcdIsT8k5C2NQDP+i
gPVFRRCVWT9TlLiByt/eKSSHM+ymJgWlL013vqy0T5eG4G7CXhsroD/fSVngmr0j
sNUWWt46yCEJK/hArXBdRBeznqW5I4jE2jp9Di10eQ1fp7HIauwyWdKhu9M+Cv0W
XGKkzgSErmL819AIk0r6lmhLAcvnUi78vnh+YEFRbr5kn7ObPDmVaU/6U6JzDlq+
1D8E8l3FW5YgbValyacOXH5ZCpqj2L8PRw7cIX6YbWjB3eZD4UqHamwDWev2sunH
XKjj3yPqO3+iWv1Tzif79MQJdo8YOED0A2xypyJYQuaH/cQMQHK8ZRfkW+RVBNa9
xEvMrk9wsE20yPrJCpdSlDWTCcVTg489RyBYpirdIwOca33QcPxWdzs9MFYHm7AK
HrQ1WdM1t44dTD3HpsKbv2A2WVo5/Fy0n7lXgsO2qMAIDRUNUwKaz4sIacshhz+t
F3oze1LVm1FEITt2xB9X47JwyiUJ4x/60EZ6QH+hKroxYBBP52lg2SqBN8LsKUpK
DlUwd2ngsXi+dWpGootFZ991aaW2Sgk3BeuRdFDMyNB172eDWtdPQtM++XZevpJM
xBECmf6K8wB6J2ZRlTTHjXI0SHeRY99wQyFfYHekUJ7AUs4VVjacRKyaT2QS/P7I
yvwnLUCEdzW7C9m92fAMB5tDdnv4inINtjE/YR9CC685dDKzlq0ynI52foY04H16
7+jurb8WSTp0gCMF1Un5V9NoWYm6b/+iwMWkM3Iw2b8gseEd4vIkMB7g9sjYvSEZ
oh5ZoDwbN0uMtxxb4llaRqVJNkXMV7mG9vnTdBsdm2tM/FZ++3JWqHRCUi4Ii1Rf
HZMbv00YdEBgbzK981Sb4EMWjkBi5R6uT4KJsluaxW0krlGp23lwTWDkPUSiMmMn
4bbzsu3jlyTPKL9QFm3yqi9h58/pX+7rAaOz/OJjO9vAzCMwxUd+6vme7s0npskZ
dAWGJ3N/w59WzNhN5fTc9/TuZHD1gRAR6c0v9PTU9coAuf4lv+ziQA01dUqlZeZK
XOuEfG9O8YN1a/FK9a3e93pUCeccDlaJwiWo12WnggnqO83atMxG1o/mDXBuN3aN
7Hkah4qblfTHcjazk3ais5KJ+Coxlw3WIWj2XT+zI0O0V/r2z0bIxOFZtepha8TP
tKQvniFjXBGjXtsqXWPG+mBd6OF1TuFzyT+JukHW+k5HymTDoEpHUae0VxuMKHPT
tnlDMmg2HUgIp66rLziv4dcCWC2WN5UheFoaColZh311iVluzjjMVnSG4FltUAtk
8bKQCuoE5G8SjoSA9wwGdktIIGfews4w0FQNRpYH1MN9l+s4qfRR4GgchT6cDrS7
SY5HRwsZBLn+PqddjMExo9CirR6YdFFQQzGbQRgsErpIEHTlZ6BHiOtBhB8BVSsA
H7xJfwdWCMJ6IFLWO4dxvc4539dMnkvtuxU6hdY1okIgl+J07Tw2NStoY2fRyVu7
L68sui5s2kNbaTKs1U+VP6dMG1cGRRU+Ah1EuF384Gwz1ewXe4PRAYYsKsZSrT1C
3gtrA9ezbckVUA5710pF6Hjhqoy1VGmVl0/Htjvn9XUBTR1bUjTbQASK5+7dlmSQ
LspowNybAMGdTiHd1Z1mF8seSQ7RcqMz0uMvXlsQd7A4UkZpGur33gDe3cDYfiSz
/0RUKDR5XwhZWxFAYp4jReNNJt3T1Dnh/0mg5R9S6seeLSZFpU2799RkmQsULO9G
cM4KdCNHBzMSZHsbK8+2K6LjSfmMjZ7ji7TByptrfTb3Y83It4QXfguGaPtMTPsE
yFQIf2QLLfvJXTGtK4holmJ1VfA7qIY9W1Z5/SmcrYu69v/fRCM6CllNpSfVKjDI
Zvk5gZmu8ERlRAsZkwKSioleRaI3eaf5Dz6RaITs4Zu4INR6FWE7YD56zuDoLiFG
y2sxDz71ONju3ils8lktvgWSY7pnsRw9CfmbBRt9y9Hztd3F1YObusiLoOFvrY0g
gz+xK5AKJ0hhyyU/j/Nvn6Io0l7H6xMxtNumQQ2jr+9ZDsrIqyKPU18en+9oYRlL
mi1T/1kDQHl3hT7LZmnCQdnafcpE6Onbu3V2J+A6V4ENj8tVC93w1I2BxInLghYY
VF8L3IRdzx8QqjV+QbaoATSuAl4/tQpMMcRF3L/uFMIMt57ZJFMge7sjK3DHSVzc
DvUBH7tVZtobn2SQUdZQ6M8wgoaPP9b4yEqT7IlyKZeAMHdRrGEy60v7BWEqxX8A
rNZrYyF52MBmJz8tDfJRcnwVSGnCCpiQYV3xFgELwN0h/gqYj7uJjXEavuCvOwDL
q/Fltx8x/erRWWAY+UOEE/9eaY6oIGYyjsXxPw2ZjkhXsQlm5iUh/sF1KmX710SK
qrpBrQNlr4XCNXRew34/w26ktXIScazgIni0wMmacoO6wOmrgVokk3LoUwTJdOI3
OZFW/yFChOHQHk/qOQgpXabSpCjlN5xKPBhq0/N7egpk/vrLUpUTivoYeuX2noYY
bAfx3JFZSwBKmcTq7ni57/tFePRtDK+05PFFM+ia+J3zdDv/SYxpxnOwQo1DmDpG
CaYuBFxprcCoJomGPNmn6/6ZQ+YJhpSDsJ1OjUGKHzcckyczaiAc0XtRTJLP5N4Q
OIVOHjcUKZAysW8OrE5j7X3UegnSver8Jz8dNg3qWoSzu5uuzTzk7t0ByBvvltHy
tCS5x1oj/y8Zmn3UIlLrtGhumvkv58fS+/1xtyA95RLfhuBd1EMrEGM3DU428aj6
SIawriSBH/khB6ONl0roapvDEMKCtAQfGwiec6Fkl1mvjEIHEXTOQz7T8LD8Hj4E
/R9OthVtjhZXhyeXrhp+CabHpcDXhoQvzmjWZHyqzkdUZ/sRTQp6LALxiu1k8kkK
Te+Eqnr2oAurZFz1coPPbhX4gYrjtUv7ljCb+7ZUsTO3cG45FMC3pDDOwcAMz9vc
XKCDK1Kfby309w6EKTSb7FdqY6WfoIoK+R4+8UweqU3OLfBhT7FZ0unrKwRVfu2c
GLgdirpEfP6iVZWy+05wbfdrZS42RD0eg96088avgME5Dr2xduSdITeGCG1dRj8S
ma5h0/qcasUSIlnXxsF9Y1F6va9Lkq0/rL41xxekdmpUfSKs9RtSW5AxLDQVw2Ou
hLxFwp1l8yP+FaLpLuw+ZNPOWkNe11LHL/WYEJwTdvTDJX84CUcw7/hZIsBZ9kVH
ymg4sGVSUZSROXmKImWgkkHyRRYyRdx4MAScIT6v13HNW40UVZOAEjCCMxMwDGZI
Wg8GcFA7/MtaezimokMAcJVNvOVw0hAJDJ524Hu2RM5txfkXkj8lZhz6ntnqZbtF
BGXzSl6pfqPOgghU+r5/rpzUFICqBeaCMTPUXFUpR6ZvBHWOqe3wofWlH9KCwD3D
48TpatOqGGPQND41Ht9zmCdCH879LM8pY5dYB7WnI+rAOfN5cSwqtp3B+ou7uktU
G/ZBQ7q+eWWjW3vndZlMgHHcT74Ks98Vk7d/zhU3DJx7Z7fVEdadDB1+t5YOwzii
n+FGH2ypfqILJ5XbZEjvzwxDhf2O/3MQ36AMZUYvq8WI/ZKBuIi3f+mwcKj+QwBw
zP6mFpSQwgnPF+AaXHv8sBmennY3rQ7V2Nh7CXi4eCBoev9cTbOfIMnZ7/ZphZaZ
b5d82V7a4y/1Ci+kxkGWX2jHzTSvqlTKY/J6ZQksVITg2uHmahHKEsWQYXQ4RqU+
e0Ylr1NhZEjCuuR/QmlvWaYq6YvQHUUz+jUMuGITqJBhbkP+aG0gDdVeEnVDr1+3
k7mVw7CstWV6U7yGNC1Z1dAaMfxCXeSCst5iZBC7vdfvCfiI1VdoN4RRETToJrvh
oGfrgEbmM9hXWu7qiSq+xa5hK5Wojk7HHev/+D2BUzUUZOvUmFVv4X0nrG/FAmB2
ATQL/PwYxODOx1RSl6Tq77MoD1xnYpEJdu8LJ5+Oy2E23/zVIFAHGUUvZgQlTbPt
0k/3RI4vPHIcRBbf4zXrSPOxRd4Ov08drTQQLAFXusRNss8jrd4g/16H7RfFr5kX
A5ZOdiztqrhqtHeyz9AH7HFrRKJZXTNyhdgSiJOJUu+rmFlTbUliIXy84RQnVZjQ
mAjKSei767oJKEeNNj5GvSLgMdabCZBjMA/qsKh3GCYhfctbRiwv19lVJACMF5oS
`protect end_protected