`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQMPUn8hJ5NkADzHaDE1+rdt5YMRGZbKYq+zKXRZdF6oU
tni7UCUNnmWP3MQc5epUQzxVpp+S/Z+L5y9FA6TbgyUqBUWbyHar37pxP60azOtF
wEtAzsnBl3+LtHVCwSFw1ERZ7TC1zIAAO6hRVklGtk0STAcXRIs+TSvfTT3dxg2R
oOmHaPnLPam3O7lJ2KNGO50+ka8sg9DC0+1Nn4DcFs4NcSNsnHweFi/9p6Hzcg/a
RdTPJewhxitdcKQRzlnXyzofAYiVaRMIGa3oChLj8X6wI8EmCMgjxGO4yK7QAP6m
qX4KBG062ove+QmHkgWKuq0yz85urRFzzXiunuD9Ek0yCNuG4AoFpgmwtN0de+sT
Zlfyf2kP2tFftNqsp0CYtMI0/1QDCc5pnRWRwJAnZmJTeMJBdsE29+fwO30dN4Ss
l0HQrhzc7wBJzIFu316/fyF/MOo3ApBoP9KcbAZZ3P70v4Hm/5pfrEUtzBqI2wwu
oHmqsUfDrnWIRaxLLwH2NQyBIDuMYfvVbdJhcYOuOIB9mWir4d4lnyEM1tp3iQn8
RFbAaFHIWyjRQF5EEPrM0XiB4/CE/K3l3iT2q5B9LUbYDOywCQ4JLYoR7lCgNxPk
BRUeTL1xMJghPSv8ShWY+ZfwQvA1JTTiOmbX4Fa36VYg9SfMiQRlWTq9cdMMUG5M
64hgaGpmKm941oC4EOiXEnZovhd4ThdBEI2tOuT1pWohTPdR/HxQIsg63VvvqBv5
JIz+i5VHVqJc5lhEeHyG1z2cz06wTdI+p2qTxP0hS/O/I/vl0krfK/hWULJyIWWl
cO3OB7fonjpOog6msIP8LSXk7jgC9u47LFug79+RoZ5ea+Rr+CY6eephv6XB4VpY
YaWs4pqGzNaf1Pz8Au4bhiL3I0WeKbJHBmBYqjOr26zu1m5ACHVOsOd2ORL1RITL
a/J9UIQt51xkhwDiOtakoE3l3zRmbxg/lc+9fYRQVj7kKleEVRejTITVQV9RLJrk
AtSsvDx6RXATGDxB+DIeE7cA89cVl9F5+cD91LB6kX/zQ086gUY46n54kMmK/dpF
axZHJnnqiKJfeYEzn6nmR1io3bX7v6fFfY7LkBzGLAktb+GOiFT+Y23SG8HOd+pn
jXSkKjdJzLcyqoAWliJzlLMvm0Th6KkimaQQ1VMXa7rWhbqP2AOnVS0W85BJGje9
cxsUIXgC1sDWr2GNx5pJALVPuMcR5UUYCwf4P4dNOJewAfEI5EEt1Da1mm86WM9J
l1z1Z7KBjQU/sUnA9A8GgDz1V5jxQbCzmnz74mO+sZ+WyRIWei5UXh2W8Yl/0muz
khtS9B6yRWBTllRDoIlAo6tpIXVInwPresZTwXgJkWyzqvWDI37nhMus0nIwFiZ+
7nzlSzrDXC/Cjazdc1VW6RjafLvnNx2E39BUknkhpxfAm6sOV2XBezi4gB79QPu2
nh3KGAChywVp+VNLeewK/+o5UVo+TaXINKTb4vkKWFnaZiYAmrOcPa/baHPCRBH2
FeNezd+7rmFB1WfGpn59e8TtacGaFZkXAR5fCs8Itv7vwuy/evNhogOYYaQ1jsTF
AicnPR95dyFrdL9ibsBAqWyV5Jk8GZL4xzLVUUML11YCjuDj1A7brA/Ui+HaWvPN
uIeWcNjSVJWGmzZafGKlYdnxBZhBTl6c7BcvbSz9g4HuL9gvh0ky6sW0hlXNJzUe
lsrIa8eNjn6bkUPLgwsQmWrfgmMfPLm6JB9F1HKRoaG/PSHW1Vw3tiyMOZXzsFFq
ujg2pDfwEw2VTU4woqZ0ta3l0XeSv/c4+wG5OZS4T74TOzpmmbAjYUCySAGmv7YF
6KusEPkLLhcZhZfjDLhgGS8lw+lCMCv1nG9W27dcTBBXeEDe/Xp2ZjReanq6tyCq
XA4cQnsFYYeCqJE7Cmm6e6K9JZDUAS7i0qg5E9dW9D0iJ2STrN1U9L8CXcLTCJTo
j7lWiAFQNes2cAJXwoPHwuiVqyCIiPMxnSQc+mcnQW0vX076d9LKFfhsZ4yNkhRv
AAq9dP1kcrztzlNKD/jyToQ6joAiWAgnPk3YzF+vOQJxfjHwpKLB0RvqnBQcrSPR
olEyKNQoEX4GzzH2a9UPSqnE83RjOGQfBGrs/YaSVRWIQ8bu1OY0oxtci1a5f0Ad
+hXt49suGmS7Ja0DUJKp2dnJK1cgmKWWNo0HnBUs8mi7NNEiMhwj8NwdPYNhJ2Yk
SksYhCAidkXj59G7qrbSSflQq5g+EwrTOXBNluTHIpybhphWIUtJL6FKwZDMETZ5
mdebUQ9ChifNItSyrcgOBMxbE2HD4WLFo3yxyzjZiu2SOFNZZtkkT3W67776Gz07
TU2hEtaxAGF0DzJ+3IObC9Vm/BGKWifz/uE2UoNh2cOJz0cabRLQBbWoxtSiAGyt
L+wCa1/on4NUMG//w+sAgL3YPnPnDBdJAfg2igz/xlpx5Qm7DgXz5O+WhFMLQv+q
AkCrdapyclUsIgD1M4Yc2InUCfV8aASRs9ZJo1Q/whtPWTwVPtYNDd/Wot3o/p/J
uhF6D17J+M3PNBBMkFhZQElmxEkuYyPY42h1MfqXE4ngF8m3ss+GQXJNWw6LiIxM
Xuy4DsIbOacoN/bODBJ3O/N3S61TB4PSRSDCuEfdDosRgPB9ZNP4JpXk1N6T+BcJ
W4VHNiZvcrR77kwnga2AdShjHmhHt6toIa+9AZcAun/hx3HrPr0YL+oaT4DL4l/8
QU49sslvVQ3KReRvwV2RKu24k6q1yAenvcGUnjheE1aHzb6VnFzrJscFpt503tKa
XAvWg7bfFcIC8wh19t+ZO6RhEFUsHX+0IjAh/PaVgDqXbSr/NVtai6wTQyJnDtbj
1givrUkQuAL1QfDu0QQ7JA7smieDAD6rrxG4WlR7+tkxSvLy8hvFV9jAxB0JjSpY
AFKNEh64sMZeqH9t+it4N3zy17w0DbWmo5lQZz5fW8Hz6WZS2pPIlxXE8rDt2p93
BTrBN3tB5Snz1mPLgbgBrYyqQ3Qz9dAvy4neVpVTeJBEmmjGZKjEKzoO6Hta3GUj
4IX6Lp/DiF6BvghC2VQBI4mUuiZA4/Wa4SPnEGaBI7nq5lpn3o0LIVcYp2CVxF7n
2K1HJ6kloXHX8qnVhotw+nUpPXL8AczG3301jcn28HPCm8f1ozCvtoDAznM7IOo7
Eu+pX4b7upea2CBEL5/hu2mItRIOOH5at1IlPC5g3YE1sIx50qjYUGJ0s6HBIj8r
SN60wKsqEjWd8umIV+0PUAvzLUk0u/gUEO+7tIUExR2YZHbYCd23zxZdjHgJsTg7
KeoqJFTEZb9N0IW74kwVFeDp5Ek7U1BhsGk+x+jD7ENMAY5ctLI5nScvxvqHeuo+
e+I8CKnCQLR0ANQyJElpoRMOrsYMai4wNX+Nk/CJH5GOMXMvHKTq1dmJEefPf84m
CvZMPtbF9aMTi4ZWJPfWsa4plNFRxhCWiPnTxrs88PGd5q/c3rUHVfaqT4879VVq
orwnRt+PUpuqguZyh3+8KZqzum3hbOxmB4M6ClSYFz/SKELN/hKfdKuoGygFjHs+
+74CtKTRWRT077chaJm/gGusD2pwgx65fksOdF1WeteFnP7KCWfhOrwpW06cr2tL
B2YO6yI9LxAIrI/9usFPnYdusr9jqtA2d9dUWYO+u6gbNRlo3ajSDqdcm3ZP5Z3L
/LtlFO+c2CUggq2DrJKNCGfLszKuTY9lgxk8IG5UkLPBEynILdLaqNKuTMd4tEoE
kxpG+e4IpuCimqd7g5TKtufH90DTiyGlChT+FEjEdjTCP+1IvCrc8j0pSACw6gnS
rNG7gKcilgTwsiaD2oUt8/ZR5EdjyAFLHD0A0p6Q1pmYN0aNTCOONiJtimidl1mk
V2nB3b/OVOoak0X1n3jvv0ZlS2OG2rlI4CDjh8cZjyfssq1G0zX/OFXsJr9REu/T
JGxevw7EFyWVZnDJlJSq+G3GhViqNjkLxL7ntwMY/LzWJFoUQWeYHYJX5WQMx082
AZHN3eu4G2jZRe3Y6/XUyrGttWdfZaKpXLlSKjNWTf/IGkSpO4l8XybTwrbt/g0j
I9jvgxPk4rIAp5LePrd8aDOYB1bEJR0TGaEnbW+EOimFDgieFN/sZio77xvBqkN5
aOgIGUxkSM9TEtqOOJx079fUNiijm0+Pc4P6G/QyWO4ejbYJCNUTlYWvFiNl9p5d
KURBoovNAajCKVJu9Tgu/EQ9adhn52jE1ADJt/vhCnVKmzvxHpCuyGsCvUQspbNB
4OzT9FU0QJNp3simff+LjCXgPpQMxJ02oh1DREHCNrTqMi2vqjd/tkmcafjFZVvh
7bzb9/KKTcL7E2iR8x07Y0HzjMtAGfOQGmGT/X8Wyp1udUwpIk/G/+bdrjYVQG1L
hxKqxeHIFcEDx+HF18IWh/DBmtE0SNhgyBUX6Lji/yf9PCPGXr/rXV6F4352xBDB
+lP5tJPrfH6jmj7D2vd6rBEjQ6Jpaa6zU6XXj4nqUycVoYyL4y95tsrMvlh5biUX
gZ7BLysg06Hbn89p9ewdguVoxYdn47U/vnbknafuSWdwlqkNMyKzLtTilhR6deL1
5UJsaA1TXRnb+C2oMuGdejjV8VAJZknUNsTFN9uqUCamH7BVbDbgmoI2kPeVKAzm
UFNbMZlQBEm8ezr31mtzx9isuBkiOCFW3fchszWtZDxw30MMfj1VvHPSpnxneJhF
I7d7kjx0m5DbQadKYHm73/igVZVGBly1bUzmWQNhdRAt7xNBHAFbaGLrsO7XoZFt
qHQhWB37H5jGgyACeSW7LX5s1h445OpZXEQxAcTV/SPWLGQzy5TyJn4CLDDnJUAr
E+ZjD1WTBic8Vjsmnl3wtbjwwTmTZPEwJ7GOfAg0RPeCsRXUNbrxKI5AslOdv7lp
iUFk39u6Ie8UXTVUkUva/Cl2YjIVNFB4DNZuwcX95ZV0Dyp6hdY6+BtIoN+uSlfS
8Rlvh04hP+8v5zBFHnLJXxVwX0RwLi89OO7ze/45biXEAoBWyv4ROXp/oB8D9lUg
O/YmV/wm2MIvNGd0Zzs0vsP7veLGcr13c4kJ2DXKHGZWSFlyNBbAeCyu3zxEl0IW
269S3JX0CHmpBKe5ErXPgS0BYj/A+NJj45tNs5t8x6QYVW1sPxYZWoW5zgQdMZFg
D8J83t/THsGZDeLQ6xSCRQKahj6YgsjWLROlRWACBQojI8DpJ3TEKS7FmeY/p8Gb
jIc9X9jgoAUnI8gJdGUkwwnun5hyB/eYLYtphWE+bm/fkScDAvv9fUktagPEe09y
ba7wzFd+0bcyj6cl30YMQgxbUUXAaxyT82nhVeNH4uNuVy5ZCStxqjGnhemqnhQg
Q9kvxKqMjr9u4EWw5RZ0PBfcwJn4tLGYjfsyRK+sKg86W4ZEih4gnYfNN9n4fiek
vXOGRvO6PiF0pFcCewMttw4/sjasHEIJ7rN01TxWdhrjZHDi7tgLmoBD18vynwDK
fAKA5jtPYGTMHNAyemVsNde9fSaCmV0d9PDs6WW5mG+p5mxeZp15en0ycJ7k2W1j
vDfMC7nsd01pP5GA4+jQf91w3qIjQ7PBr0ZXgPceQ+j4B0M8H8Mva48iMrhrU028
NNSOm3DcC8aXZ/N66rHvQyY4ecMgPQJrUoC1FTjw1aE/6STPPp87x08pjUISUC/V
5i+GV9+4VHJC3QWH/Ehw11z7AicmwWIpwwTfB7/gBxcBKXduvU++nWuIFS1Kyo6x
tbh/QSX9Z3aoMBbrrBiwEB7lbXkhE1x8PZnQ1ysq4Br/fr+QCrDAN69ozB9xxhPS
BQ0i6dzzvIJubG6XXgEXWRT90TaaJLGWMZjbi2JZWA1K2RUyyCNjhAAt4h2M+P68
jkqEcN0A286OsvemwKbFOJmIG/VQhK9p8jFgSWctOoII5XTcO0DQKTberDWo1bzN
qElN9gmODswBGhhLAXqYiUvk2YeXINj6ivs+gakcUH8Vrv/rETwwCHMx65EI2fMS
GbUFfHibRdb7CEwPu1bePGiASaSBTD9NlsBgkUxXM8/7KIrIDM0aclcXRDbxnmcw
MdjTL1N5X9jDP9lj6KuHU2bmJBChAZKQKXFT77uHK1buWSmV8IDwRB5S9I1EChD6
W3D1uYjnGzlwz4eunin8KNydRgiHRgClXISGESbErK68RSY29Qa5HWeBBTvr+BjI
qBN/uJk3Ds2r5FBz7Xy/BRBpEjUh9neSbQGOh8n5/LjJq+BHzgtsQs3N1f7VnqJL
gXFZH7/WKZHygKRM/gXeRYJ/N1Kd14vhcB+EGZkTrqyluQ3rcy62Nct2iJmVT16C
MwRxoZSbDRZ4FKZBff+Agl2ds0MBXIliaIgOnWiRF5XTBG6auA87RACxjNUF2ULE
Hw0qEY4BdzqvmJFh0mFMPCI8K9kH7auhXaOAksXYHm0lMUrg8fA0FfFJqYLMqoBF
NfucsheiacfrdIdzMYohBHVe5PYsyunmSYHa3btBt/UIzMhIEgqulRX4yG+BxXhx
oqe9vacfUl7lKwxZNg743jZrCYl9b9AqMVj+uM7yPk0swU1aoxkNcYrpe+PpitlE
zZJDcPDv3huPztY3t2TmXuRUdQ00ctHC0vQRsz87Gke9TJL2pYP4B1YcLi9EFHwm
Nbkf8l4V1IL88gfobIy566HsxFMtk4C8fLY9GTIiWC67L1+vVFF1or+kyKt8BB45
vCFmua32gOKvp/7/cvIjdJC9QrvFDOBu6YusSNL8/FTK8cJmniP82+dHkZpC8qTg
sEKZqEn3qMKLu1yeEbC1rEa37OZgxdSAALJkHHURHDlu2i/9iyxl8axv01nU/dqz
0vh2xcqPFOW+2bMc3eBuo/BLHWEpJiownXkbo6ZN9PlS/GFyK3TOc2V1yT/pGobd
aaCS798+WW+mjV08W3fH3VwdGcli3IhHNKC2iVggKsT2paYQKdNjtw/8ZItL1Alu
H3S69kiETp9FdLQVf3NIjKeBGGJVvnSI6yarsb5q0puqCm6Pwm9OWMsgaXf2x6qr
g1g2G+4orDCtdA+QedEGF8r6QsMhbjBHIZZoLIkFb3esj1mvfKopflrjwwEQYDBi
Z/HhozFq3V82TBGK54dHxHq9QY12MYRJzaewxKi/mm+V2kV9dLe0AK2F837jfLpW
/ty4PtKF4xt+uK0vZ1PO4zC3KBf9Yq7x6DFOo0k8XMVMKjIydb2mI6OA5FVEGh6y
JLZOdoI145LCeR7VQu8fwQftjlCCpnHZmbN8815SAKuwzAMEgr13BysdSXbCEsAq
L13uveaADdsnCG0oegApWlJqsXFosJvwUW3a7ZGebuQLb9dKCgKy5qa+WpIWY90P
n4dtWqQAMIY6cZS72riElWZJ0Zzz5T9cQqJTm3fHfkDvU6znX+GOQKdgJAXATnPZ
AyswHp+AuiojQ+nRNG/9W0KvrX88i4nukOJcoYDL/jMqBpxDJTf1NHE2TAQ6lMAe
W4VtoWeeE9Swz8Ys4EU9qykq7bzSK7UnLarEv7/pEEYQMz6QEn2waT60BWlv4Ary
ZxAg+LRvSaDkUi4qmCg//xc+GGHGqI8XfxKV2D/grFkfuXtdcCp2+IHv3J4qqa8E
jbITAWcnsowNjpjWEdDEDATzIQrpc5P4OggJJBRBLyxgcmM7ebp+GpgDqXoJFXIq
5rc6XKJGfsBNMRiv7G8Fe3NP+Cthsve4CLu1Nye5VIyItdvU6AO4FNF9Wg6gObgR
fJPYKNgSGJeLl9cL91VCgXAbxcBcC7VD0L1rD/zIU7TZCIbDBLTy+RaYffqKO5CD
YGp1hD8VVewS9mE3XZfvki6Z22AqElc3yT3PxQLUiPM4C5kqcTP77dTboPuNQ4yw
cC8XNslapC9ilRKgFS/zDm+hyPZsjtJDqg0IFFOpv0US7he9zfXaYBrs8vOF7HyJ
MuVqpjlhJ1EOioR0SbFUHhgCUqTLN9ySnmaLtogDB6/+hUvcSFPR8SsEjNdiLzGG
DZhYlrgPTG9npFrDlvAtx0ck/UglwHg/BMOYI45O1zJYjCDsZ0rTaCkYscSoriw6
HzqMJDLgI0frXx29qGGRjETR/WWmYPXzLN7c+JIbnkBPDeRvK6rfb7Vt6wwM16lt
rBUBdTbYqkidnUPBjXYsgZjsj4Ro0zs38ohFUfMaB8sG4DdsCc5M0Frm8/CqxgyK
o/iQHZXo0zU1wTmfIsOMJ6/NIH6+gwfGKlSlA83IUXVdRL9OgkNb05eV955rKBIY
Z/6ipE91EfiRBeIRyADJ54XjtzsRRsK2S0izXNZOU9oPjAmJW7+8rAoVYvD8aBSH
/eW+6zgb2NrLn0ynlD0+unUQ3K9bmS9JM6BByfljA9HqX+PcJ+E7M86CWvadjIFo
oWp9wPe5y63hz2FmZRYjy50IOueKebmaOMs3fKi+tcUVxMZHT0lQJQyuvEVnLE2b
DMr080QhOq5H0qDPTu+CpNdP4coG6qJQzXIgi6Ccplziz9+ne5ZroOmYrzh5st/q
DcnvZ/7VOZttnhmUav+chQo96J7K5q/bBUW60oAfUrYtyMl6+u1hGzKQlPOJMAT9
EQLTXiyyDuDo8xIFHQY3rq09XWXCTCDZAtQ7hc110baMcBSx5ig9zqs2Cn9nln1R
4/OUF5jgt1nViZnA+Ks9n8OW5IOn4JSYHXEG1zdJ48tAM7rPPRH28H+4HBnoMobf
nPcmQ8AkI7ZPHxuTvkBojgDBYlapDGfKGuKUoKEHOdm7uf37YYhw5vwj9S2lzUVH
1lhfWg2Gr+Ejzu4NhHe51gAmGJFqhs68c7OPFeOeZFKz3JW2/uCI3Gi4XAYAQnrt
qQzlGo9OUWgX6dfKCUq9Q2tKJMm6dz18cL1tLxq+Cd5EgHA++Xl4PPDDc+h/3Czz
V2f3bcuk8HaqJqSbhbvLLZclpVBGtJMWcjqdW7crsUCVVNq7/RicGHIO3w6nChUm
2rysZaztXEjyJJn1V3dmi/+nCI03sUbXIAXxMC27rxSEGDrJIZEovb8HJrgOFn31
+v98B0aAp3jtb0ATEOcHIgsLJHnTOZz2ByOELbjtoVPi03TB3yekAXFOoFNmIcCS
zpIvt2lCtv1Bj3rxjgS+NjARbtEzo+0vSwYvCBASku7sfOXu2E+uaj1mGFv80jfm
FP6UJ7unNLWF4GPJ19uOUE8bV6wKAUa0HZ1n/3MIvaB2W8yfEYpkOIoOEaB5EIvz
hc1180e3JEG995Iotc/HPZvTDvDYomlPpWOvb57KE5bkmTG+0t73uqtEhBJdmIcA
BQKPEK1tTHpDnK0bX/9ws8D/qHnDvAa7rhaw423+3NLqbdWobzV2uHK9pBclaMd9
zPC2E6o5CQW8ABXHuiKEneGYCPlxngPdJ50rGVJlkLaDdOkVFnDzR+o/bVCoqt1N
vL7PeH4zdYPqJt/B19Ylwuif30msvH4miM//7oH7zKFGPvg85BHlzZ58aLIk2KRB
Wbt4jM1yiJGLzkVKVX3bmiXm6CbcjOo2KLfAKcck4c8T5VfR1BrusHcZBOF7iNmS
IlXzv+4UfMA8okY6oxUFGKLoc1v7OaSxk2Y2OPlki0nX8PfnND/agovd/0kMZchU
YL9mEXbv/XZ8WbN1jCmgkogrZyp4cU/WBE2T316naUwQoppGO1OB7W4Q3a8wsgaR
S4cN0gfPhXWoYhKgQfHRa2hoJIdhCOut2vb6pbvEuCpZjgtXiS1+yQ5X93IMtN8W
sZMyU64GmhWq7/ZIgbMUfn4FAGZX9ekKItJXt0h2R3nTXdpBbNIe8wGONDy0Wp+w
UqBFPcVkyb2uClbO+Bw/883QBX31+mjSsXN0mtGjig8S+6WsDaFBSB5y2cXTU3kE
RsEZJD39HQZxG9y6hefsX/0mKDln6SpemylMi5nFxjQbcIIA5X8Eqgar//jNPKzu
Cox9SNH6uBDeKYLPmWJcp4VvtWBT+NlhzcTybQkbOAUvTDOR4Oj6KwYlUFByHdoI
R7q0SHCjKkeQwcVYSZkVVAm4Tkt7titx3wj7s2m1Ex5J9O74KgMvzDcwb5LKvzCe
uulzLNHhLL3JjpkEZl3Buxhqui6EEjkJGSinYAyo0tuLX7MEBzvXRTUZinp9/Zlv
ugPjHvj5Tu18ROvf0pcGtOojAvXDtJJLg4Rg4eX2JkYw98+ReqGEGDpp4ZDP0vzC
4DFkEBDG1dLWElHBxQWI2fi1SKgCV0HG6lZCNoTMXfETzJTN83yBrACELhC65lcQ
9yxhG/H6MMvT3YDM+5f/0f3qpTWP+SWLW2nWRon9de8kyb6mReTHmBrDhraMs4qJ
mnoOC//j95U/RPZZ1/27/kLqSiRr8gw14cDCIFKnDI2J8Gsc9NsnveSGLK4kA7WK
h3FT7Eq+xw3RgwouwEbubI60lvg4LRO3q7Q2yzrXkgXuPQQLq8kEQmV5BWjDI1Hp
vJrWEsNlYyHe+zdt+YWrnFngZFLXqxb86eFyLT8Kc2e+9+5PFqQQNvDCsRJENSA4
P17B/8OtNoGyrI8xZtNNTMi9aBb1Bof89qpIHW7mCdzdmb2R54uCid+OT7g67guh
PsYA2KVDkRz4PurkLOafxVr3iJr8rlELOjfm+hEwSFl+b7Ozicd1DvnJi1sNJ3nq
c7eZmrE1S+eTDnizAyTQOtjI4JYc5EbTjeSSkKSz05JIzMAxou8dpXHgUzy/qRi8
tIpiamDFWJIJayGtEuE4gZFNU+/dYvxl5HeSIqLNYDs/CsU8433/ZO3RYK+jO2pQ
MqoZX5Feij0K/d19YtMFA6QumIak3yv352pOFkk3MqI/5i4Ddrj27eZVaaF3+ubw
5DBlZljvDZYp8kTBeXrorX81Yp8u82wVjDX6NVzHE0CS4QPeDEfcr7UJu+c8xpHu
YRGxGDZxHqmb03ABk6jhWWhTKZ2a9q+eJj4pZqie204NNUdFuT4o6ITd+QxaJyGo
+OwNzdU8WPPaA1rMlnndT+0i7Ckzz+AeLUVtywI48jPzGdPaX/pjNWlIstfVb3CO
RcNwm4QN1axLoJuYUTd2UdqzhmcPnGey5htiPwcm5wiwsrbmlkHnXL6yFiEH3AHJ
Wuoqo+88i2qAgVOeVLYyhvBnNVm65Pkrsi9aO9koZJKSqLdNaYt66O6Xt73FOYgp
4xH9e2pHuaqQ6ume4iJ8YBEJp4s8WO69HVXHugE/qJns1EKxRJ3OhfmWxMPNCNnl
rJBh4flPMsfkUo19+DWsFCjlhEKGNUX4m1/U8l5N0poxLOg6fClMefD+06Jn3qVQ
9EVv8SyeMYk0/pzAeH1t7sMXSYCgP02BByK/P812ifQbTz3ctukooxCQ/wSJH3sw
K4nob/jsgS9C6+bTPTX2vK8url2XNIhp0C3c4MfD/ksmxumyOBd0mDkcA05UgRBx
RLwFvrBQKCiyFTCx+VpbGZ3e2L6Zv9JnkKt/yvw4ZzQCyeu/1m75IgfQ9DoN/VrK
yEGuZJM4R06Zvw7lDYpZHy71dMoGe+dbMfHWRGNVVDXqjn5iaN0ceM254VXxVGYK
tBvlfxukWduYdjogsSaSbjnBUzwg2qIFpvWzpL/BUwhdc2WKl96Djb+9Am59dsOf
gFKsiDulRWc+GGrTQQsBP+m0khNoTZJNhAhBNXdmPgTA50bRfmTPGhm4VjN1oeV4
VYNMOdL56e4s3GA6/j7mLtb2pM4ywvP2Tyk7YyuGLQ6VwuB20ri8mJAIIEVQzHnX
ZbJf1wYuJPC9VeE0mJ/ql/PVRVV5PsUrwbQeqgMdLv5V4hBRu6bAJ/meNYr8CgcS
Qx96knR4vc04kf+FSKzwAU+nCW+1cEav0t2nFIVPijqbrxmMKDOtUM4BX+T2Jk6t
9yj9VKjerCTRdQeBWddM+NLOXg2nWPKStrr5A22ijqClNRtdJKU/RjVlJLOVx5gl
0p7oBzOpmzKF8+ThGcVBSwC9kgLIidd7Q+BvcjByofuBb0T78I7IDu6b5ncaodNn
Nh4fal8VEYrIUVUp8JS6OPMiDk69+KmBZHNTkBr5xhfsPx2WN/5u0s70LpHRd9X8
rrknykMMmvvbn9dVUwroHdWFULFeIH32y0SYFNhdc50yJZu1eAOZWQqKWhnpIy2O
TswMrUSRB0dRfBD0b160ri/oom8aBZzJcAlzYRnE6DqCuu0JOUgV5eJakCJHGNhA
lrQ2rxyWSzC0q3XXUHGVBBFKpnWw35QwaOFo39yQAxdEeAdAymCNg3kjZfTBoBwd
Uj+d2+NEn9t4IGYHnngQIYkvlozGCel94BTEWCiK+1f9Vwy3pOuMB7vvO+fTIRjp
17SIVmkUtvuBQg+wbdfVtv3CcsT1FCvEsBViiWHBWm7y8HmwWNiGut9zbz/5kCXR
WrZfj9IeCcTrVLsrigGwwcDwlzFlwLhLcuG3njUdfhN2j5ZCwUG18OmAHvBzmWfX
Otzve9Otzj3ZbqGgne9rb0+JrHKQCvxz0Z9TIKncts7GhL6Lwir9WwXAMvwWLcHm
5F0bPp/x7Ajfzt93HFZHbEH4LkCNLYwa9Wh3Q4t3hJO68hia4FC08TSDKuYK8NOk
ywVu82fZCX51v1JlEG9BVydwKrVsPI4K6znRD/Xjcpjlvomtomo43+X0GYYhrBEt
8Vw67aQA2p6+/l7qC3yfDB6JldWbkv0x1TkQTIdEO4cQCPuhftBkJgmBDaCKDH9+
efAd1aNjFqlulmdNAx4Jauz3bsy6OXQhmjg68zY/wmeJZ5hijNwubpplFso32Jw5
HW/RIZHGfFMuoM4Y+uObSBFZKvBH5C7JjvfEdlEPtKhrDoLVcTtt3H/nTCg6gHiN
FbTTBQuseXsNzF+nMbg3d2PzCsZ4jrIagZTGUQx7iiObqD3CdgZ2qj4oZVW62+hn
uzlzPWqivafNzlfOFh+EhAZI4K6xYa7j9jj6UGi+JnYmpwHEXikPaRWPE9DnqUDa
eHf/aeYwKBSP8Ayxzr9xdCgBTcfhOsQHc5Ic+UsziuSCAm/t/9+aAhoQQLs8TPXz
GoTZar8yy4F3X4GoUWPSmQv+IpWfsdQssu6H7ChHZXuZh73GdHcrtZYf8mblYPDM
f/F9XnIz8LJRn55eiU/28lrkbXNbR2bFRe2huNMzz2b4Oc0HWMAg3/KJDOl6cfmF
UTM5E/tOUe/lDZE2wIyt4Fmq16E0v0aZ91x4ey7tCCytPmNz5yI41q3/foQI7b96
y28uUxFb6nSWE+NsFZ41UvDrRhxCIETz2ZE3gHf+ZecrBc//rp37f/jb565npUeg
e5KOTadzhCSmA/THNaMIpqysK54vll6L8+20ZlhIGAPyCdzqedW4MXygNX1gpIGS
DpwFW3uMKj9dYhVLaUXCrvcwSJVK7wHaenJV+VtrWDQ3RjoR7m0yyNkYDTft1r8J
tyDBgTYDomUYf29iE1Q82xEfQQSkHAmbdHqJn7f85/NTE5eHyiDjoIyNikjpXxCY
y5mrmVp40Sdccnsjy0ZcsmwR6fhjffLgp4kGynuprEmKfYTdYCguibVgMD3gevcz
yyNZyHunHgcwT/caVxpZgGd8POPVaBze40/VnpBGdlykdKan+g3G3WQqSOSy9fQN
RT9vebBKc69aXVSVTpOxiA/M+8tAeJ5mVp32bWY+HEc6AhMnz6Ac8xwLfgUv1IWm
Yg7U98Dxh6gX2ouPdG8r8BhDXfc36EZ7JQOb1yUr/YSEAD4Ejeb6mnHSKW2+kABY
p1rrEjZUVqBGCrWaGoQGlRsOeGg6RA46g1rQe8bYNkkkgDPrKMVlEldWWPMHL+42
MsIOWPOjsk/bGX+4Wyl7tV6RzL+1dx8kUl++Ddi0OoG1qP8G5ZggAeQflIcGOkj2
7hFWYaE8/FLSdDw+qA4fozqheSmiw9knrX4d0I4tE5WhrJtqzj6jRHezv89sOV/g
key3U/q0xCGOBpIWgW6yrJLy5yU2HSkMIkGBY3KP3qb2GsRhuFoq5sLtrrRtRLBn
TRt24+Xa4dUKY6azbKYpLqEZN1Un+qnikpGnLbfF9RHPamxL/0BOk4sCLommcrWF
cHpp5hxGJWaUt3ZbVaw1fStIGyROF7R3I8O5YAYZkifgs5cWQzMUX/FK1+TWisGh
ohGIeg+r3t+AGZhA0WpUumAV+2JCotPZ6Mkij4trwQmQKgf/OHTXHXTQgxMPDwZ5
5urVzYPZdSQpIuZsJCBI148APDMMG4vENjxdA7S8KFwEJcybZvaWbj4fGDMXQxWW
9fHnNBoffnSBTXV3Eqmv+90XOJbfL4T2VyQC4ukRba9Ey5pprvNFfTqguaCmv1KR
6sA7sJNYEnQLznRPqc4d47FRiwIwZfpYcSi5i8YLv/bIHc61xM+yasFa0IPJ6lZs
P6TViO8ldjTiP8paH+RDfAKpbzlkGEMGZZvcoj/AHeo5GyMqRm/kcK1VgNkvxQgw
OzZxvEo6ix5RsV96zTUX/Y1RpzPp5rqwmzew3VCdIfCqeSDaofyfH3IWvLoYzC4G
A0UgThfF816yfuZc6QObD3CUZt7HojiG3yufYKgeki+ayb+SxCrB3g7ZR67u1Bg1
t3rF4utkU81u9qvgfyiPUtktkjMiKUzqKDYclo8vb496JcqHjhNsNgIouQL4M2IJ
`protect end_protected