`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
zZSxD+gXg/oJR5jdsH5AQ98lZJJ9TPBKB/KkGLtRI9hq2BSj1kjTV3z8bGrzm86Y
PirbhPPTGoZkTKLVZJ7bPDi5T/QB5Az1wuH8FWh4OXDgT52z91kIJVwtA5ldN9tQ
/rZ/7LGzyhR2MhqC7jAPakFJkULTSwxQG2pgpH7wAS+m9hmB6sQvQRTXmpDf3zVp
DbdKZ1V9FY4VVjssS1QNQyp8tW4S5BQ0X/kmL97XRAiNrXpEtq9V0FpBtmGhFfPy
oOpct05oodDLSFLbLMl+Lh4SJQn9/iqWo34nE/MhEOFKcYCzm2ZNGWXn2Bp59OUc
EOQqiKLh0dqKGwgihMtyy+fnHULwsX7GQnHZoFg2FFetIYdnaluQ02tQAO/6Of+J
Jht3kaOHfvCh+YQe0+7tCVxxPA731I3KZh+KARIYIfA+R4NzKVTWDkliLfPIRiW9
JF2gSotjVaI52bnJCUGSDqJClbOEpCCBmscq4GBsiYbl3Mr92ydOzp5MIsX4uYxQ
wgpsCQ6HZMtGH/QyfG+mKi/b2T9Zv2a1hjHDcENkjk/F5dTJqls33Savj3xy8hmE
V5gTBra4wXb3bx+KLlIb2+5XPebV4ENV4oQivbFE/w76H4yV9R/MKQkEyPJmvfFm
7hhoMtyMYMDUSA5UYCKShZRAoxN807haEAUiQAzpBX6ePFk4ZYJnJkLJgr5MPwOd
Sp7gR2JsiXGjT+kGpy4hX2OWVzTiQ0V5LSuzX5D/p5yXJisQMBlzApkYldkQLOYa
3uHGj6U/1ez8xYBu3EOSdEjguRQjpVM/zkVWeZvBqzozHnj6+Gb+9kUtqm+gDiLZ
RakPCvCGbnBPIGB3mrcusFJnrz/IfE9+4Qb1MkBQ2Fy4IaqgBRIQPD+1+0q/rD3x
lI/q852f97r58rePfGyNUjGIUelO/6WrDQm9oGDk3l2GxG0lVSs2XSq3zaIbbvPL
2K5CZ9l+kzw8YBELYCLl8LNpAZ7z2wUKUF8TrqYdWZqI0d5NcXZQZz0n4ThghSw5
PadwBfkzEziM7l8DiXAdxnFP7lTu77SazvmTAAnUmLkCa1lgpzicQrnKeIK2GdrE
hW2+R5MenURrOCQKe7mchVnN/3PHuEiamjv3u2rzHy7c+Sc5cmrB33qUgAMGNMRQ
dngoPN+NpJ5HkDpt2Wv60/qo+WkLAW0n9z7WqSTwaZM+HH/ZKxEU3lu1nOWEObum
jxnrRPs6pPkLtp77uFA3WqPkPWhvuR/PzXhN65Np3WpDM+xk5iZC5uuBfvgAGPLU
BpMa0mJEmnvapUP/QAmBqeRY8It1MQRtQG0VgjrweGKgV7Iews01XQlTTzA9BSCt
0WIViK2QfmwzBpnVxli0Llx/jlJcRcxRxmDopvTgkplBHzjAisExMFbb4MQWkPti
lRc3Z6KuGhJ4cfu3x/Kp1hIPmbqAOZ0Rsy5hdPMAZPgt+Il/LRlvWFnrsh9vrPmC
qU6Zw56CnJeRyVdIklOwIBj4WwYSQiss/H5nnQX2bBrq8+GsAQgHpCXlpFrCDjjE
P4X1knTyNDudl8FfrHGFrq4ey/y9UmLoBjKvk0PPXb2sfnlI0mzPdFlhwTtJ9ZoF
Q47lnOtifBWqVI1+fDGCOD8cpeenIbzGFEHB+ry16kU1O6eMgMiIixeg6hG/yFzZ
wv+ZPDzbTvykUdXS+WeckLNl6QunpwIw2Ys2QR58XpGFCKgBhK8Q/hCACPcUxEc+
p8uaCC7mVG0IjFupwBBIPapuPCYFg4XicT0dBpgagbwLsp39s8yaryNoh5PCO3MY
E91aNXEW1SXAQni8Ws/fNe5M8P82FSqm1+k/pCyiQ1l/MkGfRQt4bxzbYNm24o/p
JcW/sDUdqXiFSNegRgjJIT8rjWTPSvO7tso2SL6p2R9CytN/M+4daeVnYPegIZua
9ZaY94ljH+in3HhzqbuVpfCO4w6n6fq5f2WMyYaWbiAHmfuAUEwAgU3W5xvMd1Wb
qLbzfrw9Tcx0OD7wm3tEhHl4ZL1n3mndtM905hVNai6CG4p4mEIbK8cPOKv7RlQr
NhUlpfctsuQudobBbpr+IzxohcJ/QPXky1SagJOQWa/TZsdJf/O4GiSYqiVwEVsv
vxoZei1gEFMt7evPDtlxZnZ7BCw7ibiksUVkDO1BakuwUVsWu9WRo2fiIgmqw4Rg
ZQ3d8uURzWRNnPkrEiS0WOSsG5GAQkpO8OWHufVOb0NJMMLQ8ad1q/kgpfxwW76E
x3fd0HBCkUFwEGJ2o3feqFamzvKHl8MJYlo3glj3hqRI3+R9RHEKAMazfmtJsmAE
x5iYtsiqVuyY9punh+ntawG3mxDVs9fGyYAtMQdLkcr9rJraL6MM8bqI3UgWyCQb
wADRLTUKM3h9v+Um98leq5LKokkwZXST2ycAvMyFNTy1UW39My4XyId1wtOEnnUf
/LXtXXnuow7cCiIwShE5K6ht5B3E9mNTQj2OYe/yP5morayjLvL5ucnfCkIuYHvo
3bem3outIXtcNl7mvhi4Ug5R0imNtETf4mrnvSQjcojozusouuoPwXZixVa/wts8
/6wBY9zQ+5NLkmOAo7WOw9dJNuZUOhSrE7sdzwM0iu5PKuV46CbAKmBxLSump2Bp
H852PI2kH13L++jEDYPARip3T7lKwkOwV+tXInF36Ij3LJBiAgvDTcwFyfeAkz2s
2MN1LhukCmMIdHE+l9CrrIF1f6qbDrcvPiTetx6R6Y0k/EyAJRrrthkBxZiZtRLi
lDSJjW+gJUIxeTkE17kO7Pl+ZM8oTM8LHSV0KZ1svgAcbG0VGve5ReKWl+M5PCgo
WYeFRATEask4hnF8nmD+NAO9oviY1qPv62SV4w5pD/CrPzPi8bMA+hVwlIrRZ/O7
HUBa02p7pjpafMpCcuwcDvdHvyjSYZ1z+hx05G6vzk6GGw8nTMEPVZKwFFbYozIK
FNBETQghM+yitp4ceQJBQ8DNQFnZ1xJbckTX3rfwZKZIT/xjn23Zfgjjm7cprRc8
qO2AkGLDg+3QRIXNl6sroTLfEe1rUTnSBvG03YlnyKpkWzsq+lDRMEoeUI5jinaJ
gVLzcifu5wo7a4tLtyIRRfh2F4i89Tru2bALSJ+nnCITo7KbdYN7FcC82JE18poA
xAwj1qzgEFFD+LfYEPltbc7Yn6XcfdLNkKrt7/fDp9Z4jXxx5XJJqIbCdU78+JKf
Ikp/lwJ7oR2GghSPoPWPolV++WdJ4zwjsEs3f4wiC1zzcEyfyiR2Eb/HXCvn2Xpy
PTNEej/oNXYp0lT+iCbf/6OasiJjXU5Ua6oLytiqwqjMkZnz39XwsMJzafIkKbbb
u9Kq1C1yhfQ0a2qYg4AJ8PfT/F6OIGzOnO0sfKd3vXZIg+aNA23adtMQJpYp1z+p
pShTeMwUMrqjpvc6xM9dUoOWGAq6JT8qOrhMDYKVNfG+oEpWv2N1+TY4Ka1MzcIU
C7KgeTWli8SvPbUkMI6tsFHhbjTsDVJHUzrdz7+IskH7XyKmF54Vx861T4gj4mmf
JCl6v8CWi3g8oI8GdzXmn8TyJvF3F8QDMXl5EoLQ2pmq1teSjdcq7onSGAWeSage
fyEbZOfwj9eWGuHs9yPXns9QACuhmBMGiXuD2lUQNvWi8TqU5Ie/Y9CVVIsuxNaX
r1CueZ1fGDMjHSaZjbEVwotAAiBXA+PLj3MHsqLrRjyyq8mZ8euuDFbDHgroRlTq
FiWoS2HeCGLoas5nLYXK8nrIx8FosbivRUrKhjV98s/L5kq2wtrx0PXW8Cj/e27O
IX/hRzhAPqahizKw2rxu7ywqiUj0Pk5tl380bRbQ8LnNXy5QrH2unFUxH2RR43uX
oGwfISAGbeJGbcChZDfnhpCUAd9YvexjBW1Im2sQBSBSEy01cidCkhLYlKvJjgwY
kI4tf91pw8BgP1Diell4WehfH79kdJNWrzEk3/wlQ2nXZdm1IVKuVcydhk0Ctj1D
SVB5tvVVhWLqqpIPv19gGtiseCRVda4p2bnBAMqsnVrPh035BEFnpJFHqq7cNaXD
xV3d9308PK0ZOEsAS+IuPs7NPIGac2eAVKc1JJOBuiISdqjDBX3CS/ElTc10HxW7
JKjmgjaXBrKJqtt3b+4C4eCV+PDN0VeTtXM35m0hinRDGqn01eOly+xFyxpPc8L7
S2tCSHHpieIDP+HuO4K8yMU8sYbLSSfWGv8xTCVRfLYzWIdY/jr3HJjfjPmsftHL
EnPvyX0I7g19QGRmigy76NwqtQ6IOr6G60ENJhlH23hOHOFcGrrU2VL2YKddI82i
V3Tj3oXqGeoXBEKk9WonHt6pKSYywwnfZZgiK3I2YVT6Uge8pnZAU/DNqRAcP5mz
ODwd8v11v3J4zcoDX00DRYh0GvHPPodVRdxhuIZAj9K+FD8Y901+BMP/754y3xwu
lqj84YAdTjsUOZxFqz4eht5UIAnflDj1cxY8mOdKyiTkyOVzSZJsnCEWUfMFgwRZ
DYXFcDTAyxczyx8W+JwAcUS+2bl50Uk0q+xQNkr0O2c4nMj2cgQ7iJ9hcVZ25W68
Z2he0PF/eGC/gBudlj+Y7Lix7rZTUf0DepYK5V37IX5hpiNjBTtmy0qdhcPQPjII
NHaqZ7hcqt2f9tWAeR4vR56g2InKb1SR1PpoRRKHYMmdvb/2+P6bSnJ8l86akf3u
IwMMMS6jFSvaAgrUrJKTzQTSqM/SEsoO3GKLaBEzV3B9CasLwuRpojsQJE1SksZt
jVf7ACeWh6efW6XJ59u1G/TMNi83UB5sehJEhkYfPw8YASzXStykkBtOrHRKtCdL
3xEx99ApwGg1NzG+MRjF4KZHRG83g3/xWxqIZ3lTDrJr7AsEgR2OE0sSjWuXLs91
FiMifwjUX8i2VOn14ftv7kmd5/L+DIUG9J8miLAJ2R5hPjSDIOCtN1cIFyZRzQY6
+PEXmzeKzEqbf5HQ9iTXseWs+Rubx9jw6+LefkPg9bSXV7jrZsW+FV8hwPGVQJqw
THM7b9Eb988Y5IbvyqGVrlGseIxm2p+PPPt86/WHiLBlJ4hxAcaqfdTOiXQoJ2Q9
BNCwRLmZarvgMADA0X8RQGNweE/MjmGPNWMbv41eOvGcFKb6+Is55UKeHJEK4c+z
ptN4E0O//aK9vOjt4oVuceGN8ZHbxog3phMmoi47xq1HTsGEmiP8O+dDiiRaQfYv
YBYapKYgLIg16mSGzJusPg1eawS1zmNc8XBrd+u4NLgAUm7Rhkqaqxllfe3ewM3v
3bjcgtCN2x+/TCcLmHbTNCOovBygrHR7pxUINn4yVTr0uG8WQFkdDEb5NIeppJ5p
vW9q8FM0n+qwsIKKa0AzyFKwrKLAM3tarGPPfMkuSlFep9OBcQ0ULCJ55KJ6xEdu
Uaa9V89dmrrjVHRN3pHU1BA2/GniwdPPr8+VmaVsPye5fk2yzkKfA/mKlLNW+IL1
7IKd3KpNKlEp4BxyrTXYwoK3Eo8mZpb48XKjoawKvsabYZ9FyKng/gQKv2K3MKBz
kIjrgAkYBs+wxuU4Oz8rE7QqF920on74otDVqPrP4oCJ6l10Sg3lLMj5nVNO9EFt
sv5mFjjBeoi84EcJ+y0NmCo7M3f0ehl0N5oMSgbD9YKjXrDBUCQEsOuUQwYV9ML5
vncXnYyPszGU5WTsIl4s0iUbq+N04K8FQbhuf7Xio87jIz5Y9pQE8hTMM65ocPHK
hqQgRzd59VNqPd0qAe4sxT6/X43bZNTSoPMupLq966u1CX055nhvhxG05xuxlUBy
lQ8LpgEEEdJo/aPj12/809MG3JZvTFV+6t18Lnyl9XeJUlmVF4AYQ0d+OFZ5zMV2
uhQBSuGuxpbJDkoUEt092aJB5+mcsKM6qrFQfaPdoA8EX1BO9QfhrSJk+Rj1XJPJ
TWsgXIQvlamLzpXoAZxzdGeV7HqiUpd3zEuiSynaGV4tOSq+gT29cHYjsKf4higd
0RiwIndeVYYevpxCNE2wKKaC3BroON11jPpvy5do/mt+m76wFp+wmiqHY6Oi736j
J/qfc8hi9zf3ThTzfS0JrdB/DH8o8OzKbtBPUjuy2aT9Ia8i4bGk9LwVZXYABKkA
Ua+zaecBk0++wJlMwQByoUq79+xrmEtNEblSMGJpYy8AbnE9UdLHtZ6EBk2U0waE
8nbEvxJdg5my5Cj7q0+/Lqx5SauYXPvujdnlajcM/mxWcUmIaikvlgSbA2XDO0oq
7OBLek2smFHcV25PpfXTcOY0y0ymyX30giXPdBv1vHSEEj7IuF/1opktudG1SJ6I
WNY1OSaRMSzr7Gmt3LsV9vGne5O9xhy7m9hUwYMj6tQIEtWfGjHTTltnyYCcXvsV
2xsxBnUPaSNr/fxhqO/HYRxPXJjEthxgBg+l9SOlEKE/pRIKPO8hMLhKAB4K2OJG
eqMfnuV9MYP9v0fDtbUhWsQ/XkhdW5XWCZSAGmW6I4RBH1XTdfJAbYDngBKCEP1E
XB2lXaFBriqekwTxePJUXBRzKQ4TjVS/GdrzgP3VoNFuUOttRxXP1m+Bn07Syge4
vr7w3+iGYu1UHoa9DoKwtSCqfcICb++UAwXKyqOx9loPNzt2qGyx4QdGvN57xOwm
B4oBoGYB/X9Db78BLV3X6k9YVWVN0kGK6LRswMdxkQ+0HwYiRaPoqIbUwOUDk3tL
5Pc0DYO8AOCrdhESAMayczuVOj+Ib9/8/5UptEgKNU8achP/8kEnvj1PQsltrDLK
p6VayZWn8CTp4tvLLXfVGbF6IztrLEQ/VlwSF388TFXed+tsL2ksyQixv1gUldGC
OaH7t1m8gRwZOq9Z/hhTwm7VB9h+sjgJEztoFF9aegfS3zawcDlE76/xUtXB0DTf
caAK1h4yJh1Hvwe10x/Z37b8zJNH/AoBuhUFmUYNy/CIuffLWquipBVO+fubdlDU
riVPnwhvGVCuXLVRJFgTrHADiJqayCrPC0pbYqAA9BAKU6AkZDF+NpO2ZfocCqjP
DXxCzCmACS1Rlba9l7ppyEQ1ntPsKW+N1crH81wfXP8oS14tRP09czOYbf0FOQMD
dgM3YP4DM7Ts5Q5JVFy2pr/VSNEvyBZGPvD5pMRu+19cjnXiedIx+vZE1ZAPQkSc
Fr2qzVu/clHi69RHJy17rsrTxAgoixvUkYkR3VXJoQun8BfmxtU78M/0VvDwiZfL
K6Eq0JeFroCEoiIelCR3Z3m5cgucZI6wmGWutWwwAgs3JtIh8hBNqabPoYVhnEQj
SMxTO1T+/tAivCe1RGINWI7O8gNuRQYAvPX3UH7GDSA2xl55UFyu7ZBFW7pFCQdI
JJliOXexpCBhsB/3mvjswx0CxOoQpS9z1vcIBZwPctSDngjZkbJ1iAZ2/r3ZTC/N
+xClev/RXUyrK5MTtOepphjKgxltbltnwdSrgREoIWopCA/2mex4caw3+qhUkOAA
ABIII071GfCob/NANS9gu0mOOyMnlYuulpl0ykHgvBunQLPE/yfandPLzL+QdqaL
MzkvlnYg/dWYc6ATniC18WswoWV6VtcTlbRahWpKRquX6LXhfyQOmmetnK4xtLq6
/PTlBRpWTaTRpWGoaPsoyC1NXmS7Z4jVhhF9cPae+IYgUl/dO6E8MtlkcooCYH/G
qPv+NfILM4oZtcCBfZKly/zkDVH7r3GaccW6j3CMyjCE8IkhW/IOCqbyX+wNbIqr
4/obI6G/owYYu88X5RVvzeEnJZZYkL9hNSD/RLzgVDZ/1zFz2moaLEDvfWvdn7EJ
vyG2jumT06h7NojZiVT9KgxR32OBXMgI3bxuXvydvvpzGSd5VU5qGAbs2iGojofU
RcyMvJzw1y3cd9bq/Iza/U86UIwMSguJ8dRi9ed8PlhGjrGljSyTA4vJpd7Wvd9f
qW8WX6qPIu918S58ILBNm4/pjnXZgbyoI4Sp7FeePUuK8Tf80tv1CXkZQjQLMUCR
d/IcwLyu8nsak4fd/x4dFuS1K26KQWNkrLaF1pT/aWHJmhcySMl10vr5rVR0HVs+
yDlwYrSmZfoweYuIH8BvSvzB6AJB3drNdjh5DKrDJ8dnG9jvkleioQSbneTTKy0p
PYrErslncvIaQKBH0wJ1IO+qBmNMVmPWm8y5Ak3canDhetUk5rbR02/CrVB12NL3
jaWjTT+CAoA/s0RBCrijTKaUTpCO0itSex+YJme3SfMDDI8avd7iqN+QEQYxoVbF
69COSD3iW+eeqE0VgLHGoLigrOSI/79KoMUmh7L2pR1W4LRLuJgnwJpoSyPJaDeB
e5TGTcBPll+WqT8/1N/JYujx7BSOuqfFe3FtBSZc09uqsxnxES/krF68JDG/qezr
AgcZqClsYX1ryUlEggyCTV3j/KmFjm9qiiJSd89ER/qnHYJya5UCLTgnjS8X+u+S
4bILoZkCc5mUFcVkKRqfRkN/YN4NtQTx8eRD104dVm9JL0scv2dzkHjYGHGT8uwW
MKr6nj9QAGiT1qMyASrNVBq+4DV3bRODlH9jCX/oQ4g8Anjf/wg1yZtaubhhcgdG
ZlFsuOwK3WVV2jyzlKKQfTOxtgLZM4U6Q25ja4YzurJypkh9gFoNEWGS5PgmCELZ
KCtdZQM4BCEmKZ9bauJTHcUtg5+kjsKHPlb6yfELKJPa5Yu5Iq2DPsg3CEcsKKa+
qVI3Ygx9GtRWtar6nGRt+EaKYvcgvAji8dyKELkHtiFnpw4x4t7iJ0gIUEsZq6zx
mxw5h6361Jq5zPDyeL3hxlXVqx1kGnEl5vRXHTqGok6d66A0RH9k6oNWeOVq6Li3
zqbRTE4pQCH/cXg/6PI59km35JJOFFbWQwKUWq5su3qTJXfcOphDBdTyoxIQafx5
NetQQvfiThZafZ7gVEqkm8BEr6rwa+w1s4HYTBH5BQSRP/dd9fMdqPgFb3zYTyon
rMSPUVX1POyz92JAf2Wi/f4oUzNsKCucTCV0RquMTekxJTyEPYR6zWj+cIGFmOGN
i5k635U0PVguKRpRadlIHmf5ZJ37p+cEc6KD/rIvV/BT5LnPbPLMH6De2283y5yM
a+pV7aBP5UWlSmr+xRDMT8x2kVKg1/QvngIJC8qCWqhq/gw7XCFOGLw4DGfAbSkW
h/zSBsfRxA/g9nax7mwkUzrbPvtiyq7Wgz5T2uhfqSbKteKgk7/DhTG/xpCJr7JY
r3cNOSJI3F7I/SDoeJ8qWdjWp5voU3VKQCKtLrEUYrg63X/4P1xkh3H4PhcYxH4y
BjGBqbbr2rEBAelyGsHlEPqsrbFMgYCBxtqN3asNNrYqLKnNcMQha04i+MjQgPjt
+0Z5RMG/85YFgpHa4Mt4psmU+0bEhSgl97RFpPgyVW04oYORyHaUQBN/LYU3Z+VR
cKRtVVzqknp9qSU6sRBMNE9YMKCx8CnroRstgsHaLQ9GLhz9pR+W7ULXVd7zf1cn
pVfwJApgDXGas1NUnXiP/ys03mL9PYx7+Ivi5Ws/ACEfI/JI5L2j/n+fnjerpDUA
d4/jtJwEUdC0tcz9SKuBeK4AChcGzoQyqHrN6+l3YR5LsYtZMDfdzPgrdsZOv6eU
lfG040T8kUser/1v0sCmXbpPZRHRvqBdsCi2yLFtdmv1jG23CpBN9PFMcauqIUh4
SeGgW9uZxAqkCO/vmvVTOfVkDukYqCglbWWR2DcW05cxBmfBMGvNQkKCz4GI11li
oL2+xBIREwCeSjUDApkFY5iPiuPjIZZ/P+jORTgv7J8LEXHVs+oO7agPsxgI1mkn
NDU4wak0XTpxbk1xPVrCkysp2lbEnIqWIox9NfJFjZCdBjckY6sj+MvSMsNq4KdF
CaG59Vpo9O/xcEKKiefXJ2+BlWLwypZTpy0HP1t8WJHmrFQd6c+Rc3jAUIJKOccT
M3ZwVZ3nIHPX5xiA3yBX29dxH5j7xiwv5JzOF0NLeoGrgGHWzNJht0hlZ+C0FWtj
EqDi5V0KXz535qnKU7Pu/r2qtw5hX/lRt/1R/2bGEO2hQYH/gZDS7myWGomZEfZC
SAESGxT+5XHxckpjF4jur5Y6ehpVOhhKMmWols7I+TTAaFeQPPBcKppon8wLeQcC
dxmld13ac5E45lm1ND0T1O5RTQvRviNh5qYGFKzcsA1hJcvVi7apfUZH61FVPQkA
JXD913X5SRLlOfazx2OjemP/s5zNSnNlI4Mo9QDduKsrgVUMeZcwtFE2Z/QUd//j
PEXTRZbbNJCOQfEPgCnDVEHZ2jUKiDwGwDpnnybnRFcaUaSDaGwr+qnxx9jO1RlS
bahlmElm1KELrPlKCsfm309VKVwPhgTxpr826Yip0FCCehaojjuRXu9OxutqZhrU
lDfvUo4xA8RfH+LfQmUb+IEwIAGR4kkMARBE9FtzYVXOG/O+Bqx2ucmyzgZ/P0bd
ARVAjnmMTvEDmXN3rVClf8QMdP6qqZjKxD6bpqW1BR5gzGVbPtDH8umvNwqY+Oqd
nK443T6NATh9UYUUsJiHJN+FviLhMbmSlsus5ZJOggW+ujoKN8ZNklMY+catCyby
ABZ+fCTpW7NPxG1yrBruo9A2rf5yTYUobXkYLxex+lsyLBAYUaTBQPWVSt+g2lux
hrFHDEmrrD2ibDQ0FqKZo3qJaHNqnW5xf1wX7YrYHaee68NSJVmDh7ie0AyHlnLD
t/k/UcOnUEQgyaRenEi8FTfUf7MiRfFnJo8mYusvoJW+egBezDRXJgndyCDerTLZ
Ao+EJ+J/LYF8lTTUDON4iKqpJvPAUjnPsP+cc9LRomMMGjQWbVkDtswlJBlzOW0j
aA08q9MRwDtT82JTn74GT2H4/7sfexT+3NAJ0QM6MnQQXnxd3+92YMN7oEJJr2Gf
WdHoNnJg327hIY62VWjinRNkrh60jm4V11G8rnQn0ajI0TiIJgksvIaf3LCkuVQC
Hh2k2L1AwTQOg5OtYrqcaITPKC95NbFJDTIXhJ9VCjLgM84sK+w6qDEjf2+OvRIm
Q/ue/J1mplWEFzT8njAGztokGeMtVOaJFuaf1zja3U929Al/zOmI09az81ibikHW
s3zI/1bqnkkdHyfst1DDzuOhW/iXGc++8veAf08Tr9WfT8nMs6g0ooZqGoLcnl2m
7sMxg7rU6D/uF7DT8QAKiLSEBfDG2varZtuCzm/MMq3eLGy6vqpP2C42udv13JWv
XXKFtMBFT6JETLZKene5BxVXI8mjXGQGuQ1EJpkV7Ei9UVNMuUP0Su3dN1Xwf0F/
3fTEhb8BqYJw6EIR72HJKNAuKXh0gSdIk7Vn16rYTS8Ty2Vqp4kvImBLEd6xQZBP
6/mCHek+/tyLe1Lu6ASA0XzVgpyQWc59ROvOE9BpWM2sHS/58nxHxdIItcDPtZ8C
jWPtuQ7htBt299ivv3UYxTCfj37wTEuIoZNWvJkm3FmE3FFbNxywZeDn3f0myk42
o4sQXm6/BNKWjqqMEUfTOzpQ3mbA8YHcW2wjmQwhCQR2hqs/ouGiE59ZfTKualCI
dwhzoVOItKwL+nQkTLtpPgrWn65SLQRaKUp4ngiiZTfwGEN9XznThtG4BwOGcPD8
CkL4zp4211W05V4MVxgwO1qPnN0HOvOiEnuiUkA3EOXXB3T7bdUdfm7QsmBju8os
leB2VB3oDEQ0Krfqkq6DfSDebUVar47Kt7RcLrqRm3TSB7p8I8+AnufzQnyvkHlB
vI/zbY5x8rjLK0D7ofTPUJ3Mf0B0Sn40lnC4nZptlIjZ8/koLb7C/W/JAGfdU3yS
snJ/E05hSZwrTGQrlCSAK8aDvt/27G2AAG7V/EUVyijbuS7KtNArz4xQ2VIjiwZg
JgEdGi8LqGIg9Uhc6STAsg5h/Mb9T/SnteL4Q3Ho3jmm6H/rMSkokOGXyWvtnoZY
Vb/K5ghmvaAOERGGTkacBKCCOeoayoMu6jPE/J//XgG4uBOlELdi+Y6UO8Kn/83p
2rLfmnq7UG/oD/XBGs4Wgow8wlVGeHi0TfEwc6Mr+x2j0BHhVI6rY32MX6Gss9h/
hQVGBIzRu9kBtS7dwPWZTB3U0oun5kiqS/F/AywpaVpU59mITpqbIcefdgij9pw9
vhdXh3pkjbUBFhzZ5xduadcxkoX8MAVXkTQZENpTNz48enbGW5CmfVL7uhVODgE7
lJPXNPW5lpvO4XY6VEhhxz6V4siX0MFiY+VUu84KIRpUzfvcHCfKdLkk3LqMEgMY
ipnCeR6e/8sh4C9OffwTq/YM9JYzT3bilpxwtpnq6F2x0twa3lsMgPmQ8fHvRCkF
YbX9DVUzGTXbHgg3anu68SgshqBMTBjxe4aaWM6ay8odKflhEDkVQMDcGi+bJd/k
fW+SMIAxJiTtJXJ+Uks1S7yAPbwRy+UsMLEfCIrnS8I+wHTGm38pt5GRaBPtukJk
6+RpHouHU/5Vu0OK26u3tvLNkJBc8deVKce/+yBbYfjiyxuk3KhyYfZHC9GvzM9r
ilgd5M9OKkf59m08vI4pAwk43TG4s+3dCHnGHKGY7WRD3uUMU32JNHk96ylTB8tB
sVe8qWdEaQKlsGfSfmI8kFBl6vNkolHf71ieKYHjsnsW/phlWJzJmS8Ii5tYK7K2
dwMPGUFNLTRTVQp1V2Oq8JqMfDYA1Rcyej6EofZo3ZDzP4yMTo1oCfAKltwXfwU9
FQ63Mj4EnvNuwh8MNZ13AIobzYLVYrOw2t3HvUsd+ao4ATHa4Aj17CATBxvNl0++
7hoEpW/XuRtet1jIR8OgfRgGfXo9n8kGmOD0I6j9jN0PVaFkQD+a1pGbXvxlRgw1
CAXXglFmsU79LHwxQqcPvh4uY2bryzTYhuZ5sRC0sJfsRqOtxdkIV3eVGs7f2cEL
Kas7LYnpfQKtanHFxGliOE+XYJBHLL/TBRj1Iji6Vc7PmTh/qd1BHoKuAvedFFx9
wdi6LVZlWN14SJZbxlVyT/b4FdHSjdpkdF4O/KnASgy3A1dMLLtLNKUKXGAaTF/V
wm8tB/R+qoPWpGgLW5tOGfKRzFDyP0BiG4MxRkaUmLeedP8A64oESRdQUegu3j1A
NFFd66bM4Z2O4sA4OcjvsiaSovUEPmAsUnH7FYOKGnK6ci4ezQr/Be5raSY7qRyA
6QuQL97yXh13R8FFENrx77OUX4hUbw90LI+H/Abvp7vC0q7Y1Wk4v+CabI6nRrd4
t/5dFny5KFpul77tGiqImQyh91Jl2D53sE1Qkg4ybpjPwr+AtoEnU3EMQ7taED6c
3V3rIARj0ccz6pEI2E583jTLT8dHVL4ZbD2ZE8fgbuX/ttkTmh/PyCsPRLz+h4m8
GYJCp03x52FKpfOi/zaexTBb+JgXUtOe1fm8NtGg7QzsXrM74z4Qwi5XDUFP3e7s
BZ9bNtxwPohQ7RNyBHHRBnt3QWDGgHFpNvVVJ7AL0d+JcbQ0/84af5ta2FZAR67F
hwZJpc5iSiokC+NlXNEDXfMO5VDkG/+XRXaWbcE+f9AVhkodSnkv7641YsFAlyWL
pDVADOlXxXZcyHDzLWOOOyn3iatq4h/cVd1b72Fxsiy70RUy4exSK/yMKURoH02G
3RhxEHnAafoMaAbYfq+0b0AnkT1tosJSjqpCfu4b4KClEeC+e36W9ipYK96e7B6Y
TdBiFtFMO8tUPjdDOYwS8PhmpHrWsE7siGB8xp9fGGJEq4MouLHomyFV4F4uGKyd
qD87Dd08cn4TIGyKYGM3MlogOvrPVdehQL2wa5yjpatu0tvogF/SKrkhHp4wTA5M
yyDmqVG7cpZQndMOLsWzPx/z0dDyoJaIhEIl9bxTeWYR+r7cJNu/Ju2ic6K1TiEx
YGWHqpBTXc0BtRCbinf4VCDuFlOoAs8amS0DosXGA1PluSGQjH9HzG66v82wHXXH
U6h96qLf1iasQhpzb48ttmtOjuWj6t/geiSGP48ZPh6z1iOTq0TExRm+szGRYxIW
m3lhAncMnSk2dsivoTGY5YmroCfoHERdqW7I1552HnxqpcShNYLDAqB6lFSmeSbd
3QAphKu+kD8dx3q9V+WLS0AZyiInDGpvzP6Tm/k8fCwNoOGQ0id9JdHusR8LfKks
y5JBkKyvnCPpC80Ryh+vluBe4BNwdkr3GDMAYyG2WgC0YWcpYJhw33hD/S1lhdij
Zsy2kddJ40LmprU7a8tyVQkRfb+w3DFmtMMi+O5S1TwyyCQX8elqYCURCqVBAXSw
5u3eEIlbZNJ1NRyktA0A7yss82lPl6mY2WXZFrkkN7W0kOM3lhum5GlPJ7QgEBPI
4xhxH77EPV8NW83VIfeUbq+axivzepb7rWhSUKfiXt9OkbrVwP0yNkVMAZvvDeQb
hy2vsQkrxmievDZO+Sa5nDlM2hhFPcfWBgmN8SxG1Elbkzs1x4tL1BA75Q0WTIts
VILboLJbHbhbF6URCJQEs5woG+rKLaefQrpalq48C0okOOJV3bzOyhQ8csMJnOs8
vhGQHvyoyhSi5i9BSQGI9Ie8qqLg4TjTjpcJpbAWIS50vK0jmpm5h7wmCwPezXIB
cKp0HpMjQ3n7YSiF5wQVwleYHbEumhOM8E1ywm8e2iEoBxZJNiAz/btzqo87R/d8
Cna2YrSWnE3z7Iggxdzb2bqvxseCIu2WFsTYTE1I2+/FOJZuSH3mH6nxcfjz2iI8
IXfvMbfYpvUeV6HTllM6ZMwadj5jkhhBZT6jeqZ3d78IWxzc2X3fO+/lomrcbVFG
LNqa96/RRiFD28Wb3EyMhg8+Vr+2+uQyGZQO4Rs8DZrnUdz+QAeao28g8mWiotCG
BjZInqOCM+q1rB4anqKT4nGRmTllYX4BvQYRBtoX9kvySQiZbRCfa37IUQ6PGC4K
GSHWkUSQYCSRjJU//fWXQdsdEK57Ateau6sY04j3nYs2SfgmSt1iDTd3gU7gr57Y
4q1fr0B9DQevWBXsXUMYcC3AZcGNdurz9yphiBHuC9CBYCkiXXBXpqCl8/KH4q7R
5ou2ibC4XBjwB/3qYoieFfrAJLf6qusCUqcFpuyh1/q7J0cmpNG+G5bnL/v6CzQv
AIuZMl27w+qPU5N/gz0YD/4woqY7BNX8rkp9zmu0Wp2d2DPxZoo7A+Wr7BGzAnXp
DYcP5X1gDcoaVyBHPpDWTd2k4dZ/4eNUS6NOPD79QZm307vDKnLG5NhS42BSy94W
C/QbHpOyX1MZcB0tVwU73dK0ny+lPs9fpkokmjvt2lNVF3mVPldPhp1K0N0dTNeb
RfssPlUDs1eIjSVjM+MyRAtzq3JVtQYAEILJSslQ5+Eu52qqp+IZkUiQ+x5UueCI
3V30vCE8ll7z41S+eQW5QoutoemSdU1gm201EQENVMJZrDooVIPmyxdnJyhXt1GR
J6bfyBHMqtsvKiyMFbT0tJ9iLUkXXbSLQliqvc9BQy/xOymN8UPUOLZ7VMZBTTGj
VJq2HBSR/xYW62N5jsvVP4zlE0X5tzi6nnRwS0+O9tqsCYTVU73wNVUy9fw9bT0Q
6BXuemwBpWM9Brz3GsRAaDPe2mZAHIvicHv9lE7zSJDK1NqOA1xHnj/eXKsfOggF
spkrRCo2tBgCnoaWXMDacpVtqcD+cD/ng1kEPX15J7pUXQYQSnoQK60sxIYDUw3S
mfrnEcNg1fX/ZFSVQPFjzmQrls8yBFpEi9cmkBOpZa7OHTGKxqO9sBEt7d81fCF9
fEnwTvmklV1tuZJZqhu/bLY5oaLfs5MnG5qND96TZPxCCZPlSsIqUEUl6tDGmEfW
oeI4EeQ1xZlKEkCjdk0zP/Ct3RCe1go88pBT565coQeetTWIoz4Pt3BH17I1wAM0
gYR7AveKFbg+wUgXa+ENBdIgt6/wdvq69F07aLhMKzC+hxhLNfDT40cZyyTkN98D
4zfk7b8E98prPZB/o/QLtJQCkVEsYXa/66MLV/YdcwSRZwcvkIRZuiT6hFBxMTz7
I1avlPNkv9uVL9kPa8rDheXa5rdbWZrV+1DX0KVD9ZZmakJIgg8NPzacNOdJUHfR
rwk2Q9X0SDtMhkojb9yiOHuVy45xknQVhwbWUIb1YXeHt74NtTw7J3j0mn/VrlxY
ExxMrEM9H+T0UtYPirPsEsaBZfVnTH4mCOtJiOc9cVQRkRe5FpBXf5jUC3njvwQZ
SEuAHQCoFnk1nsqHxioAElBtye0Zo5aNU4cP0cicIHLA0KOVwzApeJjnC6fExBPa
NL673aSbBmwUsgRX2SNp/9G4rsSs2+sLQGIIq1FuaRIGWzi6IM68fVKmEKp6bnO3
PZedig8QgXVBl3qQo453b+Acc46hFjjVLA5/iNGJA1rIHwaT7Zog+CP/63ZUtE2z
1rGrsMAv8KnBdVBg91zLAsAuLD212ykK+XB2nlTsyiPc2M7Fo7pyzUN7IOyino96
0QndzRivQDy/jYGxdHTZqQ8no33hd8aGc+v2GjLPGribaDTEpE4Omy09JykyQ2RU
BGrVdMfudkt3HHrauiLzx9VNlJjT37LhlK/yO/WMdosVF+K2L4r+et+PB4e6AgoU
+cg/I9u0mTsogm86NZK9JYakvDyeV+1hEygHDg1/PnC9swdMpCAhY+jXNh5ceteM
f0vDBRtQSkfUX6mDHo6mAvaYTPpwonQ72tgxRWvW0q7s1B2GrOiCjyccGeM4Vrnz
slx63qcNRdL5Tg4Gvl43SYYSUgYk6jqqkbsYsxpH4MsxnsbHltUHUnIMy1YRfT+b
1UROCx/lspIMg4BnhfX0wUKeE7/ge11vgPRqikwc9BTkt6u3iT3MGBZ4MRghIK9Y
zf1pq8M/TiUqMqPRc6sO6tfzg6+ur6chkQfncrvEWzz/caDGHBjlkwcOSSGjVnj2
PdI1odmaPiIQgLT1j5OQiYDj+6oGyLmm1CXUnHL+NTc3mftago6CP/90GLJvy17n
IFkCprBNAwMANPEWhmmYYmvo3aCdKAIt+TV8NrJ7/VLczqELiHJMigjfz1IFQgNB
IbX6fsMKQZ5gZUNvde9OiHOUBxbJzo9YXxuoD+DOnfjKlwUKQ4yfe6aHBtayzjzi
nvwkSuIxeht32Zuzp1nm8gLpNccSYI3aAvVecs3weSUbaT9G0nfcoMsPeqs28CHG
cmEBiG+FW2Eq0yNv2DDSTf/X4vF4DhZoV7tRfS7YsCjCerva3jppmH9gDBlSMXRU
PqW2+NTProX5q/gXGOL2i6843wnCZ8sNhRd1vrfnqllpHJXXdQJyEiIQALUJ884x
/Z5HtNWyRECYeng3Ar16olxgsmFbm0CxOX9ILBzlgV65WAdi99ixHBaxxisxO3vn
yeF1DflVUhdG1w8CpOb3ljY5LA/LRWhfS19JefKg/OtxKhmL27Ls0HE07L8rh/sT
TVp0x+37YWmCXH2Mr+LDp84T3t27Z/NWlb9dv4BOBx4azrTUeEd0acrAC/C9HPNE
ZOaxB2NyAKC5FczrGR4WwVjV0ArIN3Y1cfOOjqPB3sUtBqSRtyF3IeOyVhrBRIng
8KOPI1Em12OLiV+BdMQ7FICOr2kOV/2zKY2fipTTR0sdaj/F2rxwWe5PaiEm9Itg
SEXDJDTxqHvFewGoqzyOHSa7a6nqUUdC8w3xfSs0R3RZCcST03SB0Is10Tr/HdWe
Mr4hwIII/SdsfJ+E6vRfgVrA5juUZ2Zsd1SHO/yOAkCyupiqqS6/PlJI4Ca10w5T
C0O0urOyUM5Dm9qPSHyPQifrtZwkDM/JABnK6d0FoP+XFiE6iOv2DwoISvuIlFtp
7A74yKUKXSOYK7bjIvZ8kHBI6D4B8u5IN5Z+gLCOBF/YL8I+H9g7inQ/BFdqxdFe
5yB8kGTtPvsfX/lA8EoYrKyUBmUW11P3w/xMPMMIzxfmNV0Acc05EZj0r0blQMHP
1TeDCRV6LT+2iUkiFfZIZP2umYaoUaMLxfeakipGQqh5cGFv2+/Q41KgdLBGg+ib
irx4A57NaCC0DWAzgTy7EUEBdfaPudnQSRhlVlCwE35lP2nhKfPirj+/orGuny38
hQ/dxaUv0KpwLhMURqgaqbZIhQ8LMz8O/2yYp7q0gFM+cgywSu23fUpmJNGt+EsX
a/eO0v4+F32YvVzhTH49Dg36lhfxlpWlQnkI/4Ntw5Q6DjOusCqdFYG9waemSuZf
+v3RI80F5ZI36dbNfIRhNmiGNIOrCarZ7hPXINrS59pwhY2OM5pErNOo3/4qnk7y
OeTKI+GGANT4b80qE3VwW4rSPev2n+WArhbzPfcu5WxoDby1DtAJ05JdExAk2Iqg
nGyWXTO1p/dW1JiwR+N/E8yAoQjtWI/f+QQJRUFGf23C7aPJ7CbyXAc5sSdA0Glw
XpGFBVg9NngLdQS36QX3BXtOKoYMccrZpg5vzV+6d4l/oEG2fglBfCHsbDI3nK5z
jdSkV/hopEhhVfdEERIRzBsPhz1BdO3yPu1iLMuY+D1aZHBwPemFVEzzJrkrQTyn
1nJu5yuby6zA3E8pygt8XByl+/zdh46j04/9eyNQ+/FjfcMkQGIG4esjp5MZkeBT
vm0mrBEq48OBATwYYzQCGhcMd7vhlV2HybmyQQS4lz78YzhMqZdgaiEI26kklb7n
q84jC+YFqhHd7xQcXZX/ZwlscCA5lRWjitGDcI6WStJYEs+nvQI6Ltgr/erxY/UY
wyAtDSOGfzEQLN9gPtl22ZnWFX4zxJLUg50bK1xU24cJp20VrMsra9wkc3zA0KGl
dYcYRplv1OsSMOE3/bw21fbIMj0BP1RjMaJ9QSfnMkOWXuAdjbjXs/22oMnPRrEB
ETjfLHWqxgePeytOYHZKU/unZNDd8QutsFde2t9SaF2s6vWNtNPZxx5tOiaX7MQX
luv8yTV7BcEHk5KXieIse6CB0P6nnthOONzd2GIprLJ05TXLDO3e1xLKlZf7Z/Yg
nrPOzvAho71e6erVXH0LOPkQ8TODo/Ui86LNraHKiH851OgM8ZAMJ9TcTMGa9sVj
gw1XQhbNKTv1fklh8IIOT0mdcFImGvhigYNR52lR8C2k0cgqJAsW1hvf8r1RlXfF
cSBF7kg6SQDvo5dQfRyUkOP5gIFysVZN5Yaimyhn0Zmms0Mur1SOktNVAkHT6QsD
9CUFOxML2otfPKYVQw2C5FAKveDqjrxfCadUR5nk7L914c8PmWG69pz8ad2XO/sR
uYJRffmltitnNWn2iyalc4bdoPQoypR/PXb8cSBHgWaZppi8hrzSS20FeMIjogvj
MSrwqJ9N25X1OhhL29RWuaXsx6nAO9/JRYQZBovPT+hArEyhDEBA6J2N3OL9tXVG
27ueAfgEqVxflC75ngnHeUokoyPZcJc+veNog/IMgrGVoFGOce75X3dli9a7is1T
3ZdX5oFiQCakJBgbPGBL+zF+jPVaZ3Uu1qYMfh0UOAXCfmkf8CprmihKni8AUPc0
UjSvhWfzIx2jHC0M2qoTLiYucJTQJWWulPDYRoABhvAQfKdZ+iUp8kPI5GZeYZ/k
GeXPPTnSC81rOye8heEnYu/H6SMfAOh1Sc9tEWF1girumxebSMMOlSbqKPymhtKz
7pCR6g7EmmDxnoaQSebTxG1s1o/qJ2EX3l9G59PoZWCZUGCMmJ6xd3aZAhz0xf5F
WxI8YNXJJojXEj8FcY7ROc1C88MTTzWIYXQ0uoZCGUlLTcGW+86N+RPpW19mtikW
oZI7SqkwkQjaDY7vE7SROT25+TSQMERTG0722ZTAu3Bl/8PAxZgf1DAfp/Nv6rkz
vO9ODcfiVM821S0YCVAqe6hzBNbmSKThCJarNXSTiyiMxGdCLEslfkcOYSr8mZay
AksTzqAFPKR8jbJWxYlmyTTzweIRQjqjNe8jI40H2v/V88VvFh1MhNbdTehDONNv
/GirufTORLxBN6w6PxqEg/+O316oPIIgWlSnRoCmFF/UN8s15klqJKXK/JyzRY8e
n7BemQh9/Vh/SY4I3RxO66jw1PWq7A4/4bLE6xgQPuiV1gVo4Lz02jHScAKYMOpi
J7qlHQbL8yBKBCszJdNM6y3bGkBZq+oqEggU0C2cnpPNqPLGgiWrviUC9HfRzyeb
R67JK64lSmxf4DH1kVUhwuroSBvkme1IeXRmCGBNo5Bkh5FmLefXkIMomI+9btO4
AxoNnNmcTrXfRiHpGlOlWawy0YuhKT0z1VoLV1fvP5U/PQIzRq4vGwlgA45mlLsa
PPnOfNwzs5GvNSjvFi/p/nn9bxPBJ8DCOq1oH6mJlYChfJD8/aMve6LwmUy6T8Tu
IEJhuCRu22sYJyY1x+3hDv7cYBEAMzyHXQO0jMckns96pdDux28pA4vEQjkpIuq0
ueY7n8AevKmsJ9rjK//rPQcF1sItnSZFpt7/tASWrUg95FxFyy9+hSeSGXmMAe89
Aaqv+hyzptAIgnVOaeKCCBjpU+ku46H5LZN6wn7yed+WRLTv0ys/LLFsDSqCx5JB
D/IgjrMiFJRPgDYR/zPa/irLXOiiw5w3sjweHBK3OtakC35QyVtKcM/TPq8MWDtb
Gzg/7frN93Xl0uqMp4jlpxgmYoAdBCjgQ5WNV5t5JdsjU+DDh1OnzP7TXPMtJ4fy
uy+P8AEQPO+mbk+Dm2O9jjWaYHZWL2MeqPivJF+s1rSsJ3V9vDsZ+hDhU3McECFD
MdCRj1/KDJ/rIfcLoZL/i+HyLzVHB3Ki5yAvatJVfbWHdXzrbzeNRGn/LhwWmtFx
Rc/bsWyPXcU7QrzS5Mvb2yjz3l8ehiIZDKQVMXncoUdwjZR6ZJx7kOKtSCHOMjP7
BAsqk1kjT/oEA60kCfGU1TTximX1fBt6lsKU5k1VaCmXhU7pIFmGoZHHwlsMHbyW
Pyy6fEkcYt27wYtxHrn8A2scrO7CDkkpHhrIT0olzwyLSL9gyQtyd/hUTtHqt0JX
LRSRGvJa/8lTw0CstpnNo0H2WyvUz+AK5KE1CTEZaKaLWfFmRgOxTgbhx1S+Y2lx
grsh8mjjsxdjjowWhS6PfYIZENGcRNGwI4soskcF0ohJE22K3r6k1p/M5h8rv1FS
XsW/FNTBAlnywQ78SGRrK8J71vF7ibQO8l79dUCaVReJ3JFre8xTm1EZeSuTwwCV
HmH9O7KbT3Yon6cBQU77oj8ZsHeNvYx22B7fUcfgB7X70X3XPRaSzN+qEj7PSJMH
eJRvkchoMz8pIrz9NtG6mVh7fP5fRvVoEW7lPvMLm0FoOa7NPdH3S/Wkpk94/9mM
PnHab1hcTXZ9wTJwu3kTkQapmR/Lc3OZnHWXxSBWEmRXZzkDNipkYXEepXZwzsCg
4zUo51tdwe2VYWFGRjK7Lfmi8npO9K3sO2k7qdFFuIAvDK25/yavyKp9NaNuqWte
tIdGrnjQjbRAy0sFgiyC3jOpHw/Rv16aFL+cvC1tbThknU7+Ph7JZjBD6Zhe8nxG
cUaIh5TN0ZdgwFw7uhKYji0eUTrJQhM2g67tiY3onktQNpm9ZgN72GtR/fDKxSO+
9LoC5E9zmmzdoEAj6mSwb6uFuG0YtmX+/WD/fpVhc6j7jyVyZ6N52WaBFam7A216
UhikxFBYRtnOkbebZdt9wzEeAcKQ0rm9eIv3+MfSEOkO7PRcXrY7J9QI+orcgVy4
KT0PwWLa1u3c1HSlUqF3jjPevTQzpVOpS9AlOs0Cs9DD7F0nYNATLTRhyvs7p7q4
OW1r+sGohFzXEdB4lKesGsPxJHf+8/zUawCkeI33TrBJkYsoG+0IQ4dyYPaKdKoE
Z5JvR+75v6QC28WJhMdLIsBVTPI8EIYM3Gxi1lr0wW7844C9xcpjhRWJl8xK0bHE
wuXTd+ZKnXlC4J8wPNdMgTs5gogKuQ5n7ccioZ888Gy8izC+M6WVf7FBa/HaTkm0
xk91LB+jv7SSrWBR5h2BxJWzI5VWQDUSN0rBxZXWyJfYzAxkDMGqPuDOlvRz8O/Y
pPN8bsroARmeCG0k3RKfWQbiTcISNZFYfJpn6WJXWUclWZxdErw7nGM5rzUTQ2pH
ffrR7Ae4mJvrJ1GcIwcajtWg6AjOLXStTJaRqcNvaswTgw+V3xR5+L7yeqDLNiqt
eJHJ7mTbB2qc9KThwQlZNDQwgHPRCGYubb2o3dHyf65bjSo5HfA6ADqZha6Ns+vC
aNN721CjSjV9ZbohYGVKPzIpMiX9D9X+4Wdg8Nt9IH7PKdaGqadZA0ZvVXdiT4M4
rID2g9EXqa1F3qO7rPMaa/OxsGOCugHUxhgLEJILvlpCrtRhwIS2dOb8EBpE/Hw+
VtZwAfciu+7Adrkn/uq2rGZs5v9KjlTPOC2xNAlUFHw69X6nGrjL/MXFa/aeY1xm
zvwf9eYIREJ4zemGaozEH34tkxZqecySJYkLK2O7wu4y/KxNnag2RLvmo0vaY1wN
lMtK9VgasshebHKzbSuMj0TMp3LL8Yd3ueo6y0F63Wh618cxL6iJ1nm8bUH9WZdn
iVBFLPGhWS6Nx0VfVMOf/0xeWjREToz4XcvQHQuKPES4XAELqnf8WiGroUGvsxWZ
hntRIGYHoNskwtT4Zl/2vaZs8BGj09FXT0M08ZEO7tZfypeZpN0OFJW2XVkPgUrO
K1K1eEQNStZ6Nw8HZo1CmNP+YOziq95+EEZge0JpQj+rxzVH+rtJ9mM8jb8GkaEx
LUXlkP9Av6HurnMSzzo6dlhvB/f8ZG45V0ND175zXj44BulY8ptt1Hpf8E+xxR4o
TXMU2YTVaideZvMVTXp3sEnnpGd1IpSyCbfOVQA0QGe+ZrG1r9v6Q/2/fR1oaasu
3WeLemWhuY1QyKlbgkS2tzRLUB7ihDg4Mcjn+jTFcw9FDsjKFeRwMhrp8Nk4TDX7
y/t/lWUv4A6mfwi3/t6/id2d/FsfjuVNxeTtve6+qM8xpYNY0AONu8QsLKADgnup
zJtZPg4sSZRgPDnyODYAz3SMvA6HrtpahHr26s80ZyPXNoIB91C+Cz+TLgLFkXLv
FGXXddo4mYeLKY+D/SvQqiom2QU1sNlJJLYF9ZBkliAIJ9z0LTWmzDWmXFMcH3xf
EZcthiNR/fbPfYIJgKXGasS/yQBxI5QG2UfnPGGgxRnF3CgcPv27fo3KbNKTIaVV
F+9yaxJ/6nl7MwMVqj0gImEsGDKcz270Dtoi+W1SrTWGmAmhmRzaZOx/W6y4e/2f
c26XAzqFwEWAFNFNZrLXTj/Niwg0B3Feq8CZRs7pzZ225IrDoGZNpFybP3VObMDZ
hzqDwqKwhZ01/i1L5a9vEYWBbFhKrSU3cVyKtGia2gRoOzqEz2mMvs6p77EMpDaR
jk4oWzgC3faFiAK3eyHU6rXAq3/3y2BkbK/uLDCEIEeGJoVXbWYz39XTwW5qT2xQ
hub0ZTpmDJY1ZC/+f8bMWPxvE+n2SaY/JPrMM+sskB9jpOt3g4LIPGjVR2ye2ggD
0afo6K3BFsFQxzdHCy36qUx6oWmsIb0gMLtG0uvBnX7DXHWDX5un+aiGeB3MOXiZ
QvvRIvVIMSr9Ay7RLbxrsU9Am+BotkLRUwCNpkfX6n7BNZ5JwQv15kfuVnJr5ZG2
m7SOMPCNyRbF1hCXwh+3ZA01fpBxzYhVZ4tneP61NwxDNxaY/01nN2LcGMZW/jxZ
CZXRB2r3Y0uJ6E31chDeZN+xDA4gb14i9pg5YNvp0c0FLlLofyf/U1MOxtKryr83
gLRVNqHV9lsDS1CgaRBGlwCfbQn29+++oyF+eAJ4iOb10oUKGOBvTdTA99/yhV61
CmKcRkMrVkX5439hcsr2Mgkbn/zM+v7n9Bp9/K5yn6QaRBz9Yi5lx6fG7MYcczkU
syobOLH1e/ZUDqWzYPjiGQp8cesStAC4boZyPeJ6r8u2alNwwOVmjFewZCxuWvgT
s56OOpiQgcH1ZWjhvXQNJsOiLKc17q4WAPXnDKrbkll5T86NPDhsiPNCVgDbxVS3
8mQSj7deBKfxZA3yU10fFv/J7kZxyt0jKXvUM3vlRvCd8p1OlDXvnjEPlP8IELzj
grqO9K5WxwzrVbjd1XRMj/XiEYrriO2sEN6KkpTvGTJWjANyphj4eVlbMVdUl2R8
3zUMucYx7ZjXdVC7A2SIyunx1rmtf1Lk5RyjxigLz394rQBT/qbUFOzljkcrn9wL
5o1k5lCSeSMcmILkkZlJJmkq/yVZZvUlCZTU8fzk51jvBsLtpfyCikHGDu175PzJ
yETq0uWTcjp6hBwyIxKoPK+ajlnX21ncOltAJ0C3+8LtVIK31D5GcZwK9A77fU68
QEeFHzpv93n1suHC9BwnL0mec4VLrZRw0+zvJItT79vCi3PKIBJlQxcFV0pojUny
8pK4ZfxYjVWZGA4NGV8UJ8XNbHP3htbMyalwz8G9F9cmqamjBiTNqhkp3pq6vdf/
BVCh52AypVyMmVOI/tt9P3GJCuUGC4mkkCxqDDEXr55/PPjDdyJBh4d+5Kd95ryl
s9uYf+BXsOBhFaQ/vO0Al68fo2wTI8BjDn2vKMQmr5BlOGG4FxfniiloprGFfAQX
rwDZXF80yOj4cbh+KnXmvwqdNMvHt8nxX/Bv3AuN1ezhVMo4dOvKJXl2RIYW6iz8
G5+xvQJcOD5opdeGN0UKt2XgUeZUP8PcJ34I3KQLdyon+Il7gwcBEm9jG60DuD/t
JwAwnBzi7OMMkDHtWEgV4e1nlQ47Ki6BliPZ2J4ZRKqP/ZBVC6zHObtcYtV4wVoh
CWN40qBUSobwQVo3bNyqHlEOUV2kBQFSbXSYCbSFKAqUNXL7YMdiX9LTXIyLZ4tr
m1IYFqcRq6oDhIoUd3l0EAKrymBTXEmmmnZWO7T/xLYr+MCGymy6x1UQ7dxfgvqd
4M2B/cq7ndx0fo9axl6IGGCCdxGGpafl3jUg6E+4L6fQaCCv6MAvffiz8o+VfMlJ
7LzUMbS+RUUxEZInrb3uwPiztRgBbZu+qt3+jFlpovRnsCJCjGwIXiHwv/FlQo2k
qfQyZSKjQk1Qz3LUZDZk7eMOczT6Rt9MjUbBS44Zj0tMcw2w5b/EMmjGxWHM94ic
+4Fegrz0aj0VoIdGJMlTqZys6FM3T2WCNTIlqq1rfanm14OIHPGRxRAScY5lCNWw
KDSCjyqACn/CsHsRrXswq8V3Ce/T9EDH0KQDdMbqtUxYmmCVutm75j3yULWaPEYb
mitLI4q3Siu7DM+MHPyTCxrQoYBQcKcFB39TagnyaaUw01MTzg0dolLGGdH3QjB7
D6LY0tpXZ+E+atHa05cLfbD6WfasvRH6qxQf1ckYU+TpyGzusjTPqNwduIy4wKoF
jxQzpvwPVufitX2PpbCQuiMzyWhkZw1GpNsMfJG+SzTaEJ7lD2JsQWKx6A1ip841
cD9l+9XsERGOVHcjLSb9/lIXi6xE3mlGiVJC7CTBRVp1bBwuywGj7ljWtpdLlqnQ
hvVRzneouqGRkR2g3cKnJS798jSlfaHPypAqtcl7qKL2pWrFIGJfzH6xvnxkhxEw
CyEncaN83DQvNsVgaxbh09fTgwd3oCnSDm9Sbr6AXvTVWN0xv7HxJkR6Csu6Z6OL
4qVFxo8lgNJQPPP29KWka3QdZ+rv+nXLIUJdX3fo7azbuMbxu5WIXEyaqDF7X8VY
5hQfbyG+RXK+RLqptrI73HTn4Cc2Um9mfczAqUM4RGAsnSlp4niJiuUBvmWkFijC
hkMly0Y2OXpQj2ySX/i/PQmfq+dKMBK2KIdPQ61gKVCQXD1oIZn9rIakBlWVA0nx
pCn4MCTIT0pFQTtxFuFc8IP++DEfw4IUYt+DOz92f9pk1Ixv+a7SPO3n0FhDucwZ
F6MoLvDDXDELbV9gfvmp2L2drfzZUxhMwCwlBq38jwspLwlCOBxGaC51lcm5GKQR
b/h4IAF6pRI3fd1DstnM3K9ggFUV8TmM2CMbz9xNvx27TAiHO2y1c0KKkltlWxVv
csJzc+f3av/gIKmeYylly9V5bwhd+ONMI3kMqyTYaDrv82bfZnPVdq27yH/fPBaK
lSrQhm9m+mxslLeOr+lmasautmnRmQp/g7Vpm34foqdEQxuF3OgrqQ6hKwQWXV2X
QEzvtowW2UNs9DmqH/Bat8V/vjgZphFvPCzNunkp+olOn0lTNWOd0wtMa4/RvJY4
awP2JUGas1CauWjIGilE/gI0tha0aWOu5zJXY/H52I2eanFi/5Bs6wYv8lNeQ149
TVBV8WjaIJ0ck5jNtPf/eolE3heIY/Vw2nZHRE8wku6WRaCSboB8twcutNsYcOQF
ITgn8YajytwpP03cd7mNrxXa8EcSVk9z26NrWs/1Z9cH3rKON821bq/c1lJln1tb
dDi8DeJBUGw6ZeydtwO3oXkwqOpTQ6A5A5qkwDpiaGhcCwaUWt1R7c7F1OsshsO3
D1mb7K1BGK40iywnbaoyCdo5IxxAHH7itWnKJVxHYkMY8G4ZBHYKva2wfTsax1Df
wGdWb0/oV9it4mDegTsMoLx61mlgkFT53ZmlOBfYooAxHJLhmZ8xAvM4io/MXBDX
GIKxTgOAH9g3OjxFUbFhkqUNJy4WTdA4JXczoKFu0Dc535fx5EpT3AKQTKP1ojTy
VUdoZgCIW/QI6i4TlMOJVCGqY1R2oU8H1+XlrJ8e63nVqs//y1FHeURiLqnWWAcV
Ty4VH3Nr2R5TkTQxXGCaxhUm+yjBn6DAQmjdHd7ZDGBJCHq1sWTRtW9g5G2bklXh
5G9UWUiGAsTTudFcoCMGQZBCAOOvxINAV/RBBcnDGAVR0lwrUlAkyFO3hd9/lplI
uR1TdoyuAemrRBy68xf1BISBfgFELt78hce0+xmlDB6izIjpriZlH75T5LJn309P
iY6em6NtJbl93pEe3mR6lr3T4XZr7KpFZnNy8x3daKKv1zmTNMV7QX0rMxyxs1rv
wwKY8WoCZansefUlZADFdfVY8v3EMzcO3w1FytUwoI8FGNf40QeKthCj0jAx1DWR
qaq2uOeNJ1p2gRtRUoAPlkeC+Sh5fGinnESbBpQx/mBXD8TgqsUGxcbeAH8fgSZq
ZFECptNiBVu8n2jDm8SZp+MyCQCsCTDM/5/dIQPos6NJNvHlSh/2kMuaOHnA97tc
uAys8g/BD+Me78DFmPcWAhhKz4LlhpYpoZfFHZgL4MHCGKXReUQQzsOC6fEGelil
bTk8EYRp84POaotcYOPITAF0a4W1F4oAGQGPssrkLgW/Jl0/QszEaRXfoq5KuZj9
lPiUtDWlaZ5D3+014Jmk6eVId9NqsRAUuaoJZVFD1tncLorFpZg/xlzaqhUym+JP
tnyNAhUM7Or6a0t2V98Ad0AiXf4gFx8El/nvb5/+HsVRYZNijuuaA9d6zsUv+Vp7
1sUkBPADGZ3bvb3cE/Cay4If5NK6TehvW1GeFBhg5h3I9u9u1GCU8EBdxHKCTeWH
ZuLxUWYWca5esdZgszgzFUg70t0lsrZhRditOsLvx2vDdIfH4FAZdklHOqUMoesQ
gaeF6mQfmX4QkOQm8CDqn07Hy8c1V6OXtGWO3as/YucspftOuSEkbyO657HnZtQa
FtT2hRum409xe/Q0XNcoOO5LdQvRl3xH9lu2rTRYHi9sAmwWejUBR0nuuf+3U+Ng
MwmzoK0HNjk3esXZ+Y134Qh5SPODwbwu3Pjq87XsA9/B/2RgdHnbAta50CQy+t1Q
03I93iEAYur8ncjgF78yvzRPB1Wnjzt9NfwXKuzGuYpwf/XZaK4SgYZRdRKy3EVa
MgStHgyiorupC3ZPRPmnyW8ZAehotw2dqGNw93gngr51wm1Weo/1fIl0umHC4QK1
Wq0fHG+oy+JWzyUbH+AkMFIPmFfN8132A9OcdDviV362mgmwCtQWlnk7QxNILc+N
ND11IrVLyWFU9c67t9+Y26xyEKsyW+KofSkXlTN2e01ZTpFdNyw5zv0rAgkrl9bQ
34r+dLDHXgvKiiyAi0FOKEF3xEgGNfHpczQ2+iIl7o7PO7Qz8qYq48SiZBfq12cQ
RrmEap4zC/F80HyiBZE3G3ZXgq1sdzpwYLjX/UZVSWhlWhX0NAYJ/JTJwEyYAgCI
wvMy9bm19LW49nDjr4BM5UOAUMehOQjiYu9YnMh1dICm0u85lwobL+bsuAiqp4/p
rL4SV0wpiDFgAshd6Mo+wS23a7Otg8CW2Xyp88AzOTaeyyt66FT6+H8N2039x4l8
/YCM00W/vtV1Jwi+/cpzUE9xT0019hCEy+QBDvhBm4nuqHM1sI9Q0lYfUX89vwyN
2XWxd9bpH4ujf6CcgoXgJ5f8xtVF4tPliIoZSDYkydJkZsza2OsqzctVsTYSqbV3
inmfRuHv27lTv5yWP0AfRHgYOJ5Unjj7BhgnIP6lWGRMNE1U5L5BacDtbDD19v7Z
WfpejymezWy9GnoIMUSzlOq86MQMI1bEKxmFpXbVAwc4mVyrjxl/LhLH+YxQR3sR
BB3kuaJSn+WQRo3+ojME79miN9jeaUBa5/Ojkg7MSRGfhB06+aP5Ggib8h2Ojtni
vXBBT2dI9+xHDliEsNbpaaiFy0atbfNBH9kN87B3wfLHf52WJeUhd1MW5/ClZhc1
9YuaT/DbpzyePm468D+E41WCE8BwJODpTz7mx6ZvOSL7PbjZ7Jn4+WdmeiLCwSQH
OFH9bTYpekP0fdpWWxbMyRMTKdX4yalxy6MGNyYV4fKvvlR87IZEsGOf17TzKlRz
vEutlsjEvr2WlX8WjDhxlHqZ//IpOWDuQQa6PP8NA/cdP99S48jaIPMqQmREmsDM
zq6Cdc2fIGQQcfO1P8JYf61mAwSH3VCXt1VjSzNt81CcR8VBEnq7onw9SOkzm0Sp
6beoc0zJk3ZhLm9AEWpASOOxcKj1NPVcSzwqyLn3y6g4hYPRWz2RXBuUek/G4zS9
ykGSNXJoTMKPP9sbEPGcVAgaUGzR5Rc/qbsQiWYdgx8Pp9XPh3LvNjxsIuoVlTFZ
JNaS7KQorKbeEXXOtaxcMnt4Ygb5nlvKkDUgr+h43ZPzHTBfZmlt1kMAS64bHmLw
5jKIIxUvbr2ijTLsYWk2O7vMXbrjU9MxMeMVRSwHOY+lYYBPCZXnif7ZgRGHufjH
laPSuL/ruJexsBlFHtmpraCXpgVjqPNTaBNEowhZ+tHFGqsRTh44rNlHNFH5R2KS
Epbb20/WII9FKMYocgPnH7yXOD/yWigxBsRa88aW0/I7pb51tJZlrMHOZfJIG3rl
weeIaDm0dH5ymdljmRBtbMdQYIp4+YDpjJ/G8GQXNCb71UeV1n7WgkCCqbuE7Srm
lSnoBWtJ+G1RSpewTHwu388t7ZOGVsH7eB2AD/V/UMpN3VBFe7GLczDNu5GBSG4A
gL327iMLUPjvOhX59+8Tr0jWcMoU5L9knd1u/9ElfeZenEgkq/9b9keaCAqwYyLA
4mFKzhU/0Jf3Oc3mfi9CNhIm+l1pAF//wJbs+hT2KVSU+AxidhA05886C89T3El9
S92gsW+/jxgD4G/AWpGgWsT313CEqBAzjyYPQR8n2jOCPdQsKEF1eVRHBiFNdoQl
c5Ci2NuinPcOqmCRB4tqRvtvo6uhYW8mwwRLdebD28wZyJdBlkyOTi0FqbPbZOT1
yhUNuF7Pcmk3YHvaYB5QTMnUlAH/Gs4V/XK1cmRnKG6fHkUCdL7dJhrcwHAPNco0
CvVLC0ZDZMjN/0snzjhHna0LD3zdJ6IEMm159ROBekYNZsoId1sR97OOe49+JOKo
G/LiQ8m13LcqGiRzvyt9BjGv1y2Ahq8mkvi77rDEMjTwRgjLW5sHoo84v30vdktu
Ct3p+AMxIQHljD2bnz6eeMrWbTsr+/eubjA4fOtSTOrPjblZtAkp2mhBSWBbhqjk
6cZeJVlB8WGxDEsyd9rA39P5dOPXxApWMJuDxnd5OAl6uc07vDDh7f5i8aEzRht+
j3E/mBzrLiOwHZYI9wpYX57H3S84JXCZhhZ2GpSx5lpBm829mDVcA1MFCBLhjH10
mDvlh8+kZBP9nwX+janU3U/OcUIES7/aojoHsHbly8YoaOvx9brcOqFVQTskes24
4jmpGgthyJQA2znLF4MiNsm6PMfX4Q25p7eRCTsZWtXSE1KXJwSK9stCuUsbUP7p
92hu26zJkRVGlt5u/eg0CNRcvC23VZhfurlh1QV+RIHLE9RHfo+2bk/3xteRSizq
b74uLdjyfISHal0rCA1es0IWYpHhK9n7WIpDrK/7v9s/tFIPmndvBkrWHg95QtpG
lg+r1vw1ZYIKZ5R6sXoD7UzAC2n5RwGl3lqrQESGwZVgXmfQvv8sv/t/CX8UnznO
KZwVHFFGuzczjDNpKW8l4KWqI+sure+vKoJEFl+VBXj8ZXK9ukwTmsb1sOTIFT/+
SDc7gl7lmOwbQjzCk3waSSaepTUGTADFKJhjvylpL7dOS1ubqTByZNUooIXC52he
iVVnhfpdkoGzIQsJliFnqbZL31HGqvDBecaOsSHIOOjRSabHQ6TQhntR/rMr78fT
6t+07DEA3Oq21lwDjI2lBi6qKx2lZ5CudmFiMurgpI3gV+o6lg09Cbfzd5tFX/U2
9kd2NMUVDexuSox8AaL7B0O2y908LokTU/jWpuE79q6CFgu/03GJd4k7iQrXEbAv
qcZhxrNaYVVXhjEFplbhLC2zu2bVHAzkrBHW/WudNFX+pd8KTqEiJcJDvZOauwtX
4Jo0mHiLqxdrkxGfTWDQRpiQpy+w1kaSOWgLR5AjDBlh5ud9YgflXN0/o9QyHan7
RJo1zAdMJTjwhsXAg4VUHyzHKXIM3Fb22TDwE8Ky4SfVUslFM4nzTX4kcUURjOK5
tMlKKStc8i1rwAtfp5glfWHaAk3sbAySQQ0QKHXXApuc/+f9WcHtop9MK/2I+AtD
y/zsqQyf/lidIxqK+qwDI18Enc8yKRBfMXaZfdW6tzZ1ltIU0GJXI6YuD74NMVCC
ET7w8/W/KZMCAxEjQaetFlB6gJgMaVaiduu0i88xjyOasa5gbPYiZustGin3hhwK
rvbmq74LMfBavygLovJFfA1ZSLeOvE3dDTvDsr7Pbo4QsPmWFIVjM97D9exe2fJI
LsCEVI7PnCofJBak5E23KRzW/mxit1044GkUj86TPJ/DXlDm4mxZPTBTnwDc3WED
+z9ZJe8zp1zQz6qX7kJEhcdH943hQptZnFL+569WSWFHUjECs1HUlp5IPQbcNic8
B46Xe+TNWYzJfkAsIYbUeXlJfmfQiji1YBlQrG9fbIRv5X0DQz0tYcV1DEJ7GhK7
Mx+jTSW9JG0fwi1WNCrunlYFWllTOBftpxUwIiRITKTQvYNabv2X0qRqorXr+TVA
eT3qSoB2+SXQW7HDq7BEIjjlYIZ6v1bXKDUVYR9g7ujFmoS6154AjZHIHnqW9u39
iyblmtK0jVM/htRT110jSi6rxho56GGBeUr77GfFTA9/i/MlaL/cUh2Dluf9uCAz
euW22aRcraDF+Zh9smASbsVxCLUg93RWiQRAeGkdPNcmV38wYSjIEKK2JiS+jUMK
wEQB9mCUGcOjwJjY3UIS6oqgFDosyesXx1Di+FXticdbOH5l9qlxpzoFFTL3Uveb
yXBQ7bDezIXztlaE/4XuJe38CtcP+v/udgc5Z4WV5C651UJABMgH56uEQ4fQalOE
Q2WRFKxuVZweoleYfuUyP4P54JaXe8flaUMGO22tiUfjd3JuB+XF6CvPqzTHUgVJ
nK2w6zmNv4+NJ9PIqpHElzA8MBx+aI9zjI6HUqsaT8IKH3OlIbfj8WJj2+O6DmTf
770iGl/u2rfjxV3qVpXhOC2cevPk68W0Zdn3CdIr/t/EhhLAeY6w+aEyyEnwMY/c
UCG3NJOMYfaCtneS9ou3VIR55OfEGA2o+5/SvQQAlLwcZHtV62Jo3D4qC5JiTiht
RI21alaivFicbZf172QO1NkWCU5TKpBwmOd9tFE7Dhw15i1cL/RifVzfwi+GOZtm
OXW67IHPBe/49L3a+EqRtNywxXfUpWdwEtYtt3fWt5HpcPnZbYgbRmaImFHpP4Ha
BMfrXcy3dGgavs0aadJZTm8TD4qsfFTEzU32Vs+pambE6iZnNp5LAJnVy5SCYerT
SytCk3xcLgWBX4qi1QDndJmYkXGwWH4rpjbIA0tU5Sq9jw2aLaSgTW9F+JGHNtEJ
swtiTUIR6PL00LBVSNXiyA8Bl75f4x7zm+z+mxnhhuNeS/NGc+sDLk+LMUDXOIPs
TszA34eaRflCi5QZYA0z7fxDpk1X3aEXQ6fZeTcuh7Xv7uQhoO8SN//2AUPN3XvG
016gjHG7nwLl4bbsivUKGSKUCFf3yxpZvuIzivfSmKwOSEvStNhORZvfggTBxZuB
QkxuJte5zHkaFXpY30e/yy6btFumoxvZr/OShW6ooPBR5XEUhljgpS1USlWa4Xro
lnfaTBOD0SYVjaafuPhTEk8asl6h0ekMRvyjcudv2kwCaFoW9/UqMWhpfY+xZusO
8Neyr0ZneRQ5P9lpqLa1QKKHF1nTfBhYDDNiZzB7BOxrWHd5D/oWOgByWhqJT1se
auni6fOq69hCeypFCK0tAFi8hKzv3Ze09slJO2rNEHzU4xFCpvc4rZQv1A2J9L+B
NSHpSm71/RcqmYCH/K7pm5KHX4dgzScT8LzOE6CuDdCplXWHFVeBNQ0+QbrKDYiI
5RsAuI1DECagIeTOFNsySc1BlT8m30gPngc/GHRFgBlU6B41UCoczjp8NuZ7Xosh
Xkfy23nDEzLNHHxLZFE+XWypiFaVx1yjuNdyNlq/CpUs2oKveelZ4GCmfAUgE3Sy
N72L7RWILNomy9QCs0vIGNJvd5h2NzbPRmxAvGY6gfTIIukViFCT3jZhM5kpv1DB
O5LUIj+daRH/ldFyo0nwOvMg5DLiv8M4DdzvZe7FGSAwOVwrv7qgjqaT+aRxnkQ2
rKe+Ag7cIYIf5f1OEZ0jEX4mSkmNE9aBd3QEUY7SeiReKkl0oVQ2sAB4PMEgIeJ2
/bbuFjVwXYR4fSZ7eZdipE6+qiG9lZkTYOKvdVe0dBYbfCoefOIImuYS50GLUdRH
sHXBtrf7TJoKtNQ/xMq+A2MHKJ/gYzG1ukzugxe+iCMKJYI3APwDGT5RXWdmoeOi
IrX7UBMufgKKTv9DkoHwka+KzPxCSk5P8K5LQiBojp/h9531JHxZDlOn/LwZA7mv
OAu+PgPSGszNwNAkGU6c8TYqIOZciT3VphwRXupuO/QnB+jMQCWqt8h4yRSitaph
vgLrgOS0T7Ur/joL5OT1X/3Nkdou+gW7XOGmYpIxgV5mlcDlvx6qW0jHid+JiYUF
54gxmL5kUiHjZdGxeb2OoiCnuSVvT6VRjjSemOl9njjQpxjiF76pUbtRLZ/0whJv
lG3fj1U6OP96bOn5kCvlCkU+Z84kwYKjfWQ9whns9vP1A1M4o19elhN8HdyIPcuJ
m5fW+W5uTGMZ/atpCfY3iIflOdcyzlJoQOxF+u/YsPW7h9yv054nHshFYyaK6jEW
p/v3jTr39qeoY+qx1l4Oih7bBXNxYMxEMr0OHI/yYJUA6r0rx5zVWAASh5K9GLzA
FNUpfZru2RsrBQSDbxOpUVKK3H1fw+hDry/LPsxwosrSm6aFdVo8ilKxi0O/J46X
fghkwhQwg4UnU/HwjEkGvw3eu/5DlkZaW74Yg6OwUjpWe7j3nQIqGxqt5lVnCNZx
nO3im04O5YVkAS2yApN6MAkqTcpw67Voa95ZfgCG1bV1tcjG3hNjitlC+GX5zQtp
JORc3e0KE6JZ3I4QSGatYC83QrbWWD8daliag2VcbJPfpdjJ5Lqn1xUFrW4APo5W
cM+hJmIE8BYbyE/BTvZB76ZQjKjxzZNPZDkBpm/dKAXTQflj/EgY0kd/moeKmFRM
rIXmGPRJI59xrtIN7HnoTMhcrWJ26pJ58pT4Fw8pcCz9bZjVqZRv3WTf+ZdO+GKn
doglcO2p1d+kQORC00PzClE+rZIUyXC1ggMVYbeVfOi4w8QKVZK8DAUyfl7aXDvo
Kla46n7x9TNSEXpEp9YoCJZZpEdf2wSxrVD8A79lqQAIMTurYVNLEZaVP8DIPb/A
gKAJBEnp97jEpsJKMitShSDDRf/Rd+oLQJt1XRqsAxXknUJ1R2rbDtIctWRoxwU6
ivBV7UcsPip9WxV8vsBSi//IDDhcHrsf7Ep8Ca2JXv1ylJaouQj7nnWhdqrBdM9+
IyET7OCc0s/KkhMnArze4MGRaZo4k0Z2oXZK078SKZ7bAj+c3JXbIJCUWUJJUVzo
+IomaNTNYM8rhXh5tzP+CRSO27shoofTcR924pa21rLMpf78BEPcBWPzOJFeG8m7
SMzMz0vihTvjsAvjJT7x/ChYtqV5qmvQNHUJa55ObXhRfot/KQEmsbCmMz2izMP9
lenJM0wJ2UhBh56zR5l4qjS/W6aDCLto1RcnJ2MZUd0MvQuqk73zvispN4ZI7rMN
g0pUAXhTpIwJs0GK5eLy7PMv+Rc7LNn22CdD5SBkDpXo8FUTyAbYcLsYgkzTXsVj
nqLnTdzRKNGO7NFdFZElFvQupYNaw79e0YptzA9zLHKFKZDaOUsQ4t/rMbYl7lqs
XRz0Kg7NwY2V0obFT3J5kQEI8BOobSIWeH57aq57+STnIe1DxxHgr/Vqf0aw9Agt
KZXKzMvkF+340G9Xc8phfzOqPtew0NuA2qhDORYGIiw5UJggvgGzE22ctVpq4TKL
7QoPg2gecQ0KJxl0ip1DwdlLt0YD1+LKMTn2X2l7KUDRLVRVUhEWtFKv/g123gg/
heuI9TAWcXwSbdqSpPh4uMg0/iPv5ezl3gq8uVq2WbWFl496FPpPbW7cJMiqxuy7
f+QqJtxTmFVKhVeP3ubdT1fBKTzubhts+tn53xHjJsxvIMmt8CE5BGhsOw/XXzq0
l4E0IpOlpEocpG8j0WpyjfHTTiVl7PkOV59M9uOLLiccgNAK4DLTrLItAHJeFsiJ
ozYENpglBJ5ajOVwhrCapT6l5yfU335c7E2TQHuq+i+plwCN+12aSxECt5m4jaG+
xC03zciyudF30RXr20EVEXqLd+3YUogoAL87CPjgALCKVo9n+7aEz9jpW2Ptppfz
YrZxuqopyc4m7apqEoHAqFPsTozHSamnH6TR8z2WnR5/yldW2Eb30p1cece0UCuE
xZWlQmCptPLKqeW2b6gHgs231ipEoaSNbDcaMYYMSwhEjU9QBFKLFck0CunHLH5Q
rcAQjWPVDkxz0H1RQR+rDJ41sIHCJjzOuRlMQgYqXC7OU+HnM31sGclohOxK0L/A
VDM9GCs89km8dSj2FjuE+EslO0U5ZMy/VN8eOgEc63xXnyzs8bGHk5GLi3Fr0iS8
hQOTrt0+5OREj/3DyYuKs0/SIHKavhPZ3rBcPVjR8FrwDhCvv51z2F15TJgXUZPu
Yxli+jkYdFrGmKyCarsjv4EHdVbyWRzMG53YmC9pKB+TvKzvRTsBY+DNLJUr9s7T
ZUVLDZ+Oi6eUuX5Cw8ptKXF6sZuh3a58RzVKQvJhBBM8O+XFtLySrx2LM76cnljJ
mHyZ8PYVffgB+p+TUg4V1T2BzzR0N60kaIbEEB+AGVoDg3C9cf3SrGI7xijew+qX
cJldq/44bLnwrZ8ab3a7DCpqcXqnUTWj2CSQ/DpSdGgeLmD05K0sPQqne1y2GF6a
ETKr6WydfcHQ/pq93IpZLlM7x/6HKbjBLVEJ+HpC8oNZZxwlzQBwoXlG5z98HJ2V
BA1w+NH+Q+/2dCc7A7mRuw6Ko8y/81BBEAVVgT3bPnCjvEeHFs13A8Ewb18xDuei
ND4G9e3MTPW+ZVRkEh7qzMUzQotRDiV7d3WtkYGCXueTc/YBI6+GGpeaVcYDpiBU
0baU03Fh/Y9p4BkxIqYEFBlaJyBqaZj9SgjRelI3mSSzqNs99ToGs28QuHhUPj3z
bKknT3lyAnNcavE660yd6n/Tk/ngVOHosinMAJJJlMIhkt2pxxTqohgKUPxHQA9G
IYz7MemfuLnPmic/ADp9EREJ+i4mtn2AMYsjzEyrV00ixD2+lpOlgg4zfn8xrE5g
jOUI2IvZNvtb9BQvRfCZz4cYNjWGpPsavys4gWsSmHlGC4uuDRWonYDURF95HahH
jEs9YG59sRDJNmnwAaq3lcv0cjrR8n6UFI41StQAK5wLYLJ9yiHGW9y4wAtnfugq
NkjsP9eZreOVPwBPD6Q/zmeH+QIV512za1L7+YCxKw17dMRFLRa5bSJdmr3YnY8n
0LaKoyS4pDqZIyeH/+pB2kicQdXDb59J/nLmNB//Mdj+vmk2Ue9vCA9G3bzBZps3
MdnErLUHlrqbJR0NOi6DLUF/iLzTZ4dNvhxpcL2y1hKjgEJY9gylZI36a8PkebX9
xCGS4Pei8RnnvJptSQu02tzLDvC2Cs6pErYtF148s/oXV/GtVuOWmgzwVkzyDb2q
vkNhF3Gs2gEyv109K4h0c60NMX+8BAhFcEnVpA4qYDwS2FZA4hGhNdXYdhqHJXQ2
POXtUBzOfog/j1WuepjTl8JFaqcTo3lS3lDeBZApwiYD9sQwEsdQw1iGMbvCkokJ
M13TURFcZl+LtrW0+2UVaLvRXAsBXE1sQawVv+cNP/OOT+oSfJNusmx0FOzBChV4
dGxdzKDT9S9hKog2c4uRpqKeA1BK3GBuDrW6Dr1tjYRz5bzwb8Y+ggFy/3qGWQ/5
TT55X5ZlqyDUg4IoCfjAu4pfWpoN5Y8D2h1U5ZroemL+5hAD4rM7iroH1JnlKczP
NBoodOiI+offDIwWdlbnasUCoGRGSoKr6anG3VNdDx9FRhh5VgRZRoMrbNop7m3n
dMMM62nT2UjX85EItEp7IetBxgQqFk85/jHwrthPeuT2MCPFp+ZQeGSlXm3sLgJF
vZacUpDnQ6nf2asenoskWZTMvrWw2wV9wVxZy+3y8cadfphy88xK9tzoG4BTDCG9
LeCjYc4Ip6tf3vB1z5UcjC68xNz8IhSk5x63BHciQyHEEtooCLGj/XXsoSpkr84H
zCFBsid/SFL1tPljFjdQlWibDXb0cfut8OEloJgSSJ7stNWvhExNCgui199cxOML
QO4dGCAwhsFYtDMywt+mmh/QKsxu11qBdNzvaYkenACN3nR+pSA+bUZknWoPmCtb
RyH3X0WzBaWzyGfSDtSA0VaRYUGpomtzDhN+Up58PCOhVrDfeXv2VbFd1X+hQAOy
c0DBsGgdlxxRzKeTpWdR3uss5kZ1GWB5oCEKyVIaC3h0jq1slmLdArkSTwkutHS9
OXoY7ULlVPAW/kohCEXFzRsLEKQ5BnFFK/EWL+qQMo3Bnag46IC9o/vYFuMveISC
sYGBEny86tS/MFHgu9LBvpuPSgcbEPl7WuPg0cHcc7sdDxUXkgWjc9k0xxFPxG0d
37nEQL4eB1vr3nM99ELcw6nC/cKeJwd7sSaVbmK1HjD2rztMDTzGyueYqiJqEBBn
WDo0aEq3KyOjvIuGuA4wl5S81rPZH7cWSfmmPeVBrCbnCJI8Hr4F7ydnmHYCAdFT
WmoQZlHLU9v+R63OkC4KuSR/DyF9LsF10uNYXCTCiETf58cp8OYWFVQYMgX+3TDn
YSYMOaCD0s3lnsnAhA8KCJXbcTAJPJ1q/L2Fs9vJ1lj9jAkYG3eZAgHaNaJ3Wuqs
VMsJDi8676E03UC6c6mFtCBc7ojbVMZwxXa16jp0j2xRbsByoys+B2bs054ru5BY
UucH5DEmL8r/boVBaLS48zv9qsu6cI1Uddz5+cZ+cGJPzpyVE679M1FfUJT0qGkx
kMYfdh8rTSyMTjp5RDoxdcihS/HgNG/4u6D2lsNtaGibUy3G/K0F4v96I3tjrEQa
+7no0uNtxLr/CN9mp2+8adsDCreqXdah3i2m74v3IqOwgxyDFYXolR6cbKsROQp8
tL0+FrvXChgLm6ul6TBVhafqoWCXEanQms47sh/qeIE9h7lLAjPhWJKUMs+xLB5m
5zxVsHodu+4bvfu+/T8lkph33oCk9+KRekZN/KRv6IMCf/E9nFjCOghBPwdHCfv3
8wqxpzEy6nnXawUGp4c1MjygqaqtbDwaLOPpxhaDM46JPH85spHcIrAwedmEJnMK
DLOQSo0DH4VCXxUy5FrQNBGUZJpN9HcldM/wYSoueMrTM+w+t5qMm/MhmukbJOaP
pq87SA293ndajDKje2QzbVuoEbceSLM0ej2kb5g7cJyjp72ZyuqWhzYVpr7cZYof
DmLOGDqgmztVSus1CAA3HxASoEpQyJnpx74TFI0EmcBPEo+Vd5mx9R1/j+3TRd+t
ZnYzQRWxEcwRwSZ1Eo/e2euaPxABTKrOuYUThWQKdVmgzrxC33NL7M1bKnPbmXii
lyd+4LSCbmRYdtTsaxKqlb85QXWIf/aG3DbXBZzmZG8+eqw5DoN2lzH2wXuNUEqq
WTlacxcTc1So0lJd+MYo/Pqn8KAc4tqW81YD+E5PD0U445cLLj+jP9Ps+15fazx1
Cwx+DEWmT0YtCP8Ho/ZqBoLEQe6yhdBb3ObKbm4PIvXSEPaib6jnRiRYO0YyvnAe
wf67Z0M8yq+5vUn5/PLiIJ+GR05crye5vHtCzmaMeNNKJfnJchpY1uZByG7GHKwT
eTiKiycIrbLWlyriFcSki85qrmF2mR/hIfDxu12v/eRs96idAowiHo8tLXAOlf+v
r8nFmUyaJmiTbvReIRI44NJyjJQvAFhKT4Z/6Sng2FkMYSxJm3t+IaayDSwXS9dl
U7yMP2+fK0pCpAE+De2dAUaL9X5mN2AUXsic1rLMuFKfMAJisedkoPQc1XBjTvhY
+Sxx0Q3kSK/tcoFB8Su/2Q4YY9GGZZyltaXNdl50ttrIoHIAmJiALUbh/yV1nxVh
+Lch3ARFD0+dc0spcAtfcupNOB+Mha8jHp8wSoctj61/h0z3aXSAA+G5csCQ55+5
6ZBC0WzTab2+QLihydIxmuypL8v6c9cnOYtI1ByBRC0jHEl1iE9l1FSCamu6kVpd
+n0sTOx1fcngRkxUzf3j7ZLinptbiXsUhxCoDTBmypIHrRBWxqtqTm3ONZpVqqVf
U7fyxMKMfvmIzZv0GuR1L339CisNJfr+WB4rKw34zEPoeUaQFqSRHW6CBRmzY9t0
FrrkUAcOEGMgcs6Wgtn+s2k/EWgG7iGEJGY6MzOy8+7w8A6l1mUbBNxMeAOfruwE
sZlZxrrPVNKKxjQJccvJ3CVQ7MNNO8WkIaimJyueMrtwmtEeBSnPwILjidkVPsBD
V6dEWHM83Q5bUwwm67e/13z52cbFtvi8Ff3EDpC4sw1qHrkEXCqlbI4rC4I9Cg9p
uPxXzLsAMgll+4vd5JeaaElIn7S+rQ3sRgXNz9Xld+6LKULVBoMU28Fitswp5Qo6
s0OPlegG8i6Mck3rh0Vn5ZxiBpw8COKcMFTQqoy0rpvJsr/GLwP4uUZxYeK44dVh
DP53oa6WcEYraUN4AVG2kbLONPeoYsPAJ/iaD1FU6isodQ2moAT17Sie8cuPDdCC
aHbYFl2eFRy39rV7qH2uvcdk6rWYRImthzYCuTmZv1GyRTBzRiAhV2ZahArIG7aV
Rz35j91sLuuTbSWCIJBRBq5lXljvv1aFY29rf7UEGMzW1A1Vi5ql4h+4yM4yDXS/
QXlR+dg4mc9QUaw04Sss7ipo2f6AwAppjlUFuE9KnuF7F5oadCmUyXFbNXwOf1Kq
AVLDZOSDdYZOHeREopebasVMqobxVAWP6VGtDQ+6faWOOpwcSTKsRxJpBOAPTGsU
W/I/32G4nk7ciAco38B5WW2hF/Rab20zhWszXtXWH9f3wthjZkONqhxhp0vjIhSU
UsSID828Q4nWoSU+qfgSViyk9XVhacBeS2OBUmLdjnw6ot1MLii6jjWgAn3rZ3sf
zfUWPBUAo6YRcEHONEEtXErzgGs/ZsT+D2hTUUMTAwAAPVHnKTJeGpQDG87dICy2
wTAL8/HhNU71JCnrfPcZ/w3Tzk2iAWzd57UZ0+kkO/hW9iKMEiwiCti1x+WBaoXq
oQS6I1O7ejokRab14fzqXxIELUiywmed9/Ss7FnOdT72pVSeqlaMlGVJnaptt/cY
ZsQHh/yAsv1f9hfgVL2i/Ht+JwyXSNiB3h/pAM61CsHGWNdqtb9H8a+OKahlke1Z
hZpZkhdH265WzTBxIa/9mrIskMlfFIx0XazQMSTOI8z9y+TKx4yLKr6xNzzQMWRf
7EdnLB1sXVa788bDTqN5a6WrBBCSLDpsCSHWU4xFfq+TkYz6tL2JFluUFmQZrEKJ
u1VFGWQPv9igdWwOgn+iqGzQcVGe1LDjMdrqiP27OV9hVIJgXFeoIM7T5mjcmc7F
6XmtlWqGPTB+oXcoKpkeb+eCkbF1F3/ZwI/3XnDOoOSdan5psMkf+9cBsBMdgIay
fMvJ9XiizbhiOiosw/RczPBaeLi4oHKH2pSKClcEEbF33YlD78xukzePOTmtxhFW
vWAMi3G82JRkUKUxjDkAtdWNiIBcGrib1YcvzxB5gg/ojTylL09gWLeBW45dDtoZ
nxisNaS+9x5Gpua/7d+xMWRUr4s0eGl7+8HkZpqpwrxlKKWuzIYkIlS7yQdogb7N
L8kO9sZnrTvFfmSyyNfZznqG/DTnoYxP1blVXsyAq0rz0ktPpR++sfwnMlfoDuFt
P491+Agl9cDWpIIz2J2BGy53M0QKgUeF18NGPGmmPHzPlsiXpm8V+KeI812XzHfW
J/k0DtD5w5QXkxZ0/kh1988hI4FRf1M/mBEpd+/di5CEDjRCNppoy5DNyrNCDnGB
h+GG8btTCz/OcIB5Hqctu15a7zfgm8p0eMg/N+7ZvSJxwk3m3RdbBvsZdQpI3AK9
0E41aWB61ZxvYtJqD1zK2gvyc9q7yDLIoWc66JXwyI3hRmQM/qqVdeglaMtJ5GoU
XIrLpcO6GCBEIgK0avTdnvcW2TOx/pPbJE8BpwSafQjBWZ0p4WKv8TLiFnBPx7Eb
VW5BYH3ZC2GD7sIITZUGgSnBTfH1VHaazSsyKf4ejpnL8RxJ6aL6w/fGKbrQCqK1
0nQs1bxKDOXNpelG2g9D7dh1DsN71EHhCxIOsCYgiaown7H4V4uz2qP9VJ1b8RWs
fYU4QgZeTrtfonXpm9qp6TKGM020MaU07/XEi6XBM2hyiPdMcwugKNvD/U0zQUek
zCTfvpYyh/ifJ7vls97B+5EXmEUNDDmxevGdN9OpXi7PlTyO7hOP3hnNE6Ad82n0
3AmKzDiWn24DPl7z9Yuywizk0wUJgM/Y/pvN98h7qGdfnwlGftLSAQmp8X7lJEAf
zySFr5lqZwxLG0Q8zJ48ELyorBkD6/4hyQDhyuopLtwRTnNM19IcbtHEeno6eJpR
GCH+YmOhDCr+ieOAdvosqqL9Ym3vrPiFjBiFGnuxIaEwAx7ZN+JGrVcX9bEKgvj7
gVPgD3fPGv/xoDfPgi46l8OGcuaVpaFzwQAPlHEXIC8e80uKO6guBiacaOvhQ8X4
TZ7I5eHxJOXR/nToWSOJdsxWEd+4JILv7wXY9wH+LunSahKZoPSTEmi73CGw8Ee+
nBGDyRwRLPZHaBu/rsBSmHMdZjgOyvqjA7ML2fHEyTTnWVNfYePCXnUI5xQI2g7/
BW4UqdYHUyI++oAmF8yQ9a/CX8ogJJZl6Hl2Q3edcAyIfjkgFgSsyO2wg7Xhy/vx
uhugheeuwARQdxTptJwWylyP7RlT3Gp8HnJFamrmpGQ6v8LtkJicLic4XdVy6BU1
91tbNRBcBuc/ex336i9hCpvwFOXsqZUX6NVjFMZxlFxrjNU1O6+FFa7/WX4Mxaw2
sUIwwf9joIvWGIKtFBXr2Yx6/LZM2vgIzr7n7NOK4nCpELjUrG6d/a9044Uglm6v
pMH7lRKuVbThOwNfM7AaLKCxXx7VBr9PEo9W/FvCF+jNlpTQ0WU+unGDSDPhaSco
HU42xpSpPFhimGRujjw9oDYpbZMZ86QuNaTFnVjVfvPugYOYmrQz+5wT4M9qu2HV
d5/WmvHXIjyFt5gKZhdNM+bsZ2AB8wk+o+SDOgjpg8g4QgawI1tHFcD5WS2TdBLc
sByJdLxnxLBr0UwQNSMYQqzRakoG8QZyh6GKMBhRSmcb2M3SyMhpiDLDDmwj7QuD
E8Ky5b/4fn47zdNYiaB3JXwWy/YZ6qQRg+DrB3DHD7Sz18YPl42lge2D9kHw8fwe
KNiYgxayYwXLD5q3UkG5rXs0TZKNbSnKYWT9EMP0W7l8S7EHA8CTrVgmH5YiGUTD
idR2mPpZQ3EuHGzkiGnYR5xxLB14le5b4deABJhlVJNN7oz2UlImEXbp1TYQpcLk
4OZyMoWDQf6258SSgt/r99E12NIQEAy2YnnnobNLRMz1xhQxtEB2AKE9niIKy7zq
HdUh3yyEs50StdHa3/ko9cFMme24JbsyjjYcokxtge6M6pVky6gIpXYqNK2Ov5S0
odTmMf/4LednPCoo4VWI/ftNvLSX+8sBu0zLq8TCTejuNW71bQ3efOBC01L/CV87
sIz6K/6g4z7wHV/PeB38IwcKGhPEwZw+lFDtGr0MDn/hpvT1nFf3bjChHvshssMh
lQptOteeyJ76iV0pFn+3U/VYURwyXlSQq3xzJsg7XWDS3c3mFN7OEb26XSJM04Wl
tm7XvOwZbePLki5fMBzxEI/waaNDKU1PrUt4pp2Hf42w+7Eyhsixrxi6MpRXlMbG
H+VhUyVtH9+7KloHA2Pl8t65TTJ5GUAxy/bX7mfen20eGRCr/6tR1wCES7DTMAdd
Z2fcAh4PHWcfwkZ4+qBYMz2vwh867ef3F0JwIoNHGLwYVTXjQgxfU50MmMY52KEc
GsyecFRJqRSDD4lwNC3+pmm9oW1XmMuJh/V9fUTNWjKt9WkiXe41A1e0FSwVUJqP
dk0h3uLAdM/JuRVIyLSQh+UDSzcsU5Fm6JelRenvyf1EzPS6zNmXLpX0EQeNKLld
Tc1sBnlI8JX2tfAMXMX3VYUQ1gt28l431OJii7NV5lzoQIRe3vnyLfEHRyOGNEWk
wQYQifEZvRLM5GDjWeyhb01rG66cy8Qq8cRKz3o6wVHJF0LxjbUatHS3LVU9tezb
V1Y2T4LPlArqFLKKTfQVtldlZPO8plXCWtThTJBSpMHYP4CTonooLlvJlU4lyQtX
eK5p7SpkICN/dnXD79yeq+Zdjr8gn8bWf+N+sd0/d1/Uc1LGiBYIC3Eh2M4XwS3U
RqP3KMj0EYPCXnT+vrGAhR5+mSpY6iXYZ7viXFqnZx/gC43dbwQjMsmTtsryxWm+
MPDOz9kXl9d6XdJEhi2zESDrjJzxUijnWuTUDF+3SBwOw+bmbRHbupqOR3wpxlFi
TAQAuKgrdcZPXvfRdXr5v7FP6R5TVLs0X6fX7q3EFbQDQDE2uBbRcYLAZxOKW2To
7zmZepGGt6IPcfIjxyHcvG07U8iSVLx8nrj5ui9DkqYS7XO9l7Ix9ZsoA+h8WZBi
PnGDyT+WUx/39q56PesEOHj7YLj/ObKaYNd8R2fsz1ziGU+eYk3RuLOAUEPvK3AH
vhdziO+lZudri0E2vi3IY0nSfV++GR9hhGAMAPAGHd6D/mVJeagHMO5gW4m+5ZCa
/5coq4EUzYQWcQvHTVLbIdpKcR9QiZaBFqBKGg5KiyTo5QBDtRSEX0iUeMAZGLcP
jA0o/cvcj0XnJSEOTS/5+u7TEo+WU/Kryoog9OKEm1oH4XC61C0ZEdy0qLW313yN
pGS3qEgPPksmqyoVvoBwIw69Z9zcsvah5v9ECGNatA0IuqW5lcMUzbsAYOD+7t/B
jxqIQ3u0MRQOrp426zX9TkBC7eAPkoDi1LKKAY6t+KEOATfCGgLg+z8oJGVJHViI
xu1nW6ddkXaajwtt47TE1a3KIGBB24AGOhThoR6d9CMs9BtyIkOOrOyBJ5mP0iWP
ESIHu8x3yb+uoIVXDBtuiXsYpqfde57a5UDUw/whVF85kr2Yf+QcdVkTnW4YThrj
dC85S27+YDu/4hY6gSNfSCryv9+oXu7T2ezRVgWPuSfjT0jOz+h3/rcPA2D4/2Sy
uHcsM+b4xSccRLTCY3/QqCMb/OcnZkFqLuNijtN58W3BMW6fS4RBFtvFZiIjXNVd
jDv22U4qDZqPQ29wXwsuYYvrYj51ZegMfTnPV2jLf1qNEAbhjlQbfT3hl320yLjP
0EEfilp3IfmApsKor2Y2jsRDWhIsi/MLDC/3MwPdbYKi5/SyssuxkCRTuCHm2j1F
SY6bBdh83CTZOeLcY7rhMz9L50NTKFV4tiui9XfHbnYnlrHwWQIT4JbUVpsH7SWq
YPsMUlh6C2LOo2OP4+cVqn2ywkDgUl11eLAhs6eQ9KWMzTOa8/PMNa3HoJhMcGlJ
21pjcuvjVsjrjNuGiyb+JxiU/EhfMF5R4msjfMYVIB+2YyU4buX1ll467saTt7c2
bP2xBYpfu1kVR+Rxl+2d+b3ImoSLwVdVp9eh+6RUR5bqlHinYeNHF0bxBEdjAV2H
9e8l0eJZ9LuZwWk8S4NW636rDhYEdBNyyDDjrx4r2BHO7l5kOaqwfNAS8thucpCD
BzPk7le/tlOiI/AeZD7AcyJ57hon21LHIUPMNLXHnFTkv5X17W0y/pJJWUlHGjvG
OR6HevMhdvr6wvBlH9oDvHzj71984id6IoP79H39DFLY4XpDU/5KjIrzdh9BKQAf
9Q0ws6vBaGULqhXvFmTp20Lrp9iyLOexhDFVj5ZIWN/08BJLKSIIoGrpIGoO2ScM
+ymhY1WKu3mO0tlsquOoDKVsIvn8ZVg4c6IgIqV5ZglBWxxdkbZ++0JbX+tpzf9K
Bz2tjZsdL3Xzm885qkHqWaTNKOvH77QD6nFb1w7zGS+IZ62oYr9O62utRH7H0olU
TVhOpvZU9Re1kfgXqtWSzfAqdXKflQ9dtuMb768D80MpRUKoKsSXKayfhyscJ7OC
jDefoCKQPQf9J2gDs9HXGoiRv8Tp4rRRldPDZN43Sb6qFAkd818kcDIHZmDt4gzj
tz8N5XDxvdT7nLwr5+KArHNiHMtPRIUforGEBSdJwwYjZz8fwGlmMzAiXi3ysXny
1u1/Qk4aTwBEHQGwxcSS7JEgESS4jOoAsloUkViZ8gftdMzzeCqHtqCerLxb0csa
XoeZa6OEn1DrMT/esWbcG2lkQDWnLdjhmWUZsD/mbrdp5J4BOp5hIpu/xZ8p1GvP
ozyk93C7/gxoqVzw6Wp1bEyf61VyaVZjhxPmY3CzD/bjzWhpa5SA+VQFDONPaSLm
j3OiDPCfofS0kil/Iu3e3dWKU1PA8EA/f9FK5qkFOPotxPJXxpt4DedWk/urB4Ml
l+9iKlEvKb+ES0iuWnqEugp8ya0qqolr93Rc6/gwzkT8lANRUIUuyI5pUKvXIsau
xVKYRvMnE06MXzhCwKG8jmwPx7UoWo7yVzldZipxtI0KtZqxQcjX1hF0w2jEDAnx
bKGy873GIXcqp2FC3JQhO9/fv8F4yWpuaxroAB4FTZK1RqNowlB0lp2n8PoBxsit
fjYQ1A7ZN2RO3iiEF8zBQcTTgHUgw7z+h/Dmx/Wn76IpYuYFTZ27JqgPEZmIA7MQ
6FU63SWEe0uIlqwIhqmq3SV9+GZ8N2DUnxyFZv3woRr8+fz/DtkXgoPdP0xkiPcb
DFAkFBb0LNZcurf2MS8LVJZGVhRJX11ms1YmG90bXgrAi920l373vG6zTaw3RkdU
8TSf4E3qbwoXpx8Wcjkje2aHn5xh+gkwCKnIQLrhZfWm2IARvUsDBZfGlOng+675
QPqTfwrNHpAv1vTRL6OslsF1pllF6Xw3ziiFQzJZTP69MKlnD7HAbIfgX1iP1PG2
J8PkZf7dxRVnjCNgME/8wODCPY/RpbRTtLPMbVmFzyrcgqRmuWUXnHSk/KXWAmbm
zmpIRP0chrIyK4kVD3GwI2i/WZskZeO85QAl5Aeabo9n7NuqwNR1pTPnqayhMhkz
IjKhDJyjbGKf+zlnWg/zOlLS4dTjYih6l01NHhvS3of2e/WCvnbMMv9ENkF4x5de
Gw4v6jIY7CY0LbJwq2EYqlMqZk5U6cscDAzQo75cbvG0L01BZleoxhGTPMNexyHo
a/C9oc3M/FENS4Z+PzVmmBjKTWIZ6nPFSIKo3EMsyo7wviD2JK5P0t9iAmI9DMoB
KUPGndNLBfliouqaiUJk1fv5XCaMNH9HWbQ7vQA5d7up9x4mo0WxGSN0r5IgDmyK
WxLA+4cqoKn1aPJbj1s2b2wqCpFbBs/rjxkB8p30J3Wd7q1rk7buDofmMZ6VaMR0
BQP8FtWK5wdjBkEAfirkybnKio26JBISliDhVGNfIiynPclXjfJq9MofIW1xkftC
80kcTvj2MrQNzfdoyKRR1aKoVNaM/NPJ5SKlxeb8ZO3IDbJcdPGe1OU5Z6ZveWT1
fCHaBJdbpINwvBf6hp7zRDN7Qoz59VLuHB/G8gOaOw8g4lkC6XNziiaL82ZBNv7Y
fbkRjXrzGqxuikS/q1f4ZM+jc+MedS/bSA37kN3tH5414T2XOE+vo4fsUgoPSRs6
0zA+UNVEXvLFSdmT4gaUd5S13plZT34z2wjq65UnRGbz8zFqbJBdMmKOGu7vgBZ+
DCFUd762ARO++GIhdIVnn+iC3ZyhgLwqOLcTyiMWBBPz/sPFTPTNf5MC/Pm5QQD+
6S3VqaO5FMOfSOMgnGVh5CkhVwRkfT3sQRdeGfpPgfy9AwBJwKppRhUY8Wkcq2ru
Ig48IYvUQ9U18P3S4olkSyF2xXhUrZuDWMh4eHrLYkBMuXblivtftMwQJtpbSI0S
/W9O+RDPY8RTt7rfCOaVVLZxAcMpUh67duvLp9PLPpmH8a+v4P5xNIvylDBN35PE
atPsuKFB0xv97eQXdrWnII11jEfod9S79DOHCawxfKdMTQ6Wa8OT7iRFHqvSnk2a
B3Ye5i85SAZMl3gqLpNRr75yUXN16lQCbtfZbvCAWiO0iHn0U5PlNNyqNpLWH/OY
Z52B3A4zBSIUk5y9TUYW9F8kJ7ng6tG9XPHEnesZkHz0tGzKFz+KxyOqAafaw6kH
BzNZKu/T7xErPI9rhBEoJEw3WYLnh1LwUa+yhZmUohl3Dx/0DVvs1G3mwndx8dEi
MGB77JPpPX/FCyZ1rIKf0K+NBMGweWFw96vfKqtx4K9u8utbGQfrQhVDlM+KFbtw
rbLEUo+ctBuUnRz2vSDnHl9uBm9v87fACf6HuN6yFpeLn54pigEnGTH4IGiATYTp
UEGGLiueBs6DerJjndmWKFtBSWquseqZ75Ictz85xPv/NdijverbJNc/6lKcfmm1
G+Cj1uWN1ie4iN+l7DCpUJyKeoo55+PFleRpulDu4pVqVYkLMhdOqn8lAW9h+rPG
BAiYzrDqKFzxGG+02LQqPay6+dMAkdBH7skDA0vPe8eVoAbIiTBKAmdvyk9FW30P
UFygdZ0QHUeBKEQ56VdljjmCENtKMxchSUq2f04VhFBCbNyDHD6GTH5Kftr6UCrX
QpMsLGRYFmk/8yRfyr897u+y1ZHOGwhAovqro5u64ElhA47q8rv6G5DNpbUMtTqX
vHxSXxsWXFPiHYRDrjTXEYJ+Pj2xbuEKzZQyePonyQ8S8XC/d1Jigd9mw/9q/OXV
ETbKgmf/lJUkgSNBNhU05IUv4KCLnHVMcGFGgJQIn1aPqlu3QyDspm+e9BiX0u8t
h+/PmhWRAE9MM9OObyFetoWGDP3ee2viM+/FmQPLu+Op3V86IRzQq98XjYvyXBSw
7b3pqdUlrUU/f+uCE2LwW8hSQQrLfwQhKdh3b2HZAck/mndUFYLJ/uKQmNzlKfx+
LQxb/f33rPR4FSZjyJDFqlq3bT1vO1lumyHv43PRtCy9vtU7T/kExf7mv7MFmlJl
HPz4IP88KyvGweERPMuj6kv9iIQOSyYYltmqcBuQfVKtkjJc4o5W1FDykOwAAzM/
ml0yvjmiXPaLrK7t36ArsvL2r/xhSn0fYOm3Hlcnj1cIYCBCasKzGU7m15CxsqZ4
0BuuRwiPHOA047g7v+tMsx55343IMAxoFNiR2PVUayH0gUuy5metD8LiEPj2XrRb
/6aBNNA0BaHzRqCTPA5ee3Hi8Jq8jrBzH4pNoXfSk4z9+mLFHDpPwSCodanACshI
L8aNP0uzvSm9kchaLIIFl2gESF7Oxd8oOiu3/lk7e9yYVvWd+4NIL60eyF7CAlog
mVV8w0mxJBbi8yGbV8TovQR182aTVHSIBuje8vCYSvvO5yFa1c+cygVJXpnKfq/D
xCm0SALL3Isq8uRGv7iqXAiw+3QhR9ICW3NFUcNvV/7uVqp/DgH0JRMRwls1DNfp
VElNutjKmmX8mwb5nMrM5OXGYlIy05TyRN8X2i0wdaSJYpNtzO8CqXRK2TInm4UO
V1P4xdemLlG/IOkyPYeWps3h+L09YWorbKj9MsGCCZ6vwiYPDsNAzJvg7abHKkTO
ERGXFNgNyrXpR9a71CZmuVRgD31MdHWDY1ClEk5ypgBGmmXh0dKT3JlH61YzdPk8
Sq7G8qQ9fEIVpyBLC0fRW/8rYD5+pI1sPVoqUZ1j/XoeYsm1wPMW/68U7tpsPLVd
PPfDjcmW+zXZYcG8Eg/SyiG8syV3eAnFqS5bC3//ha1SZH5fDPNaj95PfoXkTyCC
V011zx+rAqRJBal0itqtAn6xwvvJqDsIrmRr1vmPTm8dTlce2flMA2IcV7btAI76
6XAN2xPV2405ZbBsgPs0FUDC8y0O4JbrXzKYWImuLU/IStWBvpo5/U+uiZIlTAW9
mrEICoIbf/QlR33iKYGzOzMmPkxvtLZRumZnbfuHR1+806ccTvqfJZ5cmHqUHUNC
KlM7MYSKxf7S9/kzsSwME4aDKMTQjwLKz82Q+XJDdDcDjwSQsKoIgVikugJk6PvE
1xtr5LShOHvEVNatPJK4Pa78bjFUJygdZTsGqa0dPwwXc1o7eHUQJaJ0vn/Ix12i
C3aNrKYJP17VCo6S28dDH8zyrrzJwmNa5/VVhGs84jR0ixLe27OXpwBlaS/4RaHV
zz0MlWZOBicPTGMZPrxBGuNo5gbbsUFVk20LKmPyfPY+Tqs/JVY9tXcYKfjmwolx
nZ6NJsDdzidhrfqWvZroVjRGLMqVZfEbyKoYvjlCWXbtrCrrupPVFLKZOh/mQKXo
exAYREIIove/VYeCUQ0iqfNRDvNK+XqDR9iLhYd2zgdyoj5airi+dBPArmEOPxzD
DbVppPtJ2r8tjygXzHRGSB04M1Obr4wFAFu2ZrLUJj6i7fjRFuCwQqhDWkKKOl/X
iFuFqVHmSsYbVC3fo7t0c53zryz3ar99NqGIzOD0+c7PWxv3eJvFiJFWy2HCd7Fa
9x65cjwNLYY760Tk0cFtL5tiPvvwKYV9aTWJsNR1/KhIymZySRjaj0UGmfu7WRnz
0RRb57uVrDB/Tx1cfvUkHVKXNbqYoMiEc4yPgXGhwUse1Go06QOMZnzJ+buG8Vo1
89VX91WUuGBV8UbMTSXFKNTNHmjdDAnSsI4PZXiegJ7PvAQ/HNrn9odtoIX1i2vL
UZ4PYCORNTPURpb2ca60eADR7gXJKoba9wHYFkrMdP0zzCn/Jhe9BdQdkgVc3VfW
sukMbA88HpaqRfQ/GTD5jHmeofrqciIz3xCmsqsKdeNCUC5Ane7w0lhmS3f2N4Sl
1PCsTefOTi2lmNsJh6vsstHOb5ao5IE7KZwM13eef22VppxGINIytcW1/zGDD70V
XL829iOrrqwGxq3n44+bwKxe1Hg3N+c8gCK2RUclUrnAottXVvkOJFYV6wwxgTFl
zymqkm1AWLbo/HMWSuZ4wWpaxqzKTHUyVDj6z38f81kX4oqJlxJGTuEjikiJu7nC
PNYEdmbKADbsQ1pCaT9s6bb43oh6oy143db5Z/EOqNuS6AKPzHclRX+rZpguCXGh
tm9ySfmH5fRF9Lxb6ugeiFZFKfVpr2ByUm8LmNQVM7PpG9M1r4lEU1n8E/Yp5Acy
wZ3qdLcA1GPcNKhlkCcOM+7sZC7B4ocJzVA1AUQnUg3paTmvFht3q6+4dNns03tS
3QY7wqB/U3hJZ1mWdIOxQFmZhbLfpkkklwsdbkRknrr2UaUr1oiwNREAcI1T7FUc
A7IIhSL1+NGhIdqxOGaPHQnXFTvXctGbz6/TrM3AUQYV8bj0BS8Pt+obu34sGIGO
QyGmyOb0kNiH6WgEaeitWxDDt72f57Kc3r0w4hOLyXBEPM3pHhB9ZcZg1jB6lC+B
K8/Wmn2sQFL1M0YE/FHP1MnyLeyVJtQ0u729kiJMHaPrib1cqAjYXgbpOAYcFoCs
k9w3264JE2kcmaZArregeaI2QdcBAR8np6Uxbnv0oBCOrZhBxjKqNlettVSOQ76S
M3OLkqqAtgXJanlPAsAuNfzkyIEVCuvdFwHaXOqtekOwZY+9reKLm8480gM4tXf7
5KK0uGhk8CUpvrG2ycrd1Rc8QD9Wk7b4u8qD2WuNKhRLOk2OzT9/ccH5YL/710iL
pFMezOlNdBws5bFX8y89gi85t5J2791kb8JhpTavqof3tgeEG2mDvNPjyaYr7X3s
zt7a/ilchlR8XMyG2TbyxATdqKP9ClKgemD7lfYCgwsxw4oxQ6GWSWC++xdN78/a
LvtUTjg54/fLaKpfmEgCjE0LkPon68aHJZdvTTPxj1kqTuBnvnqmNa0+wvcXyNOh
oum85Nf6KmlUiFpj2VpEzdH01zZ6DpdUVgOsI0Vt+pjWh5GAmrsexxh4RtsKzq/F
OOyCedjB8lw4Dv+LPU64iwRGe0rrBZ6VS8Z8YeDOQ/8V54j85pc/rkUmbjV76Mn5
LlGy2FYRzGvsMxLUIe7rahDVYoxaA/sRmQ3B1RLVbviL0gJ7hLwk779yifVlWl7T
gXAPZbDFt4rOTuUlTQ6faLK/52KEXvhyNRNaS9d1h/o7j9V4PCNCsZoIJJk+0mrs
dQmDRdud5cYOhKP8NACTrisWFzsX6GhV4GwPZPibMPYJWpqQC/NodFNmgdIXfj8M
PGtw4JcB1lJ1w2eriT5ceaP/i8+XEoyXEQknvrBp/KuEUIrYsVRRmevFSL7jS6gx
SI1uva5Obykl+HScIn1pcy6GxuAj7vU7JXgdE6/sAJQSr44um6AgEy/Lf/tCkNes
s6wm6C/KJ05AFyFs4G8K8O1opC9xZ/9AqNT3B3b1sCi94ishlFEB3elTHb2uRFYv
VKN4alaMueeIfxIezIb33uCMHIjFOkMadBNNGu2FzIuhhGHPeA5SkSxHP7+tt/3B
Nrn+/EG5hwg20eoglN5qZSMnQ4ld6GcLXDnQ6Vsgo3mX+NaN91o46QYbYjcNl/T4
04Pvl2oQleglesElfYosklhX38Uj4MpVRUlOShYaKgodGovC7vnNNm821ed3hQMa
8mv0kNqQN0OOTVHzD+UssG9AYq8gH1hwzWEkQmNZdf4efGBU0Ibdv43ZaljCh+Lz
19/c2SKHho4MW4wVOrRtD8sQAjP4ZMoHg8Y/5xq9XEHaqSBDwwSQcIEKYpH5QxwP
GLB32s+OKG1GTHTTMkGlvz6zjX0HI4eeH3/3yEaWgBkX2P/FcgbfbJNwEnSD4Vc8
IJDGBhoAWHLU5pef03QyJwq11kdXbTM+actshfyVLD4YJyvnZa8VkRyp/BPHFN6f
QdBHEwktQrUckEP+UdAXc0BCMnS7fiArC0Ro3LqFrF5JmQnuak6QmEWCqSyTPis4
n7YFWLBQzh45IF8VcMYKJkzTaYZY232aXWyOFaZAM63l6QpzXPY7WumTVI0v2aH4
NLnQGWssVMgQfBmMWGW5QKiSkiZUpsBjiA2Fh+4osOZ89yi5bm0fEb6sVAsy+Fo4
KY001x565lg+M1iwuP0iNGqE8FiiPEn9hG0MPUTr50uoxvugpHe+JR4XPQLqoz/k
yfgCGVjhByAJGQmgFs0VAP1OSs6VeVWcuXMR1JNuzojBcaxZW/r4qOBUFlJRAIS4
KGLvjgvMsV5yAq7Ceu0WQ9apnQ6TF7M/8wFZAbPxzpMzUideNtDaXelTtu9QmU/s
zmiZzwOTh4fUL/EZJC0qy7t+pwdpC4btb8XqoSeOI78QG/JyEmOwOoLz1OC5KXj1
aK9DrHbpbbqyeRW69BsbTBznVd9QsV+kxS5vCyeV1m6YqZ/iS9OdRYq7YIbe/rKo
SpbjXGPHKXuvxkqA5zFQV1GVOsKdfesWpVBBYHOB5+fUyc1yYimMrHjICfPCMKQr
19amE5iQEXyxYE0lVj8h2L9gQhrTlzclhIGNZfz4Cc5wH1N3vW4YBxbnzNxDXlnH
m0Gs8M/8LGH2ffZdHv+nwFpHLpWCUmxU2B9WkCCHsOjoKJUyPO7EnKmExQ+zqP5L
cZagh/QQtChfJ5k/VnTEf5rhjdPftDgAuUpPZhFNo4egvqKnD7ejvt+VITkxKgFo
L+cPmQSZHLqHSqfBVG98KVTBx8qQhz3BA/oQEKQXsNlsmbsvvKdsjvraSf8XzrIo
k66GeS8yDLy82WDkxNwVWcHiIia0OcRyXs8a0f4/Koxm/TbBGIwOgjrCcnee4xk7
6fGl7Pb55TwA5AOFJuP15g5AGg3eoYK//n8XdFyuxxJXHpFltyBsmRNdZDoaIHaL
jhIMYc4gl5MYupNHbf+bDIBsv70YUilhSmZZv/kbcAN3QkZhtTFZXPj3+ja6PaYH
bBJXj1WRo9Yz5s2uRqhXmD+hhOgjuYuWiP+8deLG35qGeMLULER3hvtq83iX/TPu
6DsebU37gpUyGSYCYEalRmbpysQ7ViATl+qdeR6CII0COu/MmIUmTXDl31zYqkcq
hcdfpmScogTICdBYrdrSamHyqpOS5G0qRnd8bJA2Uzh38uW5Ppebepn9al+z42Lh
qcKzxCoh0B4y39jvCuETMDN80FOQ2KzYh3ipQw/bbJjRZfue9PuWU3tH/4aQI2fJ
YrnjRVWbqEkgG5sOOQ5MyzajJsXM9zppEO1hbMrtV7UFUXKPwsIw0WppoFppmDNd
hSKgeo+3KeN5ltDnAORVTJN3i2378vDcrEu0bZcJr239IsfERqqfc1TCVcPaSDT3
Aa6JIrIPZOUJHQbpsC3Kp19GG3BHKNm4JH9N/zsF/UTRd6k9HFplKFpqtsJSAIxA
rpPk6R+6Qf3YFAwoDo+X8kJsb3yNPjyv0DnIrni6yZwh4vt9MjcjZ9c6a67tjh/2
S0Gv2ewjUGYwrQd3eYXmS70JNtQnVcovyvDyRG+bN4Hluqju2C4QISRfATwOkDEL
WFfs2/ogiqWpuwHpSHOjQZQbYrelc7gQ5X44pma3gGztaBo6yRKb65vCMi8tatdF
oLI7PAPTlVX48wRzXdhxYwpnFTOlnpGxMmg58Dk3CNEYI2K4RQGn6O8jkERNf/3x
CipekFwxLqlRzsbmR0slz+TdgmH1HYvmG6+W3MsckHuwYR7FoTj6LLTwaXT/WOUd
Yb3Wc+SbQs0v8tvBXrPRPhhVwhLXtY1qNG/3S81KWq/0t9It2jnPt+g4qwieHi2i
qiby7Bvr0a8sFYfrH5h7KfUIYn+8zKf3ipXF//lNRv0uDj1VLdhPy0AMhSEUwx7v
iYRkoKVeh1vzN5tspQ24/g+/2EuAKawHoj6T595gRNqVrMfGmBoInxwnu55iMVQp
5EOlau8SV9Dv1t1gvtlIDKCiJ4JS1d739ZYzdr00WOXQaiOlmKGf6Jt3z8uZ+eQn
0/cCgP/u2hbGra1CPCnPKqvOYPlYuSai9zX7D6s8nPXVWZScBlXF5wcFYCv9uIgL
ntuEL4FM7j2ByBBKF7ZqVukDcDGZpb5Gd+YThyE2s1o8pnYJiW+EMoPt4PFekQ83
tlVq8UsPAVkhqE9D4GdA2E7qWNzaLKOdu29OZqbE317FkBPH8s56OGzCnU7r3Owc
cFTfkcX+Qkk5zLepKD/KnmjqUs/TokMFFxznlz/p2tPjG7qSv8w2NwDWrGeHenmF
Y4HC6OOaY9zwQs/O2vFOi8/BmlDggTsOigkP8z7KyFuVMeHSqmtj77O3Qw4D97QO
y7DyUjZbanjH1IkxczQ3xpUKRU5cQa8JLoiWNiCv3Xctm70ygsNW1q3lVefXSVnp
PNA6jWoU3PK09aUdKsFrvQTHVlfEdwbQzmZBWYqvTVdoDtS3MAZu6XXVW0Ng63zM
XesuRsdfUVQyHAHeDZqLD3aZrY9Cur88JJc/ZmXkl2GRs4N+ndppvIdBSItZDiTB
hInSHMSN51eT1XCn0ZSUUnFFLahKMpceTj4NwukSTP2ekfMqyRqR7m0RxFTyB+aW
/FrdSYr1nBcfmVeUQruEvExavII4co58f2SPaHNgsciTukwuQYnY4Y/Hq9rucClL
rLCQBfEfd9YZvM3St9SuUmd1qRS5LzFudaKUeu6IUwyij9XEfNS1p1NXNMEm74Kz
6wTBCLoLy30/qjyldjHbx9GWJS9AiE8LO8SQ71ozufuDjaetkSs61kYwcbCJOeQW
/ETtHfCFQVVBQKGiukrp9DYVt7nW3HA51x6sBDRdI/w44icdUHIrvXoX8JDUUcex
9wWrjiecvpjkjP12763Uz9Z/jdCWUWp11bcCn1lFp33XmqB/aldbblAFssMejywZ
yPxPvHCTuwyfgtUYrDJrCtma3YN/WvzBZIUZeC4mndEfbMtOWqSWeE5EQiMTYGy9
PwBsLlR7pvCtGt6ZFR2neW2T3YtOG6PCT4K/kjJ43ckL5zyHxVQW+zIaLvTafnZV
J2Iay+7lQxm5ndUHCasdcz9msCst7XOFknl/IngYVP3BRJiXI+C+6foEDcfOdCDk
59PzB2Euo8L9YIGL6+z2zq74dD6hzAItQtF/u2gHD+1j7foGlAAQXJbNXWzT8uX0
IbjW9zDhvGZGOla1HDW8emhu0QO02KlbtprrMNfEwSeMN/wgLg7zJLuNSY20Znub
VGWVBZ/CJRjWDbWFQM720Cfxz8Awdw9a7+Wb8UyMsmh4WfqNjFSYQ2J9+DDtWHP7
9aZicgT3z8r/HumzFOyze8aD1kigE0Yb4lVtQyyVyvpM+UctvpIO42qfOtO4YH52
eLs489RTygeqzEv6sVxwdqFHsMMPS6V78evDwHhhsUH2Up0IEA0xb/gTd9NdKofW
/5OrDCetfvV+GGXJCBx8X/3zU9kU7zf6psbZEE8EuheUJ9hy/CxROOwvDuT/P/02
Bs5gReEbg72LMYVCbConGoHgcX8Pl8ZQj8WcI9I/eWEblNTtgsXRs0WEt6uMwwkQ
FSltC579H3I6IrYWrbgzL2E3uqVyLzmqQqaRRtPnLQlzXJ05rnyKZrFJG94rBqoU
kAD4kzvKShRi1Gf6otEYQNCaOmuuQB5QhlNqbozIRgX3TcT9moRKlK4ccUrSm17V
n9K66Y/g2LAvXBqvEieZbxd74T2PNi53tV8U2bEC2J97txphf4XMU2Vis4Pj6sQE
GBBYBxLjR+E2NBdCXfsXpbEBKBCvlmi78v2wWcmjNWV7vqD+YoHuCPtuCnCFZfoA
yi1ws5p31aSs8GMncWlR0TNC+zrccCu5YdWLn25QFsX1qP/XvLdQKITTphOmVa89
shU1GVPpfm+kSdqUvAYaVeuLtfcj8oAWbnMdxAOHUfS5LawdEjf5+8Get+ul0UxZ
V+/iGjXfwAKd2CoyquoGg1GpdfP1yZdIoUzNd3OlH5l5EN/l3POXVkO3vE/nf2AE
GOQjC1b8akOzzAtQPkR3LN8RmEFdKalF6shcTZQwvTMfK5RE4yRECeHp1jKct+Br
ofcC0VnGwdGEFT/+UyNif9JTmPL45hChPJLFNUpenR+ZsPcrvtzwmlHwFiDgX6o8
GliPtzRVJbb3Go8WP2LzCIwphpjhXJLKaY9yTsmrfY1c7jgq6Ek6hj72e+2gKWHx
XZGSSAKM2VP4Kq9mjk5DhdtR0bJZ68oREUtvmEIKzqbL1/nz53nu+dlkSNb0lgWX
C1KMdgyIjPKaRnKnQnz9525t34WXX2uMFPjY7mnuk83n8Wx0SDhxadDM93pBWUkm
I8HNy4bfP80Vt+Uo+CmPk/D9WSP9JPMyKJslTypm/XueLPpycXyowMBbkV3cyM5p
cchmmdwu03yJq7mxikLIFHBkEKTIveFf1gGldmX5Le5d+BRww6pbj7yXJZ87R48I
qE2RDVzyPcdOpzqwqf1dJtR+PvYi9tHQitCb5gaZgQkcN4E5yY5Xx2efKrCvy6pe
x+Bfce9ay7n53LsgcSv+uDLsLzTQaabVtvx44SZlejchu5QEUcrjyOAjHpbpgmBB
dM5v55juxfuoMlAoBOmY2ROIjJIpX2uX3+3Cda4MdKBfu1G/05A9zgKZwv16Oa5X
QSZ9/Rkz4CP1uYzopuaQ5jnfj2AmWmFZx8ouUU1pcOCrzYRFg2oIe54q1eeKa506
sY3wcVD/cuNE6vVP0v1auGz2WWREvTaMIHQMjrX254vnnMSMGqO0J94NTJYrvIyt
hsWo58W9qpqUnzgtp+0w+U32Q489cNU6UXuoi0Ym3ypS6hX0i75HOi6smBNEf4I/
aUvssBHQcykxtMYfbKZs8Yfm27jZQlFHxn0FIS2R3KcJWMNEP2FGZxoEVOpY8HOb
l4lvahvSj9rv/GZZS07ip9quALJM4YHXge8w+nTePSQ1VVSO0yhRc60zfEJKrap6
884IfkF01SwwC7vyis3lxd5uE8AwWkDfG32PoOEaTQ5sPQPcNHLgIYQcikQ8JG/9
i/AcujQngk9gSOXuWVfyQY6YVr6K5XOcRgYbEDittLfBbVWgd+1k/5XYek225Rja
JZJktbMvlJAnkYEHQubFZVGbBwzeylzy4F003EakGXhYVCfTaBxkvVDZKFi7Zgka
YgP/oJpw4fk8/EvCv2cAhWOZtgAidaMIR+LiJ09C9/BA7dBphrVLoRZenVPoYj5h
RjC0jQqmj20fAQgaUC0w5T+tvRWyWrdo+qQf4yuFxC/iQ82oKD9Gm0vXozyKGb37
N0UIIw+nVc+aBdR3zuvW8TEZX+0WEKg2Z8sYlNzQysg7TOcuUNMEzvY6DnllNo5+
Tq4SoKw6DlfPOI3nDjyEWDFNXon+czwulWcxE1zKJo0SYz7dfapX9kXRdjVc0wAY
k7v+3S0N0WY7H1weTEBFSvESw+l278Hn62qE0AmR48UxcSWCDOzW0Rv+53vuc5cX
/Mtee/cArvT3PREkYs8Eq7fzpwQYkBWUa2/1rUKbt0QaciUnjxAerjW907sTigYq
/0jclC/WnfvwtNfqQ5cvw5A2BCsOm/Do/hKf+PILOJE1zkN2EFXsbgZ/rNMW20Uv
nUVOU2yViBJkuzl24O0ILE6nVXD0KMVcltXa79OOwIYsF2TYLstbuH+UM4JiWaRu
0sb55IKco4qEzRW8bKfMvkCaoUNRPTPGMpQVXRXPym+Rg6CDkXrZLfcUlCl153Jf
Gw4W+prOc16dBm1/VKNoRfr+FnUvCajJyH+0ExijM+qU6DMNDBkeZgxAKAiSMXY7
HDd8PJ6P95fDUklmz2ygM7V3F6/iFKNmHDPEwLoX9arFOPYXLlzzW5N8itEKzT6c
Qbxc0PpmR+DxZSTwxoSR464m4XSG4N87XO1Eci4uiFJ8PAOkj2kXeEs06WG+vYSp
+dUkQbj0GvLB7cD3Ra5zZ4pNymPBWYmlPp6BsDNv1dGqLnkTwxt2d+XpEnmFrJvI
rXpNHJJIaXfhgsVlFejY/oUujWMIKLayMyjHWVzowwBFlC8EYH/ljr5AnxKPyAvA
AHAowjdQXvywhYEypoSguqLl4wWhMWJOk7QJ4+FCs13UZSC1mkZeET020RU1UEJa
XwfKwnILcg3s+HqRdMUyKk5seUkH8SwR+tgpQZrt0cjCRJGP2s4lX14/KP1ttmeg
29KhU554UVGU+G1ITRZPBr0Lh0D/ed7Cko/WfWK2lIvOwuOlbsujo6Be/poCV7zN
6G2uHJFZiK+c0kwKnrCiLolCRXcQOzZLVox+HWw8EkKf+p+TvoKISL28jeGvvQKT
yZnYFqE7c4aYK7Q2XHgNLenzkHU1QgJ5dXnnT+87itgztmmbqZcDyFiiATO6Rrpr
H/WPAqkyem7Q+LvWTXKJ+39cWeGPpBxgAEtkXt3uzyuRdI3jnxWTyXD3SVm/VEhC
161852FgvU9g86I8i/n9zeRZoB3SdVqmGXDjfiWvZJtL+PgzoNC2dL5Iqe+8X7cG
LqJMkCi8eyNw5bujnBXQYULu6YJfFFTTlLTXI9zzVG8yBdjj0MUxAESmI5H69cBJ
AOtBH6JLx6xaztQMxopTjoBua+PkpHKNnNCMGcSU2s1j/zTkcBbpJD1GDLmrWa33
apAaoP9PwhfUBOH7CYI+UQPsG7+kzBWKdbKMpWuFHGxavPw5fmQJY392Bd8Bqijv
tyRvNSDROmajK+thLHvW5GQfVbLLsJmYWzrmon9XKMFhdjHQXKXPJZQoIxppxOHN
26GC5sHnef9DH51ofyLD9CURFaK/VEB8nbGyBiQ2lWzweyJcChnUpdRV3rpSToA3
2GUOQsSAg2hC7q8QlxD/ZT3J/p17Ky2ByRFeMT+f18OtqUWvm8UwG+biKH19ZzoE
4lGp6/Jz0POG2sVQ4bsHI7i2LzF/wr6FdJ/IGWNq7oG+IYcZqEk4kHypgcoAT2xE
P3OwrrzwEZWmLHEd06+MfGh+JcIAQFkgg/4a+/s4ZzKv4YPwGhJzG2TF8kitw7Hd
UVPPLFX1blhlkKFYmLpIf+9gcA26YSa8zoMhFfMQoKH41u8NSzaqsgOdmy3G3mvE
Cg2/3pK6glsfJbUYsaLQ8+nd2ocwpfeeYESDtOcCEubifLpqFAaLPz62S0NZ6kQ0
ie9R1tgP6AHEafr2iM5I5Fsg9mhJQf5eUENA1Jd0brisQkysHF4KbVoxoK8E4QQe
LM26lNFGXZ6DkGyfgdAGtZJwzQIo9GJg8UiTG8hqNj0F6sXMb3SMSIBljGQKdX3x
QR8Zb6gDBWPdMB9BvbrQ45jNvbGUd99dPd1aYJhruqVfPO3pbMgFEcBTDjf4xCet
w7cq5QDccLueKlAdl4iwPyQpLvJ7GInGKrUBOmc2q6gAx1oYBaD3e0xGFj0mzJ/V
GG6s6l/x4XQkfbbZYAj9yt+eFE/OGvQGHQMm05cKSUMMRFkeqdgZ0OJ4hzsTJWlz
kFn0/Y88JW2wv7gzq1ZK41QLgfY6/4IN5aUWnZVaFpKfUZwjQWw7OfuzPa3bNmx6
hQ9jz6DhHPOjvjXkdGt/JaKuq20FmRWjx9EuU9Pg0KIxdtaJL0DrkVvAwaqXy7or
v4Q0X3YMM9hdTioJS2BihkSm9QZ6zVzZW9D/5C5a+m3bpJNQZbR1pY6brFJWeFdY
pewExW9gR42m58b/f7S+ix3yeCMkQuHnezkTf+RJTMKJxPykdrGzTZIx1qIeXmrC
mXXp6B9pXdHTyEB5lRgtd6xWHrRVZTGGLpDugfto7zA5p4UHQDEK3PLnb/Ni2c52
jF7x87Uy5Dz8k0jWc9FduHchxCwv90O2Gz1SoRzLyGOIvSA04fxuMR+KnwwHfrhR
QIZ6prycdZKMt+CWybDmoL9COx4iIfbUHoU7ixDZKlQgLYPNfcN8c2xoYOXRtJeq
pLkZY9IsJSYwAeaK4T6k3p2UF95kOpMlnUOj1st9YuprGSv0kAJjF00dzNVj0Ywg
FXGw7n7C1wYDv3L7+MrSDtfibzFMGMzwLrUvpEiD3WLvzZ1DgT1ASHNu99LGpXVl
mGoTWRV+Pe+mxWHm4neg1y4YPf3q3lRGpBnz9/bnFBvw0U0283rqAgNh+I2q++jh
h8alkCxU2OezuQqE8roLVHegaMgBncOLc4PCliFuFIhz+zusn7tH1i5BA9CurUbR
4UdrpmT5KUFZl86XvK3+oiIhLgL3pEEa4XoX53ZJZ1ug5+0K/Lt69i/w9+ag2JA2
/vFIPl944oPjZt1nJ8tXYgc4LA+P0PxK3veDtoPmFoTn+CaYhIwdi5njtjnYKrrV
d5AAz9wWlP0jwzkTRBVronv0oZVbom00weFb14/1lPGy6K3jacxg1eQCjPKP31iR
ifYbSp/jIcovXgY5/3A0Aw==
`protect end_protected