`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzaUNycXRd5GOKUc4xUgAG8XAQsV33wgDyZjB5GGS3nm4
FROsF4asUyAg5o4dygukmoZYyfcgD6g/g1GobTDFp3KkUvIjHGb1dlNNOd3Pt9GC
InH0fcC+9mr9LVV5pwlzxYHEgpveWKJPx6Iw61NvkxyHgKJyCKA/AoSIXKn+78Yk
ihBi9IWduk6ncBxHU9eQZvoMm/5glavkxnO4Nro3aD4cVyR1B3+LD+2mo0JiRji+
6wTd9UOk5g71JPrymM2stJ4n8NExHZNEf2lDvJtgwlXDm1KBdIEsOGqcZtl6ObGz
bFBhSgO6tARuC5tzCrj4IAPeU8erwltjMcAoIkhrSpSGl57Y8e0com6gFyrGscGR
tVWsn161EeHjY3vtmZuHyb5jz74Dn2Mg903ikn2LANMj8sabA/IFLI+/xZlmwuTW
Wy7wOrVKfY9aJ0XQaT/FbjGyB5PnItABycYg1PxFDoKXlqLMHl7N03Jv+ks6Tt9A
346rjDdR0yCmjTSxGnE2R87JoPuzRhkwpBhqivBLtSTDoPKARNekqfG0YHohae8O
0tZW3oMRtY0IXccW2xDVMBObaizsfu3xtIhS/dDOqwFuOHCBMHPMqA28EsLY8Y3p
Zj8Wp6w8vrFZj7W7Pi6iZKNgx5GBROeBR784pRrAqfaj5wDSHLSg35YdXazBqLO4
TH3gFn86bRkGNVlenljzqkNlIyY7kc838GWx9PG4zeigSm4czZ9TWxG0WDNSC1dr
He4FF+8yJhgQxlpKH4VimwY1ccJoibFkjgWoaY9+59D3OWQRXlwbmwMh+ObpZX/s
LqaM2Tx2bm2jJLV3vw916zutdd5BtfmkPA6DNjzQIVbeI6z0cveudkZdGhbsp2+m
+sjOC05vmaztCKQ/iNk7ZAGYcrcsyB08B4YZpsDD6guATM6rHb1P0EAuQ4B80kgz
It1UsADRIowxn4LoqGr6T7MID9Xc2Pp5NoPRfVVE8/0J2tvn2g0nmm07vNQgMjV3
hP+7uJu+l6zROo/8p0X7i7lnPt3dUqmzXoY6j+HLfaiBhD1oEIT96854Y5Xev3eZ
gcLO5HVvulG8z/BsDPfxbyCEqWg0gUuqJWtNJkcMzPOdI4ZXzHX+F0hkvhkkGApF
NS1mQtsCq3mdNHaT/6y5jANzJ1Y69uJF+37LZota/EKA0MJCRqgvcRlWkQdIDvfD
ScW72095z1I/rEJFRSMzlvtrLWYyz+lUTxAQnKuaQk5rxPQlLuxrezlpOK5Zr/49
nzvILwrkvxJYQLTIqDihy6siQqtjzh3gnRsatq2teOkYObKhU2cPkI/HINzUlFLk
Ukl/rrkGJeMhKz1S3PThSsNGqzlsvVHRZ2FeGfwTCDte0t5AwXVLmTIa8PoXYodw
lvjQQlPin4NnPmJUFBdmjFyT59uTzSixYf2FrH6CgT6TNUB3ryTXOixDotRv8G/H
N56B9iaF8PuMHCFtbWXvH957CZtyCwVGjAFT5SKe3EG7pNnGZA4SJhl5tg9VOU74
UVXPm2BHr7QJEWlBZegbyfecPZ5RdiyxnBVslfhiPqcVH4NVddrEOqu6FptTjHeo
k6biNZM5mjuuuLFVyUa2fgy3ZTJsjCE0qdiXfl9bPUG2YQ061i+8T7r3y7z7xkls
+b0QGUnU52vZxuI5dTA4+cFa8q9AE0mtypi+8nlUoFjcbBQK7xmLoqp7RhcebfGe
7jlgYZmkxIDf5hamKglBSr8aI5wrtcgFy22iQydChndYTSOgue9B2dtXcQMzHj0I
TZZImjkhdjxQbPkRuT8KEc9zv8ktpbIJH1tA+jz9neb4s7cOuxBGSQ80RUTZU0T/
WN9I7LRM3yY7UwAj2gmSam4nIWuO2/ZZLrycaj+Mjv6hOvubAO+iPUtKIswmE2r9
XVxvDcHr1KajSJKFQ77vFnpsDXIGmkNVlGImZbWRaMszCEctdh98iumf0GD7hong
5Cw0T4AUHhe31Lp7fRaUkCTpCLGxGp04UbN9tiWxfGFl2gnu5xYJkzja4uebqnTn
R5hOTWVFWEVlHpVIu1dL23IWm+zNRUYo+YMRfLq50WToHijJZcOnQOwiF/PMoAzG
JnQwMOrpoEiWnOVBlIJeqaPdWaqauy2007aLbc9Mdjbt0MdM1hG8ArIgV6QuZhq+
htD/Lb+v/t9g79puYVs2FLlHDg42hlzbbOdwTw/7KJblbBYcTlyHd5ZXxVDHaYPb
RlDZNapwr5KYmUYLEgbNUAzuDjEEGcISH0c6QdpSyWLsAPjpEW1QCsaBsWUB4j9W
F4VHMqN+Ak9ddDj2SygCF7Dt2X3zKHYVDr0QZh48rJ+dg2VkbyF/KDfaebMbWw/D
htWuX4YTg2A8+3p+ghVG8u898HkUang2xb3SuVsOOmUMmJrhIdtNwtq7j8klo8fj
N7pm7thUeddxBp4ufQy5LFTihXp7nc86kwlpPOXzhZIPe04kzxO8+7zCCbdsbxX9
vxlg6k/xgwpjzmtTeka6Eo3wjRA14RDTfzZ0BccRkEWFxLgKlYciimy/LVF2+ZEl
uRgQzCGu+79V8FUMbbNrlIC4RgeL2JJyT6SQjPwZxThlseXry/vuARmC6oc0o/58
08HNlH+hF4lAt+YbKe6qL6YQwhljA2jswoa/byQKh/3626ojffTKRfcv7Josgg9l
qjDOZeOmz+xA1CvyBettS7RnpL5ZaUhDWyYnpbd/XEmnC80BGz/5b+1yQzblq40p
kbPbS7CcAXK0SGdvbN4jcsQzyZ2sdoEhgCUtEwxTnQwQFRosi2YgnzEorZPtPj4U
rVhBzvkV3JiZh3tYzOyvQPxnus43zZtRTIjr5JLYi2voGmsHnZpETTRDhNeBXSTd
qnHmtUVdkvJC3QfN4hv/dtZRh1D6kKHQdt6Nhl6o9csmWg2b9TvEKCAjmVqotfFV
YqPTVEgsp3Mkc+DWzKz5RaeODdsvWWdck54yFsLZvJ8SreaRi5w3GiAjsVzwnswE
CkZUgWtzEcG2L91/F3QyIQ/SDxNL/Mh2lbTl8DUAYipIfTxs1zFeGayFBJyNH/El
1r4DW3HDlrcLngmleSZzYYPXoZwTPa76nHkHt7HokJmiUczhDeBPhqp8vqtpuBUY
07kJXpDPvOA1Y98/6SxEK2EgpOl0aJ1XEWshKirNePfN4matSbwQnUthB4yM/oIM
S7+AKEXTBAgqNqNTFJ761pFPhaYwh2HgZcEW2TwaAKAIYNWpU9dhIVqdLMz5H0Dd
qZIG3xbmVmyZ7wWrqZfnO4hoBqKxm+yetq/4JYQDZOYLaRk2RtGbtQVpq738P35F
mxH8jCcfzIqS2ZOz4rmnSuSTYIpxgDp0CaYewHD2H/1DM1mx8JpDeNwelwSqSslM
iPgc9wkwjoDIEeUb8UG9beTfJFxJ8dEZ0dkKIfDL4EpRuI7QUeF8+x1DIevkN3p6
3qIzAfEevPABFQQha0E0RoPB7AlyiHj04d8OaI4D/6FcuCWa+hMxMeLgv9sq41Y+
nBlw7iR3YK+XZcnMQdVNvoqPT98RybbpYUP1LmlmpX+pFMvbBebkLgdREKCk/r9p
el6KOr1UCmju5dz3VjKW7YY1K1d5gZD5xF5Ps0nvCks3uTk1kh6fS+c9hldh40Yr
lCKC0mHHIfSIBBU81yz/GLAJITznwWa3EVrqUpelRPa7EVRrtyT9bsmtu6UBQP0A
8j0A6z89CWKVT0mhzuLv06V4/xct8BNoInpsr6VnDvBIMwOZkOwozo8/ggOe77rU
9JPsY93lS6MK644nTpn5nb660YUElDu47OQCgxkLxvImsxZ9fv3vSTtBmsgy4lXr
qSViemy9GsDjomJ3WLEYlGRkwK8YcihPQfouisVI5pbnqlWFjV6cariWtv/IrnD6
fCsGMocS9vfOrz+uFq31QiExlKJPxs0Xa83dmEIcDEdX4eZCFONf5AlDVoNa8bKp
FRVodg+D8iGKBCDT0jYxqWDBMsRQQyXk/cDWV+tRKHpnaIbXSnFp5D8hxT1S76Yt
W9VQxwmRRgyIQe5LhN3YFJ02mnoo0S6Z2lscg/oSDyi1qCCLKGYVUS7jlEHta9bp
VV/sZfaG+jg5mHsY4XZuFun1hgP9Yz/efm9VAPgFfauuBRosjolv7dI9tYWVaBPW
Y1qfAuqUbMD+Z5y2zHa+t0tEli4gHvNYnIL5oN7OpvRUUoROOAD2ItshkWtyRRGf
w5fVRdkzLFhf44PybWlXrO5vKetzY1Yh/agrHUXjmM9ZcA0YoJf8vlE2DDtfJauO
MB7IeowJiGyvq2/YZzXiFTOYEEaJw4c8VlJQNgue2BG7IrNfto30ynSrUzQajP+Z
tfHZ8OmlQuwKTFAOIMqo1TtJWJZetOe6Z7ykbUS2edSD3WQn1xV7ppxbMbgqHTka
pUmrb+BNmdKgZ4YF88TAswH8fwrqdQ9pZDe/BCBtqZu2Dpy0m7116RBfN6U0yukb
CTXEhg4NQq6fMGvofaFVDMEOOMdou3zp4hom/ZycKz1s/m+ryKjfqmL6wmhIVgJj
lqflmz42WcwHDwrMjmnF6v3HGKUJICh9rEvERf9ttfqo4ddgCAuhipY4+c0+FwEV
S1/He77QZ35MYlPdutM0VfzwFZx45k0JFrQcblCkuaFQ2X5z9Lk6+GzPVmQjhJAd
xLSAC7hX8hxc2cxbar8zb/ZVZD++/d7+mkxGG+CwbPjUAdjy2hK9Q1EjFbphg/mN
RwxRoW1GzC3PtwwoK9VkoIX3va1hI1GFNbZynbaOcEpdVIXIeNDjwqBFxI6QXweE
O0PErU1y6AMVngUGKcxK5kh7lCyeswOJPRN93ug/m8+uIKqd5le34IwHWSv1LBOn
geptKbuk/AlLWXxY23z1nkRbVbJXlnwogW8ujmRIlIQ2y/SMo5DwKq022xX0wSDF
uXCqRMf+lfcD6aw8NcTw3OOUP7t5/KwqbAhbwE2YGQOUnUsregxXVnKE1MyEZ6RF
78zm0RlMiLKLJZYEcRVITgbDLk+wXHKuNQieDy7XefqQQOTd4Dq+W+TCPBRFMDQq
mWrH+FHYoWJr4rVLYdznjmMjBb/nhMBMPyeANgxm5FiFOh/5pwMd+nt960I8Pyeo
kVtHcSu1T0AkG3MAJ1Xwxt7htKr31L2+KPFqWkPR21BH/K13AYCiQPNioQz9Nkyu
rbnKQjxATxVaio6A2nreFgRkSyd31QpoSDvgk5YJv3J0HOaDb1zvYvNdjOIJfKdp
frbitVyje2txWqye2cuC6InZAThv8qa+F1/bOKzqtU28RHDVZshdE8LNPtFr7tMO
4JkGkwhC5okw3DvYpX7PQTpqUJ+W5Mxt6z4uqeqIDhUGHobDPfE7jop8ciBehdko
QFj3bQs1OpJsxjt6Qxu7vnTgBOfHK0TZ5z8/YpmAT2Xi8myuBk9Nze/QGDeaejhR
d5+SKetDJIzofJPM+IJ0MJNDT3u9+NeBEtT7CMQbBQXs3nia08Jk0ng65EQP77BP
Erio8rXt1h/TXQGkE3G8brDuwRAy208Jg33Fl0z2eAwGgpmCrUXTrvKgymRaBGBV
EqunL0Tl+pI0VulqcinVtZYEJV0kp+TGK6u6fUVIetADYIHRvm8HBK597yWLBx3k
16vpUMmK3WnfrsWat/1l8mh0mUf+j66TQV3+qbYMCbKJJjPhYlou+A5H4gvusdGv
2gEzFlDjn7cZU4xzUII8/BNLKCIusMIooojo/FD4/hqzo0gTsduXA25qTJfOdzOX
nBJexNCRC5/0GpN5eFN3obvxWRILhsDtDszs1G9GEHumDTwViZdPDebD/esCkjrN
G2+BwF2NEAtYuws0b8bkmW/tz3MIW+2nUdMpIs5A/hvXzBNBZKh8X2ObwSy7KN99
uUWA9Q/rU0h5e/UOFh4J6aPbaAFo7pM3vlsGD8uS0aVx7komnPadKaYEeiAYr+dV
5xeQJ7AN4ks7hbX8gQLROnwwPss8gsZYYi6ecBfsq9PvupMZFgoNQU9unNECO1ko
77z5XliZvYcQe2HTzeJmVWDgovb7c6zvu6Vk/Filmp+WsauhWBj7GIiS8LuNPPFn
NtZDYLRite3nJGaye/705srdbnc3Cm+DpbbmiPhsVo6XotaKBS4KncXjjALFDp7d
8wIfg8DC4OJIsIwp4AI/BP9kdEffL12sBSUo15an6hZfJzM9OY7kE/6whVygCDBi
k4ghUvyoMY41PoMRx3Ge4EGSwNXGHDzNTUxQ0CLcK5OVY7jwWrzQw3f2FcTNpPR2
LdBZ3g82958IF53MHK5GMvRpIwj28LtOP7KRbWsclM1hAyIgrhl4LtLaafnAk91M
NcO2xBRieMDRlefhnn0MceLTdR/BBRK5dU9Wfz/a0NRPzYakgYVbQ4/M+MDK5cac
YLq/zxWPK/RZuAOqBU1OOzqpxUDRKhqeTgtZtKWBPgB8m/7ke7X7oVzODmXWZmA5
rX+ZeQabgUUMg84Mk7XQAlxDj96d/VYmf8o5dhi4jC5sVrSlFwsf4TELotNSMget
u0P3oVbjR/GtXtnIiAAB0xxB+/UYBgHY1XOLeBgEeEKnKW2tEhPgHPaWRKZer5KF
FpWCrF6+Qe/lsPBtLxJfhCUUnb2PoXQvTMNO9JwILrtzD+JK24xCuhr139ezR7o2
xZMV7t0VlvAerWwVJt06AIpNT2Tu+25QoWtMJXWolIGsEDl5GXAY+6m8/WrycVy+
U3OFf+c2iqRTztvvGry0Papr0GSxPvWf2Amn9r3puPk2Vmr7wF6fbbQCcruFyCQX
7BbPmveIzwAcZNHi8CvhrlMzLN4DSiocVLtSHJ+2t/xi4yhMqHpOCwApNQKyuNie
OWg+5s+FpQCz5APux4ocikvYU3s+fQSwPAonyvKZ6KGpR6IpRwYK/U8wZgob58DZ
GzVp9F7sBRyVkDY6h6SRMVtMaj9VrE0F0Xwic86iR11/4Xxbx1FcDa62J8uXQGCu
/kHjUZohss9gVLHnHyInd+66EXImWi55iYpYtqPmdLsMfRNBBxmsfPTEYMeTTFy6
0Yoq/9MLMms8H3atGNLF6vs0HD+Oao0+BwnkmbdJA4VDi4EDjJO/cVBgoR0iAaWT
zz2NexW3BH15oeMJVPh9R38l3dgekVXLIBKMU+Fa7gr+eR4MGn/q6+1lqW93Pnis
5dI8MUS9JWObsVmb23McRWdiNSGiIBms6yZL2GjaE+rPXIYWpytq4lDD+GnGGBfL
tzZd0R6tLFzRfga1UbkrpSnmHV2Y3zUtoX5WxK1/0bnQ1ekPkUvtS8S6sjhTWZCn
o+n4W07KsD01lQ2wRXMLlzzOP60u/n9oz31B6vFBtn6LRTNb1ljb49Zf6OreqLn/
PspkhefQDSGSs4oW2cHWN0l0WCf7GoUeNVSsVvZuFsvQNHglQ5gJyG6UQv9xRVoH
I8ujjydOwfkM1HyXo8Jmlc4HagBF+D6t5Jn3M2KYA/RIT3ye66cZ1f2rtIYeUmLc
Sm+tCcVzTn3v2USlnM543QXq8gfxMSRn9pSEuqtFqUWbArDMEE+7Xnd3yBUIAlM9
42oz91sJf8U4z6SpP47iNZPkPFaZOtZwqCzhqHvvLz0oMOYsvzEBUBSEyFPYmQ+v
BJ1WmeTprcstHmkQighJaGTqRCEvy+qo4zZfZ73wbaofapjXqT8IfdFaLbNrahLz
+SWMtMcKy0FQF4oBU72mhxfXVA4EK2q8j2cfFRm9KzOTwVGqAEQ4iyphzn4ZJiYz
t+T/z9XSC1ABZafYMfsZi2Ih88JzGpAd04IENM9aN6JQU8VrxH7d6yoWCx5VhyBL
NfeRSfKpcA4lSq1q5JNFLRwCBKtECNCUtQh0cJHccKChSB7yxpHnruEiBzJrOzql
Ej06AXgamrN4k6D+pkpEJ/Iu2skatiCfQl5LAqkn5UXwh6BM0Y+lc9DZ5thUov1j
ZyYAs9TboVow/CVwMosnaz2CIQXiOlQDTfV8CK5hGmiyVxgJp/zcVxF+HZ9H+dII
sCU7gI+yiXx2uDrjyel2ZYFVLCA+M3bqy/UcF9imMmBmOePs1TUp8B68zK3/2Enp
8v9r+NZ9s/VNcGwDjEo5L/YmlA+6+qQe9Br9z376YWCAyp+8BXgHAAx+b3CPa78a
gaCQOWU62EHy3bDhS4h0vlESjAc2tsxO18jV2SpVvIW5HfIJBnjkmRuLB85OUhxQ
VyABdLC84k6CaHpDCCnHIbAaRGhyg73idHiWy2YFYQJnNpD1/EEg5S+GiOS49hAd
hxNcl+OLxLc9Nd8yIeFDWG2xiDbRXuSnVhhnjhVO2rkpKUIpMx+wJA+in0d0Epav
ob+QpaV0miYCZHy7BoYHeZLHoIBWy90R4P9p3Y4joeRa9LuQHLoHKxUy1Vjlutau
RQT1rVgVfVRQcuUudtcOk8DBpQc1j2RZnp8St0tToy40rMrgAZzk/VLo2+qIKG6s
lpRcSDg08TrPJc8RaWYnYRq9B9WnTsUV3kePezUSxT9cHH+LoZ7q1bxYruEFrpES
OeISgCThOuF6O9NHny/8OeCNuSRQQx1Skk3Gh0YHWRxvUkfs874rsDcFyZXUCXjs
uR4+p92Qy8YmOwlLWPxVchCCAGMHFcq1bptDQbR9pzTB1lth1CT4BtqQbzFSdkHV
b8sdJqfK9agKawE4JR3pLQTmYwry6Gq1xP6IHaj9Z/9OQ2qwsAGsf9CxS6FZNmSK
cQMyuoa3GW2JKbFTQnxCmn8UmiTFdv952Itx5CRpPtDoGlcNR8qI68H/sx52vPyS
97A4DfYJ/jgEhL6xYPSrSkZTrRmosgMXec9/ciWhesM7BCWzvEx2cpPZJMwnL+gu
WTP1xF4ZMyPNXbIu7iqIvPQCdfvL5Vl4WO/5S/kz4kCQIHHCfbDYGR/42TDtFNVh
J95F/agUPEaVBziC76pI1F0ygpJG/zs06Hku+WNyHR7IUS3se3Afg3YVBo3URkzT
Uu8JLZELZa7hQjqa7Nf7o9VV7yMaxZqG6evQ1wEQJmq4YXVTl4xKD648wAL6mlok
yaIE2YiJe7Ff3Opx3YvEw43CNefPspBXb18UfFCctrtwniyY6qs+HVsd7/XKhkhH
fr4k+9ueInVP0xCLlc9+Tue8/Gxo3Cf34z8p92PtYppJKPQ8BpTa8ai0w7013m89
tXsquoXyyQZvUxz/TXu3p++zmVk8Ho98nBte4AtMfAgZR8/CWlmHb/8jT7e8Z1Ww
j7Z7AOCmnSx031ysSPfqqeWqxSPBrSWEppveE3tjkwgz9kAEWjeSAsHuyiHPG5Fn
a0A9ZR8ia4ByEpd8iKhWQ/hzxN4JGsraxXFHN4l/yUxtlWaoIaYxWt26D4gzME5/
cOrQVcll428K0C7o9TNiOPjnHNsDh1clelsfWqUS7SzleHI44NmxusjEAEdMR5Dw
CD57se7R6MuPA3P0z0+TVsun/S4v3jQbCCvZSHWKlh4MiZlmD/P3dM1FQDWHzpr6
rc+/KITShANMlWUL1f0FgIgeYVLjSSgmvTK7l/swFzjH/GDvWOkD+RyevTREaBAB
bHP1Ncv0tMRvOeZokK4Qq973/FpzopQIeeNTmIK8qbqFgKD6IzKVijXoJxyeDzFF
asjpmCkMpo1teqGW/o4+XFlrb0EI3N/I3L7q00ZvGGSmsJBE3dssbOGHsAIXj7yL
XMD0QNjLoHMChLXfeTzw6S6GbsRdE25slRPcMlL89qocRIl+9Y97pJaN0u3Oid/p
9UpG442gisA/Ec1p+/WJdaLM9XJrO2ca27UbpI7Z5G33wwq9hHQwI3ArR9ckv3up
2veY9AitweSizKEnZfEt7MTQSYxK8fwotuFDgVcXYP3EcpFB+VkPq/1eH2lG9qgW
wWn0j1Cz6pu0Wwmunt27FbxgdXFg79RJRXn/oXcTiayLgXx627O8dlyJgddexAZV
hpp589/Lfc6Q9EEsQqDtlUQJn8kD+uwAkwqi8TZi161XUT0dZiTIh+qmo+2n/c10
IQq2mNy6f5HUFKitjQ+Wvb5uFcJ4RJzube6zFstJgWFbjdAQYvmtacVqpvTsEBLT
zWdnhBMyajz9HC4xZnu601wk685veRh3HhkMuwx6ULFWqJUHUQsTwOyksCJrq+8o
M6EL2eAgiqlYnv4C8xvDHTWP53lOsXcY94QTX7sjZC1Tptg2lksysqyvM1amZ+vr
HQ/T9CuppxuW9HEhFyrMQqa7ybVIfH6f5NdyezECSdMwUBR40uaYTKuc6uJbAYvj
aMGhw9zWLpDCweiGg1Qz7FsXszpmwLaKR8Z9XxHqhvnGtt2gtlL2lsLJ3Kzi4V9L
jFcJ8Wn1Xg0f8SuoV9AEkIMLBD/CGLkzuioX1CR7gDkG8vf7bD55sx2AxyZ45WOc
5YfBXPVw9NQazfZVbJonwaP4+pusnxadivcY/R7V6IxJ1P17ZsPWuJwMZqt7/fQb
vBLwTd1R4v7XxPS4JZU2oX3JbUrtMMK2t41cLODgaJAhUwYncwfuwpaeleGuocFs
L/I3QLiunmreEXkq8pejOe7ZoGgUKyhizExw+5CcspIIXmymFAEUz3JaLYvE92MS
WXwlued/3H65CtRBC/xglJTDAUSJx56YKR+tDVeT2OH3YgC37o9tkWU4FCokK67Y
bTqEKUD9LzOABYhR6XCZ0Vvxpk+idv7WO5tyMPLY36y6HmasHQJm62o09pb5tFZH
vNu0McC0yYfouhRJEWBhSCAzz4Ph+L5vgy7Wn6OIbrDe3rakHLk+upV4AaaHnFv6
e5rF4uUUkKf4SrBhhcfW9j3yePul9rCCmrlpKVBA54By9U6BPy1NxUlL5rV0rQXM
oVD/kbK+P686LfjYjOl+odlnKt4tAJ53fY3PKTecOqTXhZ7ciaE/PHvWoJEMSPlI
9vQdELZ4St4zO3nMCAj60d0shAuj2ZSw77+d9BsuMQ2Xk2MxYUpSnZiCN3tGT+LN
CPwP0Xk2KT2VHpvqJOhwEIEfYoq6BnZ0HXuTb8KvORAG6TYUsVPT8IPYSvQxBwIZ
xhHPDDwyzSIKhkGZY9304PX5VbsuPZQCJ0zSAm2ED+Zx3SXaPG6aMgs2+WXmFHns
ZQB6nFZ1SmEYetjd4q2twHR1MEwnifm6FM3HO1gwqYXcN4hixuBCkHiH+yzXsyeG
SbEsZIYe+zKO0vpnZUMHV/i0lDK1dhTTMGg9MsXox7y9rh03nDULe8vTXobzeLWt
heXx/zKdCySmqoz2QBfcpOhXorwXwey1Pdqj0/beF2W0ij/a0rUaX61W+GRiseVd
pM7zDHQbTkj5JPcGwbZr9l9K5iGUEJuiUnGEV+4IOxfDhBN0lNLclZ86xVw1GXGM
EierGYJzJrHMUsI4LxQJmgs8XjPmEdd47SYwB23iSGvqJFIILChgl8UTLiXbY7cr
r8SRSuGG/mqu2YOk5xo+SdlSeJ0y1Oe17DiidBszG44=
`protect end_protected