`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzUf4aF5bC3IgM/qW5fkpB+8ni05cYrTtH9gcyHje4zT5
wpNb45EXWAKYXpb8IZuCb6NAEgpTo5+3E3feiuzPLXkMwWslGenJ4DhhE4b3qgJC
UCLSGsc2nvxR7hfK4CVgFAix9FaVBxlzsCoPuvRjmzZ/n2a4m9XcHgO6NrpdIEnX
usoNPLCTwMCDqtiqp2zv3E9syTViaYIf7N7bAWPrw0B/i+LDz4Ry1D/UxEeP0OMO
kC7IizP2+FBxhxjPRp3AinieFQYcpCr5pYNEYg0aXas5N8DF/jFsPoqq0BXOqL3h
C20gmTMUkgGs/ghYlhwA3Tjkcj/72CQQuAzZcpkE8RHTcF6T1c/i2Df8YRfJENx3
XtEpeeWkMDU8+fw1+ZA1WeVx+HvdpfbadJabC0IRHkzad7unBiJqlElA8XIw4s/O
QB+I/uS3Cvvg6Sxg8ZlGwfbwKxYjwDSwzqWH3+HtalvBizWXcYGbFLwHDYHZQ+dM
YZTgnJDDg+MYqB9U6b8ahESFqBk49TcP5EQM9RTct8ErsR7IFGenz3ghojY+5V5/
4vy7jPZszF2cwD75J8eT5HDpfT2eRenj3TFAc28T4KERjI+7aNaeuvTVgkgpFCtR
205ffW25l5AlycPJYYP/y91pW9FD4Ypjh9QACditHKWoevcU10HH9Cb19g8bmOiR
rJu7oxrta+2LD3JjDNhYwqL+rDhJ4kt4Xuls/6x7/CgMeUQwOAxS89hwizZ4BwUZ
tLqal416P7u8aegCOlem8GcKt1orJqEXx1hHeBuNw6nI5aX9O5xhprx1eHzWsiHT
e+9dJtS6BhsdZVNidRhOEvXeDCKejGXRS3LCGVLYgZjfvXrQFKyRNVAs6gSIe3UO
8hP6Mv9IsD7JCHv60f/vd0bw6nNJ23GO9TM9u/Ls+hDRYAkhxgyLMwtH33QQqIiI
XA6yka+B45lvg8Os5HySZ7uf0+02Fpk3NDmcdkdDyEJL/+mZY0c3PA3P434pFhnl
v1DrwTqe3s5XUiBBeTC4N91iZZcnkJDCumFYtsEved+DFYMb4RMH0fOXZQxcfZ8W
zvkFedTCR/GHTayL4dxUNozqZvGQ2s8muk1HeJBSBVu6VrswHLTSA+3LqNO29I40
m85FR7m158h2eiuvsxrfhaU7kHVR4bK2uoeDk7alAL8gJmf5E4J5gbrgPC1TOxss
3nfXOe3TQZ+VXBAvMbqWcpB1p3qtbea58jvO7th7hi1NXqJSwOqzLvRrkEnoBZSR
SR/o7auCjKIBNiu4JNfAQTVsoLbQ1wt0jykV7E/6bfFrlQPIx4YErAAa2EWuFs7J
tIGDJExTakyCB1dMh0SyEnasMV+oUfYL17Fu8+qEP8mZS3USzVEmbXPTCJtjmZhR
P9Y90BwD2AhuaDetvQnX7/0gnVW1k9IXyKW5HVV+7dqxIWpUV9WfFbKtPBtzWIj+
KwlmV0ah6vfp1Q348lazS4rXk3G8mxM6iFYWKSxYD2fHnW9Hux6CBPUqgrQg4IOs
pLKo37mM465DXUWZmvtt6zows4lrYw4M3slO88SWmdzwYC2n9Ci2DyHN5HNo21jw
6DzVLgrhuS9WRnGXy/aHXO/0akQqg5glk2P2wv3zyGmGpkpHJ/EDvvCPy0LEw1nH
e5QNkqEhx+DPNWDyLfSBes7TKophEsdjNypUaANeQKmkKaN6K0CMosAXzeUKDEQZ
o1cLInMEjgw0wfGShRT4hDslw4CI8OIKX3iHvw1567u5NQZ8HJtRpdb1OaABzQ5r
PYa9kEoU/LjBwyjBD2uTyp+QWU7D+tCAE4tYACgS0jD5vDPFdTwJQI4bM1k1soJg
uL4sXJ+ncLSZEplET3/aoLBmYj5utgVx+s0OS9UZNp3ep+g/+p6xbFMkOn6F7kMJ
1s/4ZO6v00R0pbmpCz3+7NFtRLBhMCLzQE0s/LE2Bjuc8PxFh6NjiDZXqLNjzxhL
LCuEMLk3au6/yKLLr8FdNw414XIbdLS4FRpG2QPV2aTyAs3oxNSB7zoPZoKZp3QL
gmEOuhuxPO4SDJw4lclJsIKMkVWCGKTicaFDyqQ6IB0QkKWAnz6r0U7ZsleYTGrQ
JllYvlHqZ9804/PNWSoWECiRVDe3x2i+LG9Bc22AMwVX/X0PepghTPYYDaDopv7a
0rXwiPDRA/OsIZ1YUQ10htkypxbD+tiAmSL+zA7ecw+cXAdsmlN7ddU2JbHnfQor
b8PjKX6Zu7hXAitfkqW5rDJ2iD0bc5NN3uhLMC0pz6wWxWTjd8e38hAdEnDj5K1E
BnRlTI/KeVPIOWPV0lraUGbg/6Euzb4NzH6bpCCgCEnHhY52NGrMCi4ZAYEjjrrf
Djm2DyLr1ceHZkISdd6t6X850sAjDJNWszz9ceN4p8AOMQlJhOM27UVY76qnID9Q
z+8TPWprkX8WhpGSz+RY/qfDXRPGVsiAcO8HI8DLDZr3/nijlKFeHcXNVlGQM1Nb
X7iId/TXzUWHVggy+YbMtHD6I98UxCgTHtbf6SBrb+Cg0FNQOvsWkzvhkyOYZqnb
VUvuYxcwgI2TYDdgx0Q+IlFpnf2N+fqGmR0/kk6r/ePqHFCnrYQlCEL3zpg1xc2j
ebIZTmCuj0tpN2BpRYAD/PYOZyizlejCGs5mEfQo12URczJgKBWIw47D8ZlOxEdN
+R4fqZlNa7E4AibYN6VvTTx2pWDNvvTdDaS/skzbSybH7KjqGH13AU0L8O4a7enq
uDHtV53y5LlPPfqqoF7zH8mQSr9oerOpOJqXc7obmH6f0kDgPDyDHpQENSJe3QNz
tEY44TeA/6LdX4cV15LPeLY+YlastE/WV/I4ckiFGZt9qyEHaoHRapMYr4KNzVV1
9PQZsKb28zzrNCuaeI0cEXudkmWfFxOEr9yJFWle5mhhBTvUTpkDCnOkB4jxPvCF
JW8x22O3Cjp+rcLZP+6f3cVeW6syuBl9GHf9KAu3QTDFXJAfrSYTSmcxD+2E6xt5
wPryHdqbF0CKm0ocmjCrWUkRtW6osSy/Cg+jsUVrRxq8jOS/i/oQ0/Y8ZsGo7j+M
7SSXVchIUtyxHasU1KsQRrafoUtlyg7PNzaRbhdDrTJAw1bK8RGveMUlMqbtrKK7
zxZ9dWSwCmFlssshltBi4HbUBETk3uPiY5/yg5jTrcu0tBOdDmTWamp//AG9yMsB
rgkv6rgA5jO90Dhlteq1F50DBuK6X7n/m0Yq8821LSEQy68MrD9hb3HAbP4RYmIh
3lbkxXKKi9ov0mjqHMkjwq3xmBjSupz7YQ1GeD6efWtrXjWSwU/PwAVpg0xHiqot
Ls5Pkvp5BjFfSID20QP/RpIAus0/WdcIHkYLXQ5X1L0ZwcSY1bNMUb4mrCbLWsgs
uc9uSCx8jrVv9mkmfqr6qIhLLFn43qXmkKzpiX8e1qSY7JoymLTVxf4jhRuolmLx
13Y9ejFic89TmDlxFniA5BzeEgUrIt71fYTm8UVRSexf4ULc4Ft6qxtvDl+EAJOd
H56fpdJu4ytAokdU3CUS3gE2lvXtW+XgtzqPqWZHs5FfWYGVdK+q1RraxJ0VQC/b
byVoeWdc4EzrhEOgziXRqlmtp9tDOKW+H2KLQg8C1ctvvKvyIq3/fWfjnuvI7l7a
CznanPmlbvgt9IbE1z4W/U5U+YXOqMByrnGpEFz4uZXnfbZelyLkmhgZlSbT5Sug
xoXUJoGtwjZDMRK7wUBVj9jZ01c8XEKmtvZSjws0X5H3ATZUZ5jqlFLIvd27CpiA
VuO78GGcHwNcFo81otDx6TcZ2Pstzmeu5wt0iW7YPnf624pc0BfIVmCStft+LI/G
KaHqS/xVC+TlF1z3uh1qEl6lhpv5n1u4J2Dtjh9+NNDU5DVR0X0ICG4MToTZcVUD
JEXkwhRlm2OcPTUAdP8/otEqzuY1yoTW9//pYuxqEMN3Xn1V22UZYprgn2xG44Xl
zGyIykp0lOW/d4Xcs1meZOn6V7oMloAlKcRkz6h7dC4ayBEPLRQYHnHHdYHvnO0o
l10plkfPR8UgOuh+IXXhReuv/yF2TDSbeakMDY83BWZ27L131Wqqm4HV2Jn8gFq0
9NKyY4F8CjOceMMKocwc5GeB1qlsQVwZfj1dkZV5cdJafN51pOMLmwLRj6M7QV5L
ek5R8ShlU1wu4+ImP8VI6LBfL5KwMJ/6TcyKd2lslbJbsKbDC4vghGoXuO+V170p
bwW8TxFJssmGHahT20VFtHJRydDN5HhXqXM3px6WDYez0T5usRZqcyDYRy2lFLi+
s1xDhUVCmJCyePqP/QFrfebpbHK86iZJYaom9y4UocT78JLPrbktn8mBBqOsL/0L
pXxq8tTOYD7SQbHOT6WLQbOTlCIlXMfwGc9ek52vvWRphslIZoQu0b67DkaKjqk9
+MuQZrmUR0LbGDHA1A8W10f2StHRHckCMTFX7XAJK1TArGyXNSTTs5LhIh+9Tsy4
u2Todo3gfatGEENNdMpaX+lwO/KI5SvuLqG0FU756ofckia6Fr9ARV0H5KidY4Vl
tYn88MAiOuHCcmAKFfraEkPmN0xNsx+b+iB/HcCR41jk3EWrTUKqIoQcijGm0HJa
MLB7UKmN/bEYRaKonwCw+ymPJNnddZ76uotQDAHv3RZmyeqs5x0Snow1MhWfy+FB
tYENZBD+E5wxF1jyNfXbEdG5sLG2RXyTdrryd4v76We8z7Jkh0v4eUnhy6CHYEj8
5KM1rGPdqGTNBqv7Xnxz00hLjGITm6N7253Gek0R2ApyWWYy+wbFlMLOmiOt2qHa
F6SdSqsgftQxFwZfENG9eBz7AHfda9Ez1fIXFtNDLImlNIcrgDP89bCgvThn0XSp
tqNXP0EcqpUY0RvY+WewTpOXepbbO/kiC4MCHylTaltJZojTfeRPhWdailUtlx9K
eGMBnou99PlM7dBja+S3XZODYMuj3TVWM2B5V2daqxYbNyXIJEgUZbyaXphKlQge
yyOT0E8zE6vWCoCCD3z9jsX53DOsGeiUdANpc7YcYpFyY0ltxmMYq2w5M86GFtWe
DCf2/2CYtj19QT1pupSYWc1uSYinhkpAKh1oLDyjgwvZqylEZ9LnZhfxfSD6+Juo
3uZ/75a9py7m+q4QFQ6jp7CtydaMfecMFmr6EUcVhUAwraBG5YAVVP8z30E5qbFk
6vk2HbqGrS7oK5jq8QgTmIejP/mzX7Mo7188dtsn09hIXJiOJaPx3XLi4YlMdRtb
uUYObgO6KpSmVK4n+g/mn3X2ek09B12NKjjGO8Fk5H+EOaIOed1nEFGYni84P1AY
762YkVLZH2iweuXJCbY7bjHR851w+dwJ7u0m5ZnoT8592xNQzR9c+WbdMM6AHf5S
95GxDfjeSbbN9KYOGhC+zDk+J/Z0XNOhhmFYSAyMtsVAQW8cbH7S1EwerRPpX1Wh
6EDslGGUpPdq1LRKWkJCCEW1Vyr4pT0w5eEcCuQ9MHzgnJO/ewtaClqkckSUoOBt
zeHFgFM9nA5pOI6417AQvkB8gpXviafpTS7u4MXRTKkK85VKFlco4xRIOXRzaPSf
JI271AMyDkM2/I2PFRG8ZNpBn8bmtl0d8H/wv+VIl2W5TPREBXY4CqkqwZDw/1sH
zcbia4i+d79pcPM+EJoaU0A4yFynWvsx4CMEHpdBD1eoA4m5ASeW42abi6M4WQWb
ci2BoFCalCJ29vu2A8LK+45svP28XJdoX2PUpgbaI3MQXhY+H2nfMAmoRq6EsXrB
W+wvayTNYtHudURwPyH46OKw4JnLOQ0MZM2a5ZanKdib/62v/38ZJ/kEGuoiI2zW
ZsZn69w46OZQ451ej8dIu5PXbP4GDu7a9I6DThcY2Cp7mF7Vsz641fUyTG9ggSNW
YbO1OUFt2qQLA8qZOtUNEb2kY8UyIlRGJIQQuxC7DV99Wt/3NcULDvAE2QDjPkJ1
INuY5JQQ4xRE7BTWoiIv1VmQglUKsRqSkpkOFfJIfw3S1o28XDQa+ewIMWPButoZ
X9y1jMDyG3JOnM4pjzN4ZJxTuPzbUYq4PyqqCuR+KkvrLpyqa2n4Zr8i5KRfCpgT
zfdl8/tkcletXCNNvSmTse4UbdIdIDz5lJAOkYf6If5xMwPeHNlUAS/6+ZMJTFOD
uXBwHUvbwbzIjV8YZtiV6qxcifuCduIry1fCAULH/G/TaSxhzxNsVJG/Tw8LeqF/
XpK0stG84X6Nd2GJO1FB6UWd+fZJOnT0eItaD1V+YNxbTLDwwCpP/Y3WwIewcVQl
UAs1LY81Mg9cLDk/LVhX1/27R2VAxeP5Azd7MIDdVJW8gQtiMTuZ24G74yZZTqPm
g3EQJ033T+RRboDj791oC+1DqNH5iGsaxHW9qiquD1+7Zl10BzVlC9aOUJ9bYxj+
ff+fulnnys0BN02q1SoQaJjyHOyQHoxoFQzTnedOXg0jp0sw+MyoRC+mCf7kcGjJ
Yn+2vdsTIaz0tNlQlBhd0i/UlXsH1Bokv78t2qr0oKziO1jn2hSSmlA6wq6rbvYf
jrrHoHXQt+D759dc/+WQKOk2LjTj/WyThEjvo+x2Uknol8DV1MLfhahHkKKgbXRj
XuX3dkrh9a6IanYu+RYO5DgaAziY74JoCSd5l23WKFyJ6+BojUOn7CvdJTFO9tKV
4CbqlyckTlJY1G1Y2oRybITc3t9ZknkiH/wJcXCHs47uZah33mvBhDu3NG+sqAdw
HFj2HNLaZqkoGhMDXvDMsdpAT/jTKEP3VRWI1u0Wy2TgGO9u3zVjrldvoU81ayUp
A/qltfeNEFo7QoaunToTi6werHCBPQJ3nJDW3s0uwtyPPXtVmjKyOSgxGbMcPf4N
1vmt8k4GDxSR1nwm+6iKwayFYY6G5loovRF4101nGnIaAS6mXtlCl9NCiaJsxs7p
3hSmcPDMyuLzk2f9QzmjtMW8oB8Hu/VT7WW1ZyOzGrOiyB18GBznFLEJswfeVF6y
xCSmmJE+cJvDE139ku+onuWjUN9x0tOwiD0I8a67j9rhfyLmBif4okkqlNvsZYZ9
WNFpjRg1eQ4DnIrttvl6u2cH1Nf6/OVJ3oG+93RndwUgyqeZD7rMi9tLY2RHXyrZ
63QgpSrldhk760fE1Ozr85qlFF7FVGcdlNxjSMQfHKgv08YLZSRxqzkhhdwFMV/o
heFC+9ei2Y7l4waZhNxaKc5KovojTUloNhY2OHxr6XQzZjKO+fuVJ5bBqmRzWLOc
a15eNA+wG4ObvM4KYMORYo0pLHe1jGXhuov5FVi8FnunPhiAQ2SfqdoVNuSa7Hqs
gmS5B/jq/AHikC3Qpdzlsz2IVvshYF0l8QPMi1DWTn0eDTnR1QjH0hXl9IeweUMh
iiwV7t5uVNsM3m5ss+CcJOyuXvbWHsOGkzu21U1zcmWuTjjywi5LtUi+UWypLhaV
VbnpOdGIJYwbKufBTEE74dRvaBGtwtwbV35j2IA6cEx1zjvcii7EW4NnHBG6cw6/
bNKFLhdB5HqGOGvv8Zv8aj4oldOOjNSCQuZh6YQNx6Dg8jXdMxHrLl/KPvPCdyHV
ONDFUJvVO6wsb5De6sbezYTIsx+sS5AkRxqxH4TDl8xU2hoxUnWtyfhvsWuJ9mun
TjZRzcY2FfAvUdisdcmVFr3cMt/CKAWknj+Eq6A46thPbfyI41FtZ/559UYV2OHJ
yiX/3mp7bt68TdcAFLAcaV8vo2JcMFwl8fnkW602H8rkul6/RgKAsAq5sjzwo0Kr
kRDDLb11ip++hsAx/e8hWr2D76C9pICzcb9n4K1Bu7DN7MF/ZmBr85sS1/IMtzuB
4O9X0BTKt5+zUz33Rg6luauGKXoSIPZL0w78fPYI90EYPC08qHzOUn3xS5+pfi1q
xwKB2P+WIkieczaVYpixJeDnVlxrVpvicmyBZ/gO/NTvhOwxGdh7jtarHHjNqZhK
9WQ/u6MBuAxFdKod8OJBPwwJBcarO46zXAeJM7b3Fkqb7zz1EuE7udHvCQGVn2Qv
hbrqRUhLz/rx7cvQhsMnQku3SnYPd9BY4kwBD3EhzJSDQd695nuqzwQ9ZeCKNDc+
DhpGVSQCkGVCdWSmplbPAYXb/ZDnnj2tZCflyuEmLHg3hyiQjoav4zf88TyuNfe1
y/ZkzKBh95zBt1U+t4YI4MxnGrfMwg0XeMEmnVFBMiLM7fdpWFwq/bD0aEW324OP
PB5e22lk7jw5wG5K3dwJEe9fWpZCLBLtOEYgJBhL8jAVqatZDYPLglgTlzYFm7qx
yRVZmW+0qKkmQ816F0gKmf/sUjMg5xDkwhSs15OaxVNTv0rtulI9eQZTiVmbcHuT
lmKJxzol9ahUxVXXqJiR/wWc0wJeDKemQyfwR1vYSGkTd1Z4Ya8BE1xfgCBoNIMq
v3wGXoJeh/uFZc8ELS/XVCvrXzQaNlADShoanYzqj0CFWLCTRM6D3C+VMInspB9X
h6aBZGXgI1ZFCkzJrG1iyPpIt7zJHlxoejuP+H3xYHve4feSUEW/UQQIIln/U9Lx
4wCbdjoRn3s+xicIf2Fq3XsNqYXqZmq1nkq8LGBbeD18M9cBKukndsFTCGj5B2S0
E+wfD6SaOwmb6PtRZ//AKak1PIvVWV08vn8SMUBnxeW5cXJMFu0m8LGPWYQz18u5
GC69DxXZDBTVlOSjjK6oqw8e+f5ZT+MP83L/DhkfmlmY4FoBbJpyeyYzacCDirPd
v3dDwE0u7JIVtd409Z778xArHZsSZiFkdzvcC28m9YOfLtCFHBtpkswt42TZHT9i
7XDZWXWPuz+wsIyBZB3e0WNBnU9BD/9h2vDbIZopEpFOurNoDq1S2UF8btAv0YGx
iqSNCSqWflup1ai1BLVtrKQjEszpTIFt2gWgUyFAEipFM4hV8cw7JLed94axd0D9
iHCmQJnLXkUJpGlL/gqKmZeFvPoFcbnf41P7TgyvIf61lPJsjxp9wMMoxjQygi25
k8YPvFCMLHojtKZqDPrCr3rUNmU0tV0pOQVewbs693z9UPWOsJnrGhgfDNF03zpQ
cOxeFa9SfysXURI+RO/Q3JkI4NXMPuaiy4FhEIaljHyydVtKk6IMoY9DeYcU0sOl
OZzaQIZyQDLnLmaGQocKbWCwbbCoH1Tt/aavAIDdbANzKI4uFJ7QACwCTqvAOE77
C7mdu+ds0PQkOkVv/4I/pKVB1Xj00q5rjeP9Zr3NvgY0qNp1s2bvVuLV0BaY5APo
dsXKOb6JRc8SESTIZBjBv/qs/6vc52tfO22ZQHIzgxtcZOjC+57xSAWoiKdROUrh
OzOo/X7sOPu0WKmgSO1B/rnM7QwZa/wTRmADEomsflxxm3rI1lXarggJoFb5BwAE
Oq0ijp94PEeO9tNIaujS9jgw6DewJpitQXjBYsh6Jdy/muZSG6fWdFwXUWVSkO5n
eWDF5wh0JfwSgc0DysIdGUmlOpVwRoMWo5Ue+HpVfls7exy2Z1akFb0lJcScXanL
5IP47iFVH0ORtCu0h+3W4au9V1zvDjQS2Ry3RdAaKrs96dRDkxvQ4iLRANJ5UU/x
WmAoAAWD17+PycuZg1QZ1xPHTw8BnCB5ULRTWJHZnOzqfVgDo23zAmhRI5NzGwR1
mkf197MCiop0jdo6oWIchSzy11geQs2W+gi4m4K9/r6LCUx10kACGOHOO8vTwQ1v
lVNS0D9nIVUUYYrhamEf+b4kx78i2baYtNIop9BVWCtzuP756sr1ZS7ZS68w0fiR
Y6C1yUhGbsL6UCs+v0eVCUeu7x4FySUBz4AnCMNDiztWrCQsoPOXeDIcL9Y94S+N
L7dpOI3LPIkCL8dYvLpYHCT67xbIJW+9d9oOxvybfAMe1vnSnvdjTNp/KvD3blfC
0kjVe7DiCtPUbsDTjoujEe0B9NTo81IRkP7O9l+cgfhScpLL37EYbeQ3a0vj4X9S
rQi5G1IRwEOugz5U9I9ZCcMKBKMf2royibbjXFHHLRtQRznqxq0IbIF9Ocbhfy7G
urAdrBft+SL6QvVSqDUTwldLf50egYGt98oriA1pK/PwzQCRaX7FloGTz4VHrdv0
D4hJXBculjEuPTbqWUhCr3OJQuJofTn3YGek1U/tlXjz2Q2nJMEAOefEzhwAcpxB
k405mRkfWcMrgSvvmX0FGAbRHKfXEESl7KkNDQJs0h+aIpO4r4t4DY4GqrR0f0FO
wtzvfAmYbbS/6BVFm+S01d0mcGFeRSc52xGjm0sGsa+/NYwVcfLAsnIHPx3WpyqO
OddQGspy1xMKSRY8Z4tB1+N4CAmjn33/2pIst8rpOi0+tOYOUJiimbwDpeM51eE1
ho3vyfuOmUEDoD1EHo6JZkitZn3AaKyoYm0ctzOOks4KIZEMAn9vZAOOY/50Qe1d
RV6nFw+0Nc54TeUSgznC7KeCrU/0z43ow+I8lsm70c7s/9n2gdh6LDi1gzH27FW9
oxMF8GAV5VGgSzp3hSTz4eMFzdAbQrQnnZvTCLNNk4WR3bqPxkqnepiB0dwb1hDe
F5o2sMy9RTSkHuNYqBvKqkEwCRg7h1ygaDKyCUIt/tDAOpvNw6TUuozDOCtcLdyD
0F+eYYTyIoRb/2dN5hcpaMmm1rj6+M3hEqK3HThkiw9RzYLeEZIalkn/LIiMGcnT
CcNamTL1CRsW5tR83g1EQAnQI9IDnd+FyZI+eItK4NWnhBex5YFT1F1TWJEI7WpH
Hqz7/6T5rItThJQBpgzYrOxAz7HyemuU5b8PMuJGteDr0c33C+6FkxkYHWqqOVKB
S+kDj+yUa/dczzVqDxb+HT7hd80C8Wl5tPftz2FLBKlk/zn5vzchFd97VJ0/6kFV
7FPA2+EHixGt4gn7hgzqcXdHS+p6erPkuLH1ZOjOewfbeQGlBtx6fUAK7yE6bNg3
TZdNp2xsM9aK/9sDQVaudTJoe9ZatbhIs90UhtgEEGRs8Uhk0t9TvA2HfXNYpe61
gbbnRpxWU9HY9V+Q4L7WJzkRAOdM46+GilTjLFRNcftStiak02zf7n+q2QFcpn0G
WrQuCsdNGrT8uZDUuQDkfiUus5y+HYQ1jl5qLVgpR1SMEBltphWJmbc6EmbmfzbG
T7qyh6+M5kzFyZsOEGiypZHKrO5k8euvyjWOlePjQ4MaiD4K0xziq1kLi1HPW9IS
i+SUbL22OW5YB6zH3h0a9CYOI7Yx2GlsysS0Qi7omvZS2SiCooZuSEVhaURrw/5l
fG2AfN0Oc7royZB4zs5e/yXuyH5XKKCMZ8wRWY4/Jh/PzSr+WrN2XXLFgsvRBhdQ
DIo3+PkTO7rQkjYZDyK+L4Lyo6tpv4jgWcgYCK6QcjE7NjYz6wvqRisdUHx75L7l
6HTnMVMalMj61slI82CN1ijn9Bl4aqAzlstm17gE4T6gcTuP2te42AlgvZvgFvAI
G5l6WHyvO8ZcTIWGulwqB5d9tUR37TDBeVl0A/1yjiGr2/LaAXh5Xnpr0mezNLGq
fKjrgXysVKqaanJuLOqcWTbFEzdlTE5lhVxW7VU4+WuG+c0OHxYXYygoVGCfdwPT
XXVVwT3Cocypjo3RdL/CExhxJ97s85c73FBzoDDmm1UyCJO+FCSKhYEpv9UyVZa0
VMNnw7ge5/a0obIX71XTWnsanfG7hMMFSVAv98nustMQLpwLYKC/kYROtIJ4juXE
wglsOMchkwNVGrLlGCRBinS6sLLaYhJc+TizSsj36/dAq1HQK4N1inwmssVjo79W
yQ6G8n1u9Sdb38XPOEYg+F5PkLRTz/bNVVeEYFQrho1Jq1seRTyeXunRj+uAjDvK
I2UFqKayiCH74QddZx9ZZcyZtw6cW1vlnK9/zF6BdrCoS5dXfUcPgEGvhjykc41B
COS3UxprVdTAUNd6/IVDHGCeKACh+MftZqhM68tJlP2ERDdOKckWykvY2nvIzMdI
6hHPtfnE9gQPne8n26b6roHwNMvSHswxmOXON8k80+4Nzz7R6RBfNEI3w8fHuK/h
GR1roxJ72ysdY5HS+N20lsx90Ifi9+3EqsEL0JYe1YFKbM8trwkzPeAG/yXbydrY
TtjaEDX5LZkdp3hfcvjDdtdMYn48M0AVKYqvhDDdYBEA+50TkZ00WUP39fbq7XxK
DgFL4NfBj4udIQJ5lx3P4Spfmx+T362HzurxcD2y2cXpGXL4tL+q77mlvED/b1qz
jVV7iJeyXR3O4hyZenwBc8slcgfVExldi6gUokIHkuqR2YmXR/SU8Y+Co9RJxxlE
7/gGnzFQ2XHV0bTEWIN3gTYelZ4GCxAxAsDJ5ayfS/LY27tj5fKIaAH8lRGjm99H
GLoW0oLMhhFtzXcEWji8edSacN4+PX7tGUAZA8PHi1Ciqz5YXCGLZxciPSLaa1dP
Ss+ZwO6LZeUfgcoKUoD956I7uHV3w1N4IAThQCj3wjqyhwLXibdEZz4ynryYz4vb
0Rtvu1rq+yRlu7b6YsgmMVNoTbaXUl9amM1FIUbV4QxjSxAB3QYB5oHv1FHkGP5X
ot2F0uPbIRCC2Omz8jEL787Fafa11NK9RbXIHS0tELLjJzNPE6GyoyUivsDyO/Ty
VGvXCwe2f2EB524eajx1hliAhZhakETLX5vQmsebWz+4QBsCLJk5ziLKVPJNjR4d
ekzsgBVpv4LCGHDlmm8BX+jSe9A2ETwFX126BR9qQxV+WQvpZDa0AuAusV6ujSaY
TMc8iX3fPx55XcL0JKv4m6rZxTexoz5BwlUEINllgvIROpCBECzN/PpPXj9otDyx
cnp2lYo5mzigkA5VnbNra+9/EzENiFOoVOJstw6umEXOl8vFHgwASk7upo0ZbEB1
4/stD2b+xK0CmuhKscHKyfwxiPav9YHCpcC1G4sK3NB+v1ggBcVPARYhyKTt3xC8
vxBQvDpoiElalIKTy1ZdGETjt6t4Xn1W8AiK+D06rqE20y42Heihd8x8QShBXbXJ
BppTWzjNPaOBAaEIHq7BAN+IPG9jd5XC9lelQwlJpvIg0GHX3MNPZ/9ItqrWhNod
Lw4aswNLjk2jRlzHuwU6wVHvJjkL8k/LzZxc7TdpLPUO0TjJtW0kI0D5qSl0Ew5I
BXo8DGq9XGfaJIwqTBCou9EbFt1RPwXkvLX4u5M36PTaLk86YhZZlBhcs5QGifeP
v5h7yL6uQN/MgBQIemTnD+od3V1hb1JabeS+gBZvy6eMuGPAxG9L9K+Dp7y+aYFo
FHgZnpYN0jxsbebURWHftI9RoBMr0armxEgeUWe9AfonnjPEXGaQJSqvkibRgMTz
EIoDeHOvdR0tzJk0ByXkU9+gYb/EWVbIyWtfpXud4vOEO3QxKMfnmHfh9VCywWyr
RWlnP93ewJXicKV+QOAZ9UaCZ6hyDbhYFqOQaWmkHX4W0WNHTLbokLxZHvF1dYVG
yjMPoe1kCcpCg0qy490EApKk/6AzvZYtPtlE33IF8ItKy+NhOI9egbbu6wsKmjib
0U3lSDobCtTNCH1Yp9KEn+FflGh2oUjraFnA2hzEzIeslmVi5ZquJq78kalm9hYu
T38Homq409mRp3AB6wXrWVMsS80VSwbh6+Ba5i3NKKgcGxzxvZotoVz/t93Yr+sf
qkrfeETEKikTeixF8quJeW1zmsoWvmNeuUxRCf246/juqDFV0ANMeiXNMnQmfuoQ
cHlw3RW0zglGpITj4SaaY2hAem6U5ZUvF14uIHA9zHh+wsP1V4y7NH6w5s33z+87
Pj0+I9msAZZibryUGD0B0XXdx6QAXFQM+Oolsc/ib7aX2VB6dHKiX0cbjpVH1d6b
fFOKwjejh9lX9SBf1MKAbvmz1rnUUFCBEspg+3h1LyKiisklgLZsQjKtAVGzvcum
31ggobKjRTJHWuam7q6ASJVgdejU3jx7N2SfZlPAtO7UBffAyd17wvWB1z4pwhfP
gA/Ap8b7sqSISWaiH5GnuK3YLYktSgDUmodM0hYbALhXylQlVi35FkoXMXO5zAPf
ZrvUvTjxt0DIRYTGuSqmDGSzyopYpliqs25Cm/19O3OqVm59VjQlFSwUnVxE+/WW
DGIqh626NMt0Cl/mJKBrDrHJlfM7cjge+za9MAHYTWbbJLYQXw2Il/4OQ9VBYmkj
yxoS6KUc9NfsGeTU13YJ57x2O1OlydvZC2/MtO1eYJXHI3KOvLl9zBIrdS7LIX8Q
9ZBwyxpHI1O1M4m3pHfossRkN1mfeisyZCzF9L/8QtmLAX4WkXIkbHhhy5bTqvdE
FVw+/ZqH3FWpyTDWgsjYMGQ0l2UOACDrErMU4t2sYRjudUoZ+b65sLv+wkiar0QU
mm/P5jsYucvgCuSSEEFN0QySG6uR03QXTnpEnXsCW/GaCGiLRUzt053Sl1jzr7Cv
dutZGy1ZQK4TDRvb4qLeayMJiWu1NY69woOqRBbLFI9RRE95hJ+CT+uMBxTXMOvF
fGg8rO9xNBm+J1pgc/vPSKRurMaM89HzLnW3g7sPdIcyc+UJKjNW3GIQ95K4B/if
LcjHlYJMG1LbmXCCzfwDx5y6qpWhsDVIqObYCNYZFlxHp/uy8NHB/vKITBEqrs3j
AFr8x31i5MsqWPibqZHtjI5VyqjElvhe8pBvfKW1+yp2qrgVbIbvzNQXyiqCDKfC
vjzi5Hlou2JzALJCXp8Vk2ep/ma/mhsBKwYOo8LaDi3W2WwP/RyhooiUBPpfRWFo
T7OWx+T9CUkglvVOQrlVdLUPk2cO0XgMf8sqpXMFCm2Pb2U4cL6GWzGnJJNRXODr
55hqmXiKKgNjllBK71G6ZTMYdeafj6uDuwCl2LksDXAoIkNneY9PWjypW1Hkf9Y0
stcqSgFMR23Iy9tJK4+B3Fp0tMgfGZU1ccNxNwaVkgzyQOCHq/KoMd9RchzMZJsT
Sczj0Xl/EJBIEQGzHI+3dxZVJeDgGIrc1QDnR95xxWLSHmyXzAR9645QP7shDj0f
ZT62ri6wV50HeZddkPDdlBn+cAZ6iEQSyJajpryjJrpJ4YKqpT+SsLsYhJuS2o3K
sUBmuheGFJWNcn4p7XT9lCZYmSQtcNNncNyhWPqYHc9Pga1RkiVZC0yhK834+MeK
kr80RInCj22IYUzS6a9NAzl9GjHo9TpAjYCIt+0ItknurtBcM77UYdq3C4CEri40
1LNoWmrvfBut92o+ZZnaoJaPWcUE7UI61IweAJ0NQNYY88KBPycdNcMjZx2ONBVw
Lnpyk59CA+E5T75w30l2a0LsZyN8HvJhMJte6+5/5+neWz87NzR9FB3mKuCcl7ge
s0TqETuylvuz9QDSE5qfLyFAvHgWax8MPpZZpIR0Yoy/YD+Ir1Bxq1FRetji/Oyp
9IX4gash73KcmNSpDXFvn2lo+VQIhZWP+ZXuTKdMxeVUwJtE8IkKoGGtQGzAZ1Uc
EW1gZwtYHQxxifQROgsLACa2Nus5Sr6rpJDlfDYbOy6wy/8rdT739wiTmb+9dpoR
NlcJIcs6Ti6CmDHR71hR4dCffmkAolcxgTFJqwcrpv4aADiN5bRENAkPJ/5MKBpR
gRangaYVBKYnncpP8OFMaqUqBKHIH9j4iUiPpCsQ36/7JSUF1amDsgMWsRgIyNah
eUrya9GyoibLqUvMttcSiPhoFAFmxG2xQO+Zow2W8ObS3qjlPSnyq1RUzetEUE0E
39sjSVZWWZI4COxh647eYL0Wo/GwrJxaX1hVwjExkn/EkwbrMKu8StCSa4W2dTxM
YsW3QzHpOaFUL1XjDI1Fsv4HqKSu1tox/azwDZ8E7Uc2Y7DpbPCsJVh0xZ/fIML+
65+KwgHo5OIDtNGCGQ30htqydVoURmSrKZe61/LAaIlctX2ahIFa0m+ZMJeBLQtM
uDvwq9rfqHRuJXprLCvH85BRpaTW7SEgfRXuM0JIdS85INS7ix8fY0gLv5xmUk8h
QOsytE9dIGTZfy17iEMN8Poq4QPf+i4MxtrVZVt5utRlUo7CrFkgmodCmr1F5PE3
D4W2xihfXHA6TPC6IU/J+2Q6oWVqtbX0kPpmNIb7P2CaSGE2GRHNFij3KHAUJ32/
WMg3cwRWsCOknyIeYySYbltWNKuKGg012UX3K/qsdsZRyO0vup8xUUgr3ZtZEY6O
lLsGYLYMTweTJzyCygw2IuEmZIt7ZckzRECuXGwd+ria8BvpHQVim2F+tPzTcl+F
Rw9VF4gtDzJwUOpw/SxIoi3CJTb0n5hyUXXNPV3mpJMzTZ0ho/Gqpvjm2pOwbh6R
ATOC7IAKukviNirNJh58bbRU6GMHEsJV58Mp7H547RXxPBC5I8osFvUY88jeu1P3
q7oZu+pK1T37YtPyBVzykv1zpQ40nqgtCpwzlXGGYFKCoJh0wk+K7O6AMaWUJCxF
1clW1o/jGG/zYIygY0kQi+Jauw0k/KLZvxK7VoipPeGRT1XxD2qU7CiJWzZT+9LX
j/EHPKkYa32eNnWWKJ9nq0vSUOXYPyegsTZ7aRoCJlFfQzcnYek5r/HBHr3J4HuD
c6abfShYzp5oxha8DijvCyEBZefF8EHyw/mbXyKecBP+fLbjvfFtcBbLfT8CECm3
vtHCyNtQcAX55GACXSIQm4jKgiDtIXy1a4W+5qTMqMPt7MQhwFKlvaX8nSsaB+Mw
Wv82ctcZdM69NKJRlDB/k8hRMZc/OMTIKArI4xkwkUBmo7jfu24I/oCtPcn0MTtl
gXEasQwVbMBYOcPKKiUA4EJQJ1cTgzR44feK9zlYEpoafpIM1OnOiyVEZEIzhVOo
BWvAUMHWvR6X5LIkV9FaFw4VEqR5zzQpWS/rtf5EnixL6Cwa2w0GqxgoyhHte+sv
7J7NkR/32+dHPoOftuMM5tQdXoLAwTbtoFLkzoqGhUU1BvFiamAGoUl44rqJ+VmJ
uaro0Osc8K/jrvHP0EHNblvG6w5hzNefTxGv39IEQFmAAV50kJFzge3UKGcE8EGH
Afnjc2vm39XzAqXhIr/1sgIlpwGMrpgW8lb03BVWf4Gk+qXekpxSlNn17ju3EO6D
b162o79p8ICBho297IChL002pczj/buhAEGWjnxd9JYe3uWdDlzbgGgRvKnJR28p
Nn7VIP5l06+/867sUQKhK91B2BzUZdGw2Lnxu3ggFDlp0FkeQIIwj4LWHZSX6w7Y
X4U2ZQiFwGi7a3Pko1AcRxOCsXYUvAK3H6f5zZmhrqetbXf27O15Iuhnup9NVzSy
RLSZLHpojXCF5trku0KekCu02l/HGf8G7v7oQHarX4LtxSiCJ7tujvwO3u9JnDhl
OPlfVQKYbdSQcMXopvkSxyTs5Qa4iPj8prZc9n+R9YiP3MpgVoT7TuvX1M2rzsbQ
HjE03SKU1tdVCJB3/XPAystaniaz/elVpMPY1avfGQFlvMrlxoGCzkYsjQCTSqpr
piItsWJF8HP4L1r4/T9ebrbE0WYIlVDoPtj/H+UUEw43on5itb1zg/tgDvLx03AH
morEVa9hUP7BAm37jzfADlg3Mplu9A7giX8fHUy9zOMt5KzzWRr8vhzvxoK0xIBZ
9IyK1VpesYTW+C6RyfhFA/Ys49lzLXG6m4fPK1iDzgA+pxTUzRLYGqsdlbfBbApO
STYt+TIL5Ybt/TQRJYnHdKTZVwFdeD28CMoToaafwzpCpH41McPN10F49rWlct4x
Mn1erXd5hUjklLPpeCQe5xeJpBPI27rK+B3YL+a+Ot7UO0+nyJmjZw5Q9qrhUpLG
XA82jGxVXCXPs1djWGsrlxtZKwHC14kwMxzH0xL9eLudIRe37Evw2Wss1LXQsn+3
wosEbVVlDvktIyfzh3m4aP9bUf9mfmVhHnjPZUrBrsg2ldlDDQHxZtVVsKdtdy0V
x65LSudPlEMNP4rw1VIErdGYS7Sjwv1yOiRKkLKn2DmKjMueXihzojjSn4/R/el/
TV1mpRC+CsU9wX0DYsn/n0ggZ8ElyEYDMplFwiGJ17eNv2hDYsHcdd9AljttXcv9
X+QDi5sEVyGq9cXMQyKEBYGAPvEMSbBpYNgCKE071Uaxxur7+YgTmsti+8dFimOc
NpxjCBzVB6bJFt8TjZD4F/PF/ytpWw+YUWykNQSLcg0OsQSNt7dA5gCd91fb7PQx
RQyt70qx14nhmXjfMybce17iJ0l2lCIVYR2fGwk46VjHZ8iUQn7SMy8Zq1FmfDj9
nQKG/W2AO5MoVe0UgSxy1RJ5zG2yrlAF9LAqEEJSHFJ47XsPDDGvNc9Ie77nA+w4
aFXR2zBUkPUnR5IwnJEGds6SfePtL88zPevCYVAhM7JzJ6Lbb1/ez/GylTsd8M6q
QXiZs0B9w6MljOc58WZf9WWyruraf1w5z+82z89ZIEifQ27oVWEefqPZ0FLnd4Ye
rg2RCuPqestG6KYac9dDOxLkorEmirE9llyfGD/KmysoBc6RFLFe+T72xUxAZ1hv
bF1HUrDqh+k9ZV1VPIAao8pfj+J2U7jpKDWfydyhCHoVIZe98kh9vRs8cEyIkim7
67TmnPk551NP7S1gQFPLNpvZ6AheQ+y0pBvpW1eF4+sv8VaziskOcwVfL/e/eySq
rjqAyV2wFvaL4wrIrSVSU9qmOlWBOXt/WBpbT7dB8PNuu4kDZjNpKw0eSl6ZuEYP
kmVeoZvNH0sQk23L0dSqHas0WN6Kt/WArkcFN36wt57jt/C3Bmrj7JJiamqWsNKC
Wb0K+68D4DYVI76AHRzS+OPgDlq2PgJlfZpU0Mp6d++fgeTuqTNBTlDVAPNI0SM2
qol1SEWkBc1OrtPxUsVUVaIXqo6v6OQs77IDxlTtA84++54QLK4TthN7XON8m0sy
FwNLbewhE19BpziCy3trv3z6Scyr/oSJGEnsTTaJ2wA=
`protect end_protected