`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
KNBlPFjGuLOfV4XxjKSioWiCHyT9fiIycYTCKmSwsAF49attCct00GPbFkbaa8Zx
UVxTW4+CHoWzNbu4u0GFk/p3tvtcKMVCNylvPVugd/SdW88ID6tF10O0EVah0fzb
GjmO3c2WuJdqOzg/UKoUOrWGWm5wws1YuJaoMAMNxV8J5WAbJ5lrruQWhxcT/Wf/
9ycKo49NLc+3GLHbXtAbRJafzcaaERPLqnMQUs0KZ9FMai5VVgQt70CjJGNwzM9O
MABH9mW4/7oVSCLW0sLt26Hlt3O1bpK4mk3vB/UuhWjOJLNRctjERZw7Q6VJUP1x
IgTNTMBHpko/HDbwd3i+9pRgix0sdO1YcsJ9doujObTqLmcffL3Rofk1Ba7QcQ3Z
ZWDHUhFqLQ0fl07+rHBNescWB1RQ3+8If7mXe+WJvaB7S0tuVxyG0uqPlhahnhZc
MNr41nYtVJaVkcYIb+3/7EDxjskb6r57mZ22LwDAwGBgFeLUI+Ahwc1IpZNaOx8s
NZhE1+YArozxwm9Jw+ZoUhFsBCmzHcQcEzzbX0OSWE8Ah0tvzvoOmA8Kli1YHfPd
oFr3IDWxvrxwvS/ChzW5ty7DOKjeA1wJfkAFFf2uoMlxi5TIX9wx8jUHvR91yv5P
5U7Yr6ysKEAl8H5egbzH5t/kzfrrfWUgyZ4/conUwNz5GIIgnydSjJ7kuaunb3i5
MWl5tnLn/bNDsGLbl30VayaE4iGjKxH1F0sEZrk4UnqXakv9zqgnKw1UR9FriZTz
LdyP3MoDKtkdmBNJjl0Z7PvU3kiAdo7oAWoQpuN+lLoJASEG6SmRIb3taHbv7rFG
7zf3PPVEnmG1ZcDGIp3KHcuxNo/R0OX1kiJ5NtRWPQI3b3nA1xPr33ilrcIbXW39
k7VT36dHAxUsL5GUzZlEJULACirI3gulhTQeljDFs8Z0ujumtBOnfMF75X/lUEE7
6L5ylt7PwGi5zb/y66DTZjJSFY/J2l/6EDm+TYEgcbx3CWotgeyUOGjluUufByAu
RKe5Vkld9Ko6PxcNYS8/zgy5+Nb0up2WukGh7VmcjPYbvWBXq14fBYq1DVvcAIB4
Y5+XVX92liwHsgRQV2PpRxrSENDwNPrDDTG7xKH0bibGUOrmspIMmeFM6uflv5vD
ccbeMpbebpaKnz5Rp1tE2+lWQk+g+W0oVNxcSk+vVbAVod8R6Yy12Rl0tXWJAEXD
g8+GjXHM7hiIsG3OueJ1/r5ORbBghQRG3oQzHCorxOunJCrd4L2QoCfQs7Gqkwct
Q2B19YTIHB5S9Wh0oQhwANcxHTsPiiRxjTdilToZpSAyJPGp9Pzi1NsHkRvcbaKK
uCNbd3kP65UNlzJ/mLbAZeW9UMVMd6W5JJujhC/ImItQyq2O/DJzYGZRuQ3Pw1b9
kPFckDcCHeR6VW0lXeCF/vLIGl2+z2QlSXR+Byu2foLvy/07DBhg/lqnMWQG53fA
XFT6bYPd2Yg0fi0MliMqDanqjuhTIjkVriKiOBZCxn7F9O7mPRzkxIOFNpmzihsZ
862OJQM+pSSAGMKWG42Czy2L907WLrMTVOLffTi67nmPSA5QjakD8i/7NGJF5G1Z
8QjfqqKXm1EBrl7h515yrhpyxBoU9CTJJcjK5krJainCZoQTxH940cMSt1xj5NY6
oWSxsgkR1pT531xK+xn/a317lC2vdgFHtAkz4vqy7IyiDQXeK/nE2wS22cxOt5zP
MA2Tg3D4ngiYv1AIBHwCQx6A/KUwMFGH17BCAll23diTKAdJSb51GBNd1UU63sbV
y1Can7q37zOb+dKMdcs2kUOtt3ngIk4FFFFUUltOWMcK3E4232shr32Jxw1QKyLE
2Za2QXCMtANTaOiu3ZHLoocS5eT9wHWGqg9F3GN2zq++IJT2OkO6aqXODHdZI+gE
ueacCrCcP+BPdSamPbYBHgA8o3lEdIHUa1Iglv3/sVD21ci82FmNb533oMt4ZXm1
UE9fbRO5NOW7WprcfyXush9rEzEvheDgYug3pbEsenAr7aj5QLBrRh8CRo7o2EjB
lW81s8kPlykfCe+pesUrPIf0LeV7c7dkjIjaFO4OGc9wrlwJqIuKk7oaVZPMpYpp
CuBBXeNS3k51xajeMQi+Psn+k/LyjqdCYpSoF3M+cZP6k3xz5VElyajhilAb0FXv
3KJ64TOKYLA+3GFXCS9bjDmaBzs0z/qSxgK8xT5cRJuTZfKxhGCVQaC3eMs/dusw
XYK9DsBFuy3Z1GuF5YC7SiCSjOEQ7OLwV8GIFK1VscyCruHxnqjz9cIgXGP6EQ3h
fDMHklj4xUsZXOi34U057LZSlIWdh4A46bDqxfdJdtdIpXrDM5NykgIJVawJ05Hy
E5pU2vlI13JvoJRiCh5GdzoMYzHEyuEL4zt33Wwl1nhKdJeEaGgnZlO+f1874GaT
4rdphY7pC71QovtfxHohFT+EugojWV4ldSYepVUPeyTXM+9OB+mj1ZKBu8vHc0tC
VJ5zTWDKYBzvIAuaDWtciL7PTkuOSJSNzPXaGE8oNs/Isj/EcudCXjA7xxaGNB0x
C/voe801cSDxLW8ppi7nixm5wkirk/uBaUub8PcoIsrhu2gdn9M45utlS/8YKU6l
HPcemq+JTTNrcke5LHyxBOcsekqyzL0UdTzNk5YDOegZMIdcUaeGWXM4Bg9YJR8o
5az8VLQz5/55G1xx6ypUhWk7u7oJSYvVwdaDRACl5PftADtLIFNcgz0PYgh9DtiI
FfwBbOKmka31QthWqscp+4mhEi9tbwrjcMM1a1zLHEX4YHZqklPffFJsF8WZMERK
qfo52C79KSE/IKTpK7CF5xwlS9/MPvkGzA9PV03kj7AWnSYskT+mbVcKh3jOML7D
qiQvqUtL5BEbdmnTqsw+CklpwszEh+KRL0pRp2LCKtL1arRqYNTxWM5bl8dud6kh
X0eEywvfZ/vEpGvrH+8zCFZGz3m9eSJufCj0X4JIObgJpb2vdKplFchtqMQ1mTPy
Y2vdR47wUzD2jguCNm5lEHH091xBJx8tVdjMmaHhNjpTzO/qDW93zV/npOL3ZhdL
2iRi/7V2skm1MMgGjE1/6PDMYKUNLtab1vYBTWK4mEJrdv1m+riO4rSpY800T9uU
oJlWz0fpe0VXHa/p0SEHZsvlhdhryl00Xj8zZfSpig7MfMiJRvkGZfqrB9D6IpwB
QtuSHWVdCi7aIESVMehEVOEOamwRYfC+Xzu8hMNK9qWWj+Mw61WBAJN/EVTg7dH8
28Hq360LIjYGL8pthp9cdx6p2vszVGsnr3VOCNf2/agmMd+tkNOsvs1f6kcC3I1q
SGP6y+gSY3GxNEwveJx56tH2Muj4Eh6KgtztTUb5hz3RBfftSPHsxBE2RNu+qsrY
JXnRKpH291BlgiYZi693Lsv00AtVmAxlxpAMtQZP4OjWOLNxKO/fS7W3jsZxymUb
RS7XNEiXmZ7dgu4CS6zPO0x0d7C6+q6cs3VEnEk2EM7E15cX6tAZbXN0IcSBR4Dd
1741+oDJl/iddW+IqWir+I8vjSuICeOsfzHYU8zlmYhiIXvAYPIHjAJOpdIa7Yqo
+ptz88xK0O5jwZiCHBwLKbd62oKgzjlzoopFwFbcSDLv3rGsvsxhwdmnkLpO6nLu
F/Q8vaVG7m8UxtASitSApGcMcMxwh1GZqbjFA2xFFs6Mh85tfQ+iWH1VzgwB2CEs
Kj63J6qApmbEexTvcxn0Q+lkHtqlPhzyHi60wD6RaimculaLTQqmJeMnQcHL6q/P
9rp7L1uzbxOL8cXKgLxYArDwH/lK1rCv8wW2ZE/bn8+my2IcTi5wFCxDoL0pk/mM
jSEN1Sv7OcMDHFD7cA2/eFFLKfxHsq+eeImRL6SBus8hyZNkU4yDYnlDHmfU2gYW
IFN/+SIDz4S+HF9NDTt8JGHvdCfJA99dryGHD7djouxtwJkDSTPnd71BtidhzKyO
yP0ztandHbE8Uuc4OdHKRIldaxNpS22Szs7NFUaGoqen4yR84jkPLkGr4OV1S6eW
ld3vA32I7k7w9yin15kvdNTNBj/QOwt8uSw3DCUIi6o+PfF5WSKlG8q+AUO8AXjA
NZKtTcxqY63Y83tkDhib4c/y55c+mVT6oGdcQqn2j8fn3jolfkyHJ6dCO2Be1xq1
MLrQHyBP5QTHCP7ZPg7sGxk7MdJTY0XRlMF+5t22u4sp6/F79g1z37xd6NFuegs2
DyffE3UlQ5muOYIOF8t9wZenHB1gEqRPWYYTBixftUlEpxW3OLa3OscLwlgb66on
ESYDnCNwj6NWJ17AR0/OxJS+S45FhJ2AXhJDtFhd52Cc5W2QAI5rWpTFWpauytck
7uke//BK/ucxMXHae+iZAGdF8XkL3VVFFN5E3ZlG4deW36ACuGH7AdJfqfd0S3kf
8tt/dfyzHgyQ80zjRRfH2yuAEnwyedfJhYat/r6hhhHTpJ5ymYFcU46owWEgngfs
TRrHt13bvJWhGoctacZWF/bCorZg6IFpMc84DrvjpN7qJIY9Bn0ccjRZrjjnmpZ9
ZoTqT0s9VM1Bthig54NsehnUEc0KbQlaSVN+pbShm1be6tcTySqogM9Wjkf7DIWY
UWhcZSThedfmPP4U0P9KhuLgTGS9XEDOYmbKpiG3hEAjvQFvZ0Z+QvDQfqwLguhv
OZLpNMye6i1/rkG2UfIbaZ12XRUn1ORfkERtBUVkMyLsZJy3I0vQQEN7yUwEyAk0
eM/DuXMvaW/yTDf5fnQ3pu5kgkaSLcYdYWQocjeYBjI7Nh36le7MyPwydJsInBeV
TjsZlDz0zVfuR+GcYkhGylXKrshRGKe2J4uUZRC9agFweHsGNsYH8ESN2VcMHYkz
GhCrclHgW4laPMjLa5qQwnrKwvyPsMYfHaI7zofN/P4bjla3v9MoVmT9+Q1rSLSd
OtLJIhYgfQ07znVij5nqf4xELjzu+4wVFbeYl/44/XRfKicJIproL0T8jWPKBDCT
q0NRa/mR910bhK0ZkbXOsCQ/ZP/7jws+OPvSp6Zs4si5t8gNAvqO872zfZP786L9
9TgFWFXWty1yZLGNLbKRyO+comLH0dyio9rpo02f2VupJemys2pCYLmTVClGsWDi
LqXyVDFdOo0u3iWf/62PnTOqoVWrrTOYOy6v7FUw8twiV0oFqw1VBxNXu/4eSEPt
RGfoK0aknX4ymONLxrGXtkQJ/Kk3ulLqmVdup2QQX5B2rxy8Yu8lBU+rXqvlzlvJ
s42YGuAnLQZRZUlxHX5Q7iDJrm8Cs+BA7qn2iLAVaGJ2dx2jLmeqZ356TLf4/dnf
xeO2vAAhiph02uWyBd5cNt8nzzgHG5LnkYIFRrBXKBEmSaxUotheqBFKrpNNe1f7
nEUUHMsxSJdYrSiSH1jDAmyqWtL+rCyNL7v4e7eZCIH9Le4JdqEo7foHBitn/tbj
3i/xrSR9qZB6VSVrbCkfde5cnDjajKHr08YGmSZFnTiL7NzpK20G3s98z5hPU/To
m3jHbyiuEqmmrXpKR+sysQYkP6KKH1bTu8IOr5bpH5MV3zoqgUin72Yx8sds3Bnp
e2BiNxPKD7PbP2sMFtIvbspcezl+390bGa7TmswcmqZmqFwyDFosd+LPOsBYu78v
s/x1f1glEx+JrMcgILqIJGnDwUqwDAEvmo+sRTS6fvV+hrtQl9CUsBBdevPGz7BJ
fZX7IKny6xbQJ0FcByyjdxFtomz1j7qiQUi8NxnXJ8mg3yOqoJaJDSM67mms+29E
aJc3praIkKEMPDn7SqA5hErdqHnuTlecBvZ0mMggVKKC+uFWWkLUYb4XuOxHVhc4
a/2sAmPm/IX+0eJYiP3nz2KIKmxv30pPIoyoDSf1C2BNwQlLlornfLEpBXAd53Md
nrSda2qV2XdJcGGVRjbK5BhnxrgoPcbKqxcZGGJjT9v7tzXZyy/2Rg0bNX9bxkXF
eVxgTgFQ/JL/oHO6IWUe878hBHKvA8EfvDb0whzmUctHTrtWecL6L8puJV6jlGgk
D3ijNNt7ubst6ilSgjwW/VJQeTGXN0qdL/+mRRyu0lPoNau9KegQ+pvtZ9lONltM
VSnnO23u7Kl4e4KXZAc3cJaO+5oGg9wdv8u8kbeGI4H1HZ2hBCkS7DCbGvZLOG+i
B1cXwnt0sSTKBPQS5yMLASpE1WP0n7rRsqlfswJF4CBmoSF3m43Xriv6yXs2CLPo
MZFA6nOB8Z0JOkDv1PfoHxre8oxj9wj8wSrMICEuLHSNLLqZfwxqpNDOcmmnXAq3
i4IlSFBqJBm/ukFCbebh+m/HYR6ZYh+fYtxPXiqv+/ME2zYUdcjH9gI1DnpKScy2
62lx4D6NfytaNiUecv8wazzaEwylhfevfCWo61Cgx0H6otFp1628WAdiQ4s6Tl8n
ahgwRysLkpz8Vd3LxLfHFwxS12acccjfQpbSh1oYEdXuMQZRUx98GtkD3xCYhct6
j5T3umNcLfKu4NyU/AWuhD9Pbq48gksfqaHnFNG8R9WSzBEoj88JZg2lWl1zmwWW
IGiWFJLo/j28RLHs4Cr1a0+QkL2TLYcPcHihiXD/zUq/jG5jIY9nTbQYoaJkum0G
/sGNcIRh7IXvB8GXVNsmYvAZWerE74pbAYmhjr87H1p7sM/IAPCTGDt3gsb5Od2w
BA9BqLktUJ43jW6//NlrjfieYMNdgqSnW/91VTiCHgFBO4rJmSUT0colXr//zR9C
vOxiDecFpjW1hx/a8p5fkDg3USIbMhLbnWZt9GyCAJVH7tPerFwyDrwRjhO1gGkZ
ao+hC7/0vx/KnWfQi54Fevr3ndDNCNmPlyKomwzFB5y3Ldsp5FCOarRLo/zCpoUu
5aGKDy/3hQ/NkDSU/aLS8YVdOeY5UzzQwvf+E21CIzhLOaSu5B+hLW6GywtsqmZF
bnsty7pA/Xd/AaXZYSNKaKL/ec7vC9eRHSy96SqOemc2hFnRh3DB9wg7DNed6Vz3
OO3AXqXeAi1t0Y+Uo+i0CH8Mm5jFAlXhTJs1ZLNhTnFg0ZSO+vdRofRlz1dx4YKk
sOsTJDbZgzTNAlFQPHmoNs3NR1okHP46StLjdKrao6M=
`protect end_protected