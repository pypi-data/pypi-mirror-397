`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQL//zLF+zjKVteTVRhUGH/5+XMLSkvQTgcnYBLgJUcK6
iwFzLnIfdK79I/DMnaWJu28OqdgCCsRGOQCdxY6T26ZrdSsVBIG6gz7E4hKgUX4n
kgpcZcQ4Mxow7C3GpmQe4sGuW4bsPdQX9ioV+ppm3h7VkOtLPGBC/hDFs6H2wqlT
NOAwUwHreBabXDFJ3PCwtVTCRAOW/IsZQ16dkJ4ySV/JHydMA3LCO2vxMLBlDILS
LVt+tpR0ayGWqX4bjC3Z+iyZUz92jyc8yrhozvRDYFRx36YIOw2EqACDeUfpvXUq
9wK3nAUFXYiCxvVco57yjsAikrN9E96NM/qINekeftoOOIRI6EPBeIR6HicY17CN
BEciIag48PG2Jx9sLaROCsC1em/oQNOjUXcfFxknoCtwMNXFo8BloVr3kPpl4Qx6
IMEFIQHrQaY6Ar+RJrgI92BGUX2fPpO6r37nUeB+BlSBOBJkDAtS4hwc6sGek+V0
o3MdLuY0hS+eJ21Fgmm5a7PxTT9M3zhumlfVsCunFKsH+61RL7Vw9tri3UbXkPPY
nacFSkeoCEltUXkyhi+Bd63yYDLIvO5pa6aNhqaALQhQONMraLWmut6mf0UBiClv
Y/L9zY5D9thgInll/MOarU/QPItEUj1zRTJ1cNSMjrTCtIKTa84l9T5woUSIWyy5
XoOf6fWz0krR9SQivPbPWUA6B8L/Tcs0Xv5JXRWamERCV1gA80YNW14ggUDX6g1D
crXPGYE/GQmwsrK+VdF6ZkyHOIuVPlH/AATeL454MaVS/yvg2LbVwIKA/Wt8AA6J
3pXHEjRqj8vP9NIUfkM0fBEByvTYpGCO5cbIHC7myJoFsT9YTLRfHeCdk6Bya1QB
yaefUtIolGnDnrJiZsCkllhsnlUZ5KOh0Tdb5MXSJbdbn5XKGlUZMEIhC9/LgKMq
+wTNKK2iOX6nV31XmblytuM3u++mDocIkiK/Y8ZNKANMjPU9nqxKyGlgal8TO9PZ
hkcXwiauOXrT7o544s0N8rXSynjq9fPchN+CtWD7lLPXCSOHSrG65G7jw8/GG6Pg
wZxIJYscVhC8qNzRpDQwRwQGAKhk4Y/SRicrfLDk3iKT74yc1H85PK5aS9VdrSDi
5fQBDb70MWMmDrqjI/gyUPgJWV1pf8a6Hc7DRj80y6k9DV7+aYgipFefrS5vqn0m
mzTC7dAh2UKQkM8iPoMLYqe5fVFqa0QoZn5IQS7AV9E2KiO63JllRk+EL4TlNMzv
/m7/2+gTIS6/8m4ndiN5d+cy3Xxq9g8WcHGrWgJinzWkdf3Ka9zH9H3C/06a/cpu
CPFGqeQxxsz1FjyVfx4Nkq1yltQ2HqwTxffZlglOaMfz1yw8FaKR6OHihJRLIJBr
yFxj35T2LtMEBZQ7SNUbQCl6nOdNwWlT65SHyN50cMvAcSk/ZoWyYRD6/QZtBrZ3
DxCY/1GfgdJZO71kCkTol0AGmMHc4daBjMJSfMSAwz48gEosJmwKQ2v4Ty7/DHBL
p9WuW1npwXPF9AMKG/rnI4qMkcX9uWbEybdKFJGZHgZ2lwNc6KDBmQGaCnkhVJcv
3nrW3g13hRGfJJBx1XItRwMnYExkOaobdMWSbIEbDrcRoqa7DiieRsttXOaOcJct
+RTb4Uja9ZggcK57sYoPMSfDp8DpGlWfyyHZnox3tz8+mJzgdi6edDNPhlX+2x9G
1NF7VBcsybeDWaTkkrNlXkfxPDJbuxzoggF6r1Yc7DYOsnKCmg1RANrXU4VXwpsR
eY4PDOUgyCrAQ9IdmWFm/NQkGMzFxoJp9LKqf+Zo33BUBs6ySEn5iPourGQfxR+n
LOtw+7xJ0VBZGaGRKtqd/ez6RPwlEkLsthS+jE9E3YQ6nMdPH5MZSw3eOgPljN3B
Ew47IkianYfs+4MCF94bKPMV77D9RGSWu8zicqCDx8q2aMCOf0ICmarCnCb2XBew
k9MgMsGCglkdE24Vnpm6rFCyXO51CUaHGW5no434Z1mMhjxeZ3s57PTlCRgK74fv
9GJtFKKEYe0BZns7O4NC7LkkIfLol4F1fNxfaORJAymi6MoY5phDPtZkc8LpDHHw
9cbWygnW+XHqm0FtxFMJ5iRUUrkhYYFo0SqcnfrUvBhM6WUkPAmU6s9kCz0cFzhD
2DFU7a0SGkC5oBhUFz9uVl9ebQFrsPd+skJeQB0kGbR1BY3Cg8R8CSTVDNF8F5KZ
B7Qfnvqef1caWm0zrB2Ye7q6acZSxUNCSjW0nE/xv0ll1kyWLOjP1yHKb1IIPaT9
XAWAsJoPtAfMfZz95TtlWG7DNr1gmiVxZC4/8uHtR9DTq6xIEGsU5m1wmOzoYnIT
Qzmw6pe/ucb+dnO3brNTCAuQ6n4eiBFtHiyq8w/pC4Q1S2jJSJQbw5aA0DaKO2Ij
d7eDB0HwPpSIf2W6V1++wb+o5Q5Ar7B4KjqiVk7uDA1maosBhVLKjlWf6XQneVkC
+mQ6MykZXC90KmrPQboRHJSua4j5YVdnal01QSXcz/+kXqXhWwSXw946fYg1zvSQ
nd3Lt+UNYxcLU5t4z6uyyiJHUiNBx9hWk6XW+EubrHryH5tNMwlMOBXbBKnphBfj
Xpslq50WZMEhXLnQPUuO31lMsG6MfR+hlYzznbTTnKOLg4EPvts3a0HyzM4VSVTC
4+17XhUjpLL7ZlO+19eyHgrQrGcgcbH2c/KNQ5+OLhDUbOszjNHKYhZ8wz0MJd9c
GmFP9fPc5Mwjs+Bpw7T0vPN/YuNvOWmvSJydpSMyHCz++INiLam3oRjjTN0Vh4xe
8+GcBE5CLOjn8xKr3Tv6T/nM2kdh8yNtwiejSZ39caPmRD5s0M3gQwU9TiD6C/cW
jzMsK4aPSkwZX/q+il1cM4+JNyVHxZKl6ZTWgdwdiG/ecgLGzMcD6DXteNbwdBpP
5eFYxe5aO8nKwqfjW4IrEw4KBtAweSbpwVp7qmhAzSyectY9sYB18bgCC6jXA2NA
KN5zjEbv0IGpFETS+akZYeBIRfsBamXF8NZua0GOGU99mQzW2B0VpGtPyE+qbsaB
9WvswAFW2po1tVUmWvP3Amml/pK20RieGqRR/TBqN1AeMwlw40B6n3oE/KgwyFrp
aRUM75qEKINqSM389sYpxZX/2XvhcGN2tRevXK/EBqvALansenDdqh8k8BDOUNh1
e2ddBAb86t+897HRFfLSFMn9dyWXausVLI2le5VBjTED0SwI+g7WvlujmEgHtLhp
zNq3Ukxy6zWMZWksgqM4zXSAtdLapR+Ab+um7XgwJveOJr/bZ05SHACj+3WuKzYh
x6S6RfIyeySzj2F6bHCv+H+yF5E/zv93H2BpaSC+bZOEKusFpthRUSJN0giDqe5r
rZgDcgbsRq+vaSpbu8PLzzb/FVfuyhLvadVmMIDOAloCUno7yceeM3XHDVBcLDsn
FblBVZ0ArBtIDaTXOIzFeLGvuv06ZTY/K24bHK+1Vtq7N1V75GRxPxLfmlu2GAvJ
eNdMhNgHWjFu6mux6M+RLn2A9fSLaxMXpvajyEi5xeYSYnfpnfxm4UXGHVlJyaEA
B4/voOdahpfBU+UkV8DqfCgHH/wMarBNxAesgcaukS5+uL8k73gkMp+neCO+rvgt
8HH7L1GSJgBGal+KPNnDCnGxZ6vms6pf6xAlZoHCcUm1uD65/qJ7LebMcFW55Rix
RR6qMlUfqrKrq5yBTwHjL3gX7t92xmxGba97M83chDnVw0MhUnyRg76OKcUUhwMD
5fXXikaJG3t4uQ9HmTQCz93Si8QKAJ1x3Bq0kPC4xI7PMMavXNqYBNLzQISDL4+b
Edascu4kl1Lh7GuPJhS4f+Q32KRw5UHnMqdkfTuEqod2O3EP7Oz/I0gqGxZOudJQ
jtN4/RrYiN2AksSAHkeugFucAvR8BQaNXvjJq1BZJFNb5E+lFyHFs5c5V4lmptjw
6X1XZCz5V3C60RO73vpdcRKfhGlvwYgMWOE5FkgoRsjiWp4N3PLYmBulPn95I1AJ
6/0uff7SQMOh24oivly1okHtWpn1lRjbXccpUVTbtYatjrsEf8kiIXIV5MpB/8Xt
D5bv3rEWkNJxkDM8qSbLVGKomq4x9Sv0RXdkWmz6PBnP77U9N25QIHbcoc+AU/Hg
79yiGUx2yVIXpGGvvbyl8ikSvFLH5mmvLgAT+snz1LwVZuLsxqI2rMTux+Lk6UtG
jPJmvHDk4jPu7NUJdmHEYtgPyyfZZoORSS6Ctw2KkmN4dgUl69Ll27sPWsTirf63
oaZVCtjJR1YnDKKZ6vvJCvWg4HbCD+qjcL+aVKrZ72dy/ChZ8icy6lf28jQkE8eM
5Gr6zNBt5bP5+rNZP3y6PlIUSdn1tOhR68e8rT99Xr0G7FJ/m+yCx/p36LrWH51N
q7czgDldw6jkvJFetbI1XQ5+Is3rng6i5FYnw3sBorD51bLblREj9OuFDVQM83Cy
JGNRGC/zZrblxoqO/TYnsSCZlpRQ19Ewqx18FLD+9pYF4Y3npz1XSWOmaJpGYa3Q
sA+LUhQtWP5eQPZYqiWtChfqVGAyu9fYi+zVAGmYw4YilzwZdnJNhv82MXhKPgZU
l2fe5fgczBV8PmnGk+8Z3nqHBajlZQepO/olxIcGPd7Qf4baWbcX7GFQw5LozRr9
HmbkDaQFUmCNQvJCcFvIqlzKY9TagchnYjI+wiBkxBJwqgTBQpYzLlE4gpc2V1Oo
9eOtT8+d3dUvhSe3k473uO61u3ON03kXhiikXtFf3TqlmPlkUOuGfHLJJqgTMXLZ
Mr1Fs1qklsxPHlW7gD7g/XB5lpMqbojDKevbX5FvAtyLklZhCeZEqTejXrBHI9i7
D4uAlhZMBCt2LWw9eBk/wjFf/0tlsV4/ck0rNm/zVUTE97/aOhhnf5sHmjl+jRyU
xcWDdXsm7gPc7gCoId04Wanmh4yWahxYOLTYmF4AlpCx9ZLqlHvAfnhYg1IBYZZ1
p2LoKg9iLT6CPYHCEhQ1c2dtrmtQEd3b53CSDZGaN4LeJ49bJnCGhEQLT67Kw4JX
Qen4zL1JPs83UZSrQLMhEjOEi++hyYQibj+U4Mxrsx4HKrTwtXxONYmzIYG1MSrc
1SIBgAmwtafMic22PJccDEkNouBX6VmyDKgnirxppZLahhRzayzijvVFOOP6YjRT
4ClLDCVm/n/F7E8JXiGW5L0NS97wobOx4hNtlJVh/kXpI+98RnkGi/2wnhkpemeo
JrTjz2eduEM7U+cySPgZRLlTkW+6whRAfhV4DTZ2n+2wwS3GkQdCM/H0Qs8OtcSP
5lMSWtCZ7lhs5TG7/JyxmhnEo32nHrpadtK6CWd2ZRsYpG5ul/6xtx1ytM1S9hJ4
QPMxYyH4cCvXN3a0BCiVqaUt/Nem2VXfQ9f0NDSRLrnpbQcQ11DdewBCjQHnSaXr
DY6Xl8ocw+vvq37uDmhbkpCQUdfR8KC08Z5sHVEzgvu+ArJ+Is2nC6n6D3o8vUCH
hsRP1SkkoJcZZ4U6SCXr5ENg9xfGNP6g+L5yDiaeOagig1IjW+evuYzsJqEb69WN
4lNczReFBStds6XLeUwhuCea/r2cALgzG/OGAcZl+NPdQMTcWTiU8GJWgBApsPOX
KH0nmuAQO5HW4N7+ZQwiWENlcjjCqtyBKWTeodqSYVaF965z8Ed+byHx7VC+5OZ2
hD32RYMXbwgiSZYGuEG4Fs7iMHPtKe1JCso1xqh2Y6qCtrSTAdTIdyfmztRbB7cC
XaUIX3xZQyAjJ/nXDG69P2O8tHCeFyFFwz/vsizeWFd+PwwZyiFhzLzA6e7XAp08
XuIoXbmCg8ypZU4qZ29M7S9KTADrSPn+xABLvdRJltxDMD7bFrjXnBSUmWDlTLYe
FzvcXWHW1fa4lxjNNXYiwFcE5HBYSEoEAsMx0JqxAQsV4gSI2biT5N+Ma9sT9pOU
oisZrtM+rrMGJC+iB0VcGWf4LooFW9Ci53GtuR6hMUif7yJbcSLjZ2nQ61kc8AkM
1yoTXWR1+MAaoMAMMQDdTDlT1pNwLfu51pIiSneOjuQwL1SycHQjKpQ7brVwYmpX
xi54ihoQbeuapTHshqxKI8EltkY8IvDTCr48JxOoVPXWGyTFnduMtPU21NJhGYsJ
f4uJv0jCBI/pCToE7bAMT1ZsItemMGa0OMdX6/+f0xOKbdfmZKkSsIMqLyPlgJYw
yEAULLaqwLQz/NqSpd0yl8U9cnhYNBZpmEGVVV0OPxsd5vLgLM5EYrRSnFQWg/N0
UxQSKKG1xJYgzQwfujCMWSP9duc47uf+7tfrCTfiFDHLW3HSNkD80IN7KRhmRySC
/4h9fRCDvhFz4Y5Uxp9jAjEE61BSrvOdAjXCu8vTGrWo5sITKhfSqUWsVmYAUCUu
9WCu+FFifvHZ3shuvEGL+fzUgocjx5FlyYqRDL6qnufvdyf5xTsbbXApIjtt5S/9
4sTlVp3uvIuX9QvnpYT1DHIxFZdtl+rZ4bwr5r9bhps4pR0PVYKFxak3mFBG54tU
SX9SosmmeUQUOuQpfJ67iPgpSbQeKFVo1k//MIR4LJectGTXcl2xmeCqs8KUsaV0
JAW3FYIO9yRzyO4ILmplji5cy30fdEPkww1zYoCpa1/h+yK51iUI1edavDt+dHoK
lgb693gISkoatL8T+A+csFXndhUlGMmA8gPCWn6ALgvBbhnFKAd0JFsY6Z7Il0m1
7MUlp/UUXcqky//7oE2jFTaYO7TFtbhkbnmViJ1lR/YFrkSR3D5ZAlsse2DS+HGr
deFMwkNU/aj8DKjxjJ+P0k0WJG2Xpx4T8lMmWZb26hBhLseYlC+DicgzeebycrnX
MRDb1RRGtf3SDPqDVWuUcl2VxmouaRP/Rb//Bhoa7JQ2gNLfZdcnz6znwSDzzD5O
is0ui3hxTWW/JdsP+2KyqM8SMeLbHBjDSEltqUbqKXJf5SMEvIys5/fZKEKMsBrq
55ps9+BpPJpaligbF6Pa6TBsZLnPwqkCAPzZHFUizBUYTgbKMJkkqvAHSLUJJALR
wG1hBSfqCnRKi6aBIH31pBotSoCSw2fsef3J0atesmigd77SKKOEl7oPK6wGfndj
Q4W5T20Z+1JFhLcJIFlzKDZDiEH3StUVC2oCLPlHMBF2Zsj13tIAHLof7+eqSeMz
8rmMc0cvqyd1i1y9b8PP4JNfuqgdocPbqqxfbJ84tAyAUQkSGnGzK50R0QEXYLUT
IXnjJM8qIpORJZ3BAsPF72NlR2ZvcMBpYt7JnSc89VbBUfr3y234R74/OkY+eG2P
KckEaB/hCAQoGLfwuo4qpGAdKqRFeZIIdRTGtu1Ip+p28Avjf+DUI0+UzNO/npio
a2z87LX9Itbt4l1/laFRtizzEWx8WIaxwqaEv+4Ly64o882yOPMdiQ6qp29JWOlN
79ImgE/tJYZSus+64X2huBTggt21bpHybcyaOCBplDsf4VW2coRX4iA2zVYKTS4E
ZqckItFpW98NZkHydAXbo905YrT2ZDYcgZJcBnLLP9ZPcJoFeGZnbtzIbc1CiwDx
P9NQ4o5we1nCjAmmlYSZ9+nI7mVBjPa3goD6b6UhgYEutVbSgZQ7si+JGle4Z0xF
oAD0q6wzUG2beNMCCvg2lNL+sqvscxkcSoNyc71boe3RWN1doBSWBPS5Vv15cnl+
IaFcANFVeh0VdgTalDoXQNzwtP9PvzMj15MyzkrG3rqiHjrnYTYULqu1hvlLrJA0
+RtEZb4U945zphbNclJO8Rj2QOjlv2HhCHz6L0+XgaIdkIMY6ViOMmZ1Uows8QBX
GH9boC2QV7QuDtmGSsG6J5OLgR9w+EUBBsEMIlG2qsjgXf4i6ItOqaBKYLxkIG2I
GL27H0cq2V4wN7U0fDrVdm8bnkv073ujPxj4PQmuZJVoROC68OQQ/1Fg9SfjMyNA
2rcL1k1EUV941aHEoihjk83kCbOcgbckdd4wEST2jjdrdWrBWISCcXh0O98UUoNm
SicyEexYQaBcQHR7NuwwKYwB2mps8XmfyyI28PxjAurhJyPirkt0XO67ZsnSMS5V
HIhvui7MTQbFzieGzgZXwTaa/Ghty9Vxx9PXjhH9Gwm6tCibSbVYaEEIBPVdeYLX
L0/QOCDOJcQTcPuZM3CKTIunSbpkIg8Mb1MpM+w3SLJEkleGwNTDrtwiNzHgl575
zADQqAPHtslJf7iCa2BGz2cwqDzxRas04bMMW30C18D6wd/LqzDLG0s7GHWvtfnX
jx9cFl9tblZ895FN0VKnsRldTaHpjRbehGjAoftSfvkAnUwFWlrWKMJ3+mhZrPsP
5UkOjH3MJlpAO2xLgImk25JyUMUCl40mSznuG1ql99WGrPrPKBLaT47n+avP45tr
VQQ/CtYJholUXVZ6NR/4j23FsYvwODMENEqIjL6Dfw6HJ+Kczr/ZPCrDpV98ubq2
Y8bgW1w+zHEc3OQgV/xRpWlv1nYeg63kW6i1IoGgx14a44nduPx1fIcUAgr332J0
RpFDk5IXyHeiNyxQkqE2wTzQZnPbKspgVwyX4YsCTl4NJINMIO69JU+Sy2YR5jz6
9zfic6kO0BFHvKrbb5qqwF7u57qcuTnuwZpaCD8foSgWqLREmJ9+EiFYro1dfJ8q
/hebmHPQoQjbRXmy4Kc39GQjmTXXpAcQ6ofxxo9b3YzrKhrYW8yvA/IJgKXyfdVG
Wu7CW72cNJhEIVu/g/q3rFbtVREe2lgSyQyA2WnjBsqCYnAjd2809lRDJRfIwFwe
oGDimrhtiVk91lhooehZvgxzhsdhHXYP1VOBo56WjRkbGaD6fkYmqNfglAH+iTxy
MEl2OpPtG15XvauJP3UE4QABnvOcHLa7fRNTEmv23v00J7WZrytnDOFV8lWU0lOq
xkL3y037z8TgucFLgB9olqUyfKGaT9YW2IBkdt5qlcRFSziNSf1NQYvkQpdyOTYW
Vomu/er3tbAR3GyJGmIZOQLYsgbLIjejpt644G2TwZfoB+0FgUHy7Cmzm7hRjw8I
SUtFH5F34s1ehlx99CUdjfYV9NkV3gR39kjzvaSusgdSB2cOk5282vctN9cd4Pud
QVoVET66ZrUYcTanQAzaY4c7PVTGKRCiPs0r9Q/cl1zpu8N1WT6YN1a2Tu4gZa1e
1WOIbp5ldmMgakGJm5onr6R+0wcqKQQd8oXD23wckMRv9RmpGtwAMPtBdIEdW2Re
KKmFIN3F6bo8BN0Pyx1JZ7RqqtRt17Mr9cDS15DAQb07wzcO9eQGN1Ldo0hqnlRa
3moqH2XWEw5zVpS4JVL544vsUaiKcc/TEwh1oko8N7bzVtppXEscxFbOLM+72dq3
Ubp0zUWrg1HACj1tno9iQkmF0EiDYXps8fZJxWtXcxjLz9etMFIrIXEYBqn8MEim
T2E45zTTkgvLOZEOaznr+mD0ZVoq0PGfNBxZ9dGZNBEkxg3Ie5tfMBPLmtA1Qh/G
/ZSUN5Z4Ksp05U0XjYj/7kWKX3t51PDEYAv+dk1cUVPML+fJXjqeo3Hp3iUzoUGh
olhL5dhFgkFq08Br383lc8FMkGtYbHi9VoG0MYIyfJAoC/SistftTjBiMwnq94Ul
6Q1aicJ5g7rNxZh0NHfevQmiV4M8AdtY2r3WAQD2+jOxNeDJUHuORh76Zv3P/21E
fKgCL8U4zf2BEnfUzaNUHxocSG2w+6CNmPpSZeqIskqy8bCEUy7FfBTRoX4IhFZD
/KeUIRQzH6BKW0u/FuAZwJxkz4IoXTV8X5TwxYqeR2EIAb1hrv9/vcZ/urmEMVLL
5KFwCOu1F7dqnfvVAP/IFiibiqDHa6CDMQiTDJr6YXtr/pzfXcUarPfHCyHEeCq3
xtgWdbBkAaarne8NdeV699JJhjQRnBDcFNV2kVl6bB369A56dkcoUX4tyCmQVIvX
R1Inx+X7PvHgTWXG3VVFRjkxXbPsm1N49vy3bk0T/mi/XPsPgXyGnhN1qyt05KYI
dhTErcjFhIEIl+nIkTN1XEkibmYuiKAPFjy2VnMQrV/kDnsz9k/fedCa1JmSF4Bv
xSeNkzxAzvo7bg+Gyp8UPG/KJIPyVPpfXAZDrl+XMSZmyJcNuB/u1hjaxu47uOnb
pvdLnxoUqjAk/yej24YCZpIrHhrO5LNciVBUdZDX6rPIUz2I3Wao/iWkgCxR1hHI
6vBTpKOiVQsNB4D77WjGr9zrYzJfEdqdta6AnquNidjWKDg+fvLkMmjNvqvfEuAS
jEz17FUlEPURiiR2sFWR3+6MTAEpx4jwPoWYh7Mxmc4H26PAkrrVA6Fs2GzWa5KS
f4Rg8Kj4/ryp2RK3eytAVBLKtl8cGkoZewEe+AAuB4XcAYI8LmQKmv1uehGJDGQ+
F73XzdOOxM30Eg537AdKOzW803FG5cbdES/wKYaI6H3+gWaseRj/TGhLJ2dwtT8q
QTPxbfh50XOrYf64OVVojgJXTQlHnB52maJC+VEAjHovvFQD4mP/i19s7/qkQR3W
h2fxrsYoHkOTc4sb4SlVk5FcWW+Ku30ZAIvFKXZO4pz+AGuevgnObHnMPa/N2N3b
uCuqitcio+Fi4jjBiZZ6tO2LOvnbhkQzeaI5FUrxZLKAPKg88TnVXxUw2tWzQYyb
ToUn2SA23THoJ80U5dQj3/xe9m0mtfNK9UVS+K/18ZNZ78dGav3GjEoEBs8LfiLm
KK7+0sGLt3FlF6o/eokyfgpJO87jllahwdP2kiL6RVe7UqIwP2Smbv+hCiiVhrV1
uifgdYyefG8L1tx45JaPpQur9tG4noxAbpn6159VS/P02s2OaDJSYzvsAks2xMKr
dbWBIqHtBpNr2KH4HQY2vk1ZxPxAG5RWm6YKR44DLS8kOWUMamIx0gYWUrA3K2Z3
XjPXS3Cqam6rLzu3FaTPNbTFpzprSzS7CjIXnKh3k1bmSsR1k7q4Rl8V/fsGjTKE
rv14xBGcWm3YTIX+/Tdvdr8HERCIcj1nyUytyv3Zn9aEKeKYaQ7o6EbfWAgFpUu3
WrKWBeBVhkkWB2BIGYoh1mjlQBmXzP1K9Iy/zBwETk2C/F2ujQ496ZYnanFWR6Sg
fp12XtvXqNxjO4MJ4N6Fj1VA8iWpFWqngUQAU2Z+kgq0GB9eZX5LCpYJCiICVg56
8zezvgVu5iHsuJ8FcHMUcOzmonr31UFl2Bh/DE6cXRwAoPQeUylIKezVAlr54bz3
FuC8Ro7NspAR3//PhJgW1s1fcxsesMI5QBsxpbGGaxCST/27dCk2+sbC+iSgmJu6
21g4Sm635g1JJdN1SFAwDK8G/BpVwBcr81cxVRJ/eSSLJNkIhY9VYNegcXqngPcN
FJLYwexhICHj7bPV+5B/+mneYulg5KjFi8S/b6uI67R2wol+eoCA8Se2IX2119mg
9Gcy76X2L60hHqcHfPs0RSE2OVNCOZrYJUroIe5pMuPqxytA5FvhXxMmkPNkT70+
kRPaomFVYNaXLU/I0NzOx3K7/Tt7dw5aS00u2rhyW+8MVt7y/qMZ4ZYyZF+54ZvY
XUrtlExrRRhkJJ5WCazsDvpFraIrTdzK/d135q3FqoU1FcluE2dWJgdt+2Tz7KAT
T0cSSIccb69Yf6VR0AodSJ06LtYAbnuVF9jSZeFHEnGRwn1HU3oXzLpsXvH3D/Cd
0YBNPUAn/9YBoB01or8DOQV10vIOU4hshk4BtnTKhingAh0AboSTg5giAjpGmqHP
6yq3smk6GjC1OCn+lGmrTn03z9CATkyE8rBDL8CpbpzO+SI+QlM6Gy8BvLg+rlc7
WvhwEWwWsuQ9dtLYv8Ou61SpFHPccOA/URfS1Q2tUSXgCHRoVUGI6q+FPd3FPgOI
bhWg8Cch9pvdWb38weY8dy6snVlbpKUl49Wz757MLbGXqgywAiw3xQCkpDKvoTLt
z5OkFrueUrc2GqPvnA5JktXMVhdIWIC2Az37pkWEoy3HiXy0TM0oCzi6AZFHtaga
9XpuKR1Atda4kn94nhaHt/B2HhF4XrP82IB+HioSTnte2FwGT9EDiKWa9wPecwcp
GZVpWQZ/4mJQ9RTW8ubTD4seCplL9/QT5l/REQBqI6RzEyYo3EQH92ipyX3WlhJa
Jwf2soAuORK0xhJ0BCZ3RqNXvKPKliOXtttQLvgUek96v0FkS1BrIx2AMdIgBX+w
duehNi9VN3UuVJbxAI4aLbQCYZe3LwlyRBwS8nbz289aOgKFSADs9bjGVhQ+r28F
GnheV5USYLIO6u2UF6Mliz7EWI9IkNlO5dvkMb5m2s3lX22pTEGuHJtJVwfBT9PG
Nb7p9uggxM0H7JpLAh0ayPcQr7G2YgjbonEeDcl5bwygSHTqihBrmRe841vtSCou
nK6mbymNRiPdKY1Ty/7zyukGp/l8PQ/dGWuAJvaO/46OFv9qbCn83NTW5EiKoFR9
SkDyoaIFHIWZ1X6Y9rkUijxh7thosD19iX+VXedkDyCftX3fkft1nra+9L+6TlG2
ohdsyCIKHEwYUAu7Q3/CZ+CHmhEUFOBL0tO8xr42q5HSFMty/4A+vo5niwERmp7/
unCFE7Ox+TipuqrBFAUQcrT4S2s/AfmS2kSHI30DU+h0VZ/+D9d13NxSIrzP88ri
L5cBFscdDpYM26j6Sa+wr9VBA3aIoKKX83RF6G2aM2ghVaAzgbuppVavFFHx4yVT
jd0Zqnb7I9LBP72/oV0sW8ztrq07NwgmSzDWDEwSDWVNCDWpbST2oJ+nVnB5dsF7
Dneu+N6zvYzskZTmKDF92P9nxyGjPNmPCpxevItQekNEiOE7j581n0kdjlB0LN/O
7KkcPLRkOo5RkhrH+aPD2yGLDfk0DL6iT3oRalwI2moaVHbouu5PCH4zXS0s2Di5
vtvFERT8EpZhGpqyxQ+qjkU01z0YUUOQ1dDDZ6bpG6/+LukhR/kvf0yHUzeVaA1X
LLEA6sF5jowgKfKC1umIXj77Aap1CpBcqcw5K9WX7/xSrovCcDMGkR77U9msyoA6
NMC/6EMDrgCKnvs4x4p62Eg14jcoccQ2ncnANwWmmkM9msch04dmbdzTJxj2k2OO
wlqnq8JyfMDg5liv3RcE+aa2MGa1eCYwSgCMw/VkZMolP6qdMS4QAov4//FoCNBr
XFW9H3dyF3LA4/DHn5EZPtmE1uThf3w8hU9I/bgWVHRnWy41SXuYrvZdOjxlnn69
m8/H7WJKyOgCRVQNGJmk09zc/Ksr1kS532KxMYk4ERbUCARaAQe/VudqSL5TqMPd
rTKpv3CL79EBeBQxm+IGjXaTnNfTXiCT4A/VvUBlvmsc9+p+U0OOkEeyy7J85RkF
sSb3kDuIS6okYbgyWMXQqficS1hTv4dwSVNOrhlobxVuwWbYKDkCutZdJMbS1RTz
cuZBzpV6LKJ4eR3wnbFKbG6EBvbFxGndIE9VStKqVjmJmQoy+ipvzOOmnv2VW4xJ
9FbY6G3cn0PTAGcn7LD1hmk8JgKQ4uTTYT1GHT13rqFOLOKr6lNW5QlbL+W94V+W
f6MFocnOLAr41DfSvK89GJoA0lnSR/HWQtNf9HjyCrSPw9C7D11lKz91mXkuqQ1/
ZBq203WjJm8WuKbXPcSxum/cxvxFV3zqzt2BhVKViHr2CXau7e1HWzIGpHW9n/+o
Ek1Nc3dmM8E1HJeMZEYpSnQlAh2EgDm5VmTFPUBKUczhb7J++faAFSQLjBVX930I
2bg51NMjG/QEieT/7mG1m6vpLfL4ukxV/9rLC1L7krIPlIYnekSdrDfuCpVLZHXv
lAZcc454JTgnpqiVjzIkDL0Kzwe8v5mDHLsmPuS2NS0hfmO4DZJzQfG4WTPH1xp1
qGFQwdeU3fheHXfGwSijMWq56E7yTAiqf6lvAkkCJwMbv+MInrgqH7rfeD+tfd7c
HzOALPH8A0EUgWtNmCjS2g+Svb4+6pn3Nh8vAWQZCV7436GfZulRGaegxspNn4qv
y7aYdyULO3fUNz2R3jGs/5/RRljViHSnOwI7YN//TMTc2M+kH0Rh1OCwaWkfIaf+
jGX8hVvy6X0slu4WhDtc2HnpZGNUOgH8L66of+4CxId+/FdMutyHBbif8KlmlIA6
qGAXYtLLRxs1t9cFIINst7ON6FRoZobly5kWuduRSejITCdUXWwzwyY5Fhyb+9Sh
2eN77uWZWUf+fanqAKZ5U51awvbMxjKc+AeQ/yGH1EKTgqfd686pqlJVTsUrIEmN
Q0BfrQOD5xAnkct6Pnrihl53WlYa1Re760KSt5VrNGy0PbCNMVuykwls3B3m9XHt
MJCbCQ9d6y2wtqwecnbYZf5xj3qXkUdmuigCRED4afI3GMMZxqnaHfnA6L04OAue
FbUqMoOFtzMqMccNy3/VAVysajiqibHtK4VpLZk/GmOq+p19m3DiLHJ6I6NFEghD
pMJo8vb/8h/M2mgb7zxsvfqZ4KQ0Pkh0Zpd7rePGfOzG2ZK93QZlMTMSGfnC8T9L
otI458Xdz9E/YiCcxFFAvddm22KgSo83pMp+pqBWVxrugTJ3pi6MMfPUf6Zvfyyj
E9RHyNbHbSHbKX+CX+mFZs19vvLJTG4lczEBZ+nBxKX1C+4BidduDwXw8hTOcnV4
lgdWdOToo/Ie69jZLRYrZtB+q8DSLldApD2TC4b0EySVEHtRnlO1jb4qpXtRRs3f
fMadswlQ7+35fwfVELtJ/qTs3fvZ6AJGEMJBMrspV9tERt6dKobXm9H9YKzGuo+N
lVHo5JCMQlN/Z+fcSELch986ARmQWam6cmv3IlET1z8Zk+fF0nLEawuISHBfD0bb
8BUU2Xe4wCQom/TXmZy0E8w0i4gUikzEazlJmEvC4TVcUBSNr3NZl+I7GMcKmaPv
HBBU3vmMtSxbdWLiypdIzoohzWBSnnzxeP/vaiMAvm+dn6Uc0OIO/vQ/9Eo2yLOr
0DBqI7ak46OAVyvltjS8LmB63fTsdNm836BDYz7zlEU6MRMJB0F+Mj/Lsm5qCC35
GP7SO0gStfWMY/9MdboYYizLkE6jvRRpvWHjkLmItiWYyK//ii5b+ZCqKLsQvUks
36MnC/Q/nsGvO79g499ablxGPhW6dgoPh8wOmw7M7wSnYYOf1hpLJcEHICHnEoj7
E9WqgT3LcFCqLA4ksPBPPiIaHPVaYgPr5ShoZV7aUTs42CtRnAJ9aRM2B4Yey+LV
Vh4ckgq1CRkyFM0Nut+ptFK/lmP1mP1U7jfEjEENwTcjsYiLmpfh0euYSSYHB+jN
2iWHuvWWOFrx5TZGOvTbRj7n0y6grUv7wMbx9RZXztlkH7E1KOXOY8IYekqPj9CQ
4GGqD5NQRUBmRA4W55KCiV/fueKUxmZ9s4wK39CvFTKFUBStiYb0JtrOhckrBZP4
oulLqgYzvNToCDJSt72HYWwH2WxPFZq09NZB1rcsmR7pg5Wmz+TS+r2premnEgDG
qZFsI+KfyXE//QrlUtUwJhhGwKY6/VNCzpIG+Br6bZZFXwAaz3e2Gks4I7yWa9tu
K0Ys2j6v1YLlPQT1UdVtRvYaHFMxM+mEXA/w1/+yKbOAD+N4JYval7Ykl0ard+01
L2D01tSgFU2Zfod0UZLLWgtS4nJ34o20NWcQ0Uak5AK3nz46X7vUqpGpfSLWT1Yo
2igYZCQVg9yIYvtpdRrNtkPLQqmy42VYmO+3R2CeIdReyAYjdfe55tkeTWs6Ju2t
zvgGrLgcVqfBepVQt4SfPP3M8EKPQPbBs/1zJFaFN5pkHZjnrM0I0qX1khBjysO4
534/RoxuX3G3dFV3dNFhScc3vOV3JQS5aHUAu4DKKy4QS0hS6bqecM6o1kDt1tEU
LRK06xq7QFHlku3km+NUbCTTdf+NpbFNdR4BRCQlSNh+kALcc7qQHcDp3ZNoW/B8
sTMLJ4thQjJTjqY0HtEjr3AmQtP3qqBNrBLxD4HQMKGvOZ9X3uI6v2DkPktrsCKo
aFxMnf8lxcbHUgajG8GCJzY/iYN5GiJVr1FsjWksFt249wxIhfJ61nQ86iqpKpyI
Qd8hPnDZM3QwS67N3Z+qTO7FhOnicGftHeZ9LdJoORZG8vvvxJ1bkXmDdTDioOvS
gOiB3AlzEyJwZmbTXgnHGbnaRe/GV7QB8ct1xi3m2EsH3lRdy2PqjR4533kjqDpE
cObX5czvu2LI7BLzfe3qym3KG06v3ZNd8RmQFLPqwTBUX5rlomqKRncOK/UOQdhk
Vxt8I/SlHRlQUIyZsOzfc9QNZjaNhLxdDjmC82KyfPSYN1HRIMuslEcnERIKHHro
3FOWFvHiN1esnGH+8VWIpDDcNkReBcRGQ2mEogFGHMYcyYLNpmdK/Ej9WL5UUggs
207jp3bO6dU7PHvNeWqCvh6Kgne+dQProGJWguE/edB+Ho/hxCn/3aWtRZS4tmyJ
1ValLrkQAb1CdexhQkP7rUt4Bbk3RLWzauSsgUK4LYUtHeiguMe2ttnn8D3Mwea9
udYyVgHQC+tZGkJGwRrWqLpU8CQHH8jWhfZNMh+QbTGewd5UhY4WdQyaBW0b6D65
cnFMU6A4rpxHfFRE9MKpFlBdDDNqve/sWgfYEyiVMH3VONLGERi7x+OQBo4YPMmC
op6UgKCwKJ9u+g4GuMyBKisDEnhVSjmtjOFhakepW5C5rjJQKdl6yMYfS0p1I7RR
rhyI9u75w63MT7iEuwoQsVkjeLWb5XR4E3TcgSnWC98Wpb6efL2xkpt5m6lYmsof
yMqQ2+j0rI4nbBDa/GdfM6PEmhId1cL/4Bwg84KUTvvGl97quWAALfIVFYYIcGiq
CY1s72gwNM2l/jkN8Rlz5UF5N8Xd3bVdOW+7WyVLsf6XRw1HjoczcYGeR5oXS8s5
+qeD/4iKUzmanNOZskx2GyqtHHuzv9Lq6l2ALSvtNkl77aplL+1Tw/mr1IIBQsTd
mSJwwKLzLKnStL4lqjRk0pJ/lFmVdiNFslXUQP8EWHrGmBwVgudfj4z4vBgM/FHy
65pU1XbP4tj8YS3059zNHJUOCHBR9JS71N+q1+dy3rbofpRx4HWx+YpJGTCdupBq
HwGtpqxAQKYt4hcVAf3v0plNpBgy2/EkXB+UYG4FBolVWf1UnDRCNB9y9/6oCGsV
nTVZaInnr1ZjorbhYT0aum4ockDbiC2GUxMUYJTPZMUwBoabtRrB0c0P3zIOyEuI
4SjASL3Jg11rDocvK/9YzeY6Qug4xNv3KQMjFzryTtv4VvE6A8QRFNeef5erdf2G
dumRN+JDzXx0fToY55ThPP4k0KnBCfbJrc57F6s7Vta0k7P6yN8ZEPwd4rQtflmr
9+N1KGXRkmWNB6TBXg6HpdvSLuSb7ciT+Uu4dZq7MANJcGI5bnxWHEJXzDp8QAqA
GPHLpKQPty6dAbUVre5RSnjc3YO8MZi6zb3iqdRup7C8zRfqZSPE5c7iUPu6Up9d
0Tm39QHGxMRtH/4B+MB5BoJXOjz93mY+KTJltACQZtWVzBTummG9Yigck7cncV1y
XshlTVsIoVof/eBg4D/XrxKPc+/6CGsbcacyfIBuYya2fVQuXb8bijyKjKrtbd5U
Zraydmjy3nstkW2TR6NiISVY8hWqRx7ok5hFASXKEqT6eZeedlUXfmpPvEB2qtt7
PymQb2+9LXtsRakyEmMlMrz52dbMYh/zMfz5OmY/FG1BiRrfEIQuXUnQa/yJSiLj
frencdhVlvkwDw8kp9Q/i7X6MdUagMgWw0LitMHwrG/Jxrq+YEKWYVD8iddvyQDs
TcH6P8ER/UgB+1ahw9iMhEsCpAcU7XZ+NITvBnatX19eRGjsLQTRDuamNwS6Gmh2
/Y6JmxIXzGHbbMUJczIlUgapeZYoQ/ADjW2QJaBFvwppcKjepOnpN2Q0NLPOlK+1
5moe6S4AYrr0PsvXDdH4cG8uwaOlpJlwLyaaChqrkEERcmuREkv0OHZW74tg9IFI
0FgFRhhm9kJpzhCH71Qh1ch0aK+Gg0Ts0AadTiQWGxedDOHIhyfX6SmrnOE/iS4X
LsiCmXz5WeSMdWomxR4BcwGgGp1flMWMdhfHPxh3+1gwytguSBjxnzjO+OaKjTik
et93tlF6OXOiHwRX+6rGNr0VlZ4Xroi65ObGbPQT/p8J43govo8o+L+818uU3ICO
SkF6Sp5p8Dku/QbfQMjg8/2wmhul6ndh2bBqCwBqbrbE3d5DjvfdhX0KD/rWzMZP
4WMqPz56pNSRtArONniMPsxht68r884WJ0aqUSvBzs8+rJQTGpm6JOHZRuoGVjAQ
R8zIfxbI9lBX0IeOdGp1oOQRvFDc99Jc65gzZz6E5m6h6BW0s6rqABikRdoSK9Rd
+xL2KxUkNd9R4LLycb7GWL/SgprhiwfcM3idOKPMHcnTq8H0QY24YS8YKPRyUF0P
oU2OnR/QE9VUdqgb4jnIHmEumyP7RdfdRVW7zKn58gUaxx3dHx+PHeE622ftKH8+
fYISg+YfoA8s8fMMEeXDfm3yPCcRnkhBUlggbwNbrpPvC1+k0DToMpKQqXMndDho
reTqYbn05Dl2V50xxIAGM2QMjZDlAUKFzW8CT/L0uZ0oBJtA57ZmOaPiLfuVZMS/
dg6MSyYf101NfZ313j02ond1Kfr49atUxVAPqyul5j0rANtFezlIX5m5uJTj02uM
aEkDPb+w4xWIYgXl/BeABR1YvanSOrbOZbMfYArU4e6EZ1UmbPIhIi1rXefa2lxh
KDZL022f9XxTMCNDZjJ3w619ABHRQwlcKm4JCc/d3taGkCYN1fcHJ7e0cx7V912g
s7rd0wgKi2lzmegWRRmwXrZuGAqTOAuw4ov/AoQCUCAiUEdRpIFi5g/reQ2frjHD
LIsIPIDODHcQQ9v1o1zYEwxrxMwmhlRXStWjkrk0fg5+DEoVoddDmFcQFLUbia2M
pt8Fz9aZWJOOtrgMDfvB1NJCYdsEHFSx1CWDEUX3YPY9zRNFtNu4ChD2NVYPwYQk
GPN4e5uwlYQVf+sZ5k2G2IzUGG5SKyhO9n4XWId7iEqlPiN7m4NvRht/GvPV+gjr
ndfQWyc5qlmSAJVN1z8GwNYmdk1qV4VHke6gI2bR6qzvWwopM+HOw9P4QF4eAeqs
zYe9Zmj840TgVnhwIpijXYJjhfGcGV1qC2erEQ3oiKqMrW1GmS789VKEWmcPYD3y
TAJB5M0MiMp3sGfiKycUHNYhs0xIA14k4Ovmy6U/LoiScNxHcBZp2kPCCmYRwm3j
8fnaOEVozLJp/VyLMRBRwVhOuo4+xfSoYgH80zYnicUINaV/DCWRx1ZU+IQw8X1r
+my5AHFse0TFWJ5YWHvnW4Rxj9JwCvHUxrZ+tDm6keovw66spMYYBZEyh6/BwqkQ
HPYGAEolV5DahGLEUElT+zM1vyqrzNlgeQbeBODkeuPxnhobftJjSb1kT6pikrX7
3OkGqnz8uNX6+LYwWZvdpe9/NKrCxWwSd8MYlP4N8k9vVneVGqvPa6RvF2nxuitV
dCGiwrAvIn2cu+EoGy9dUwfx4tFMEas/HzjHVKC71BIXfRuU70Tg3pNoK++eugNi
idB+aC/T1AVBcLm3XSBfvFHlarNrjYt/oX5xWSHk8U2JeszwzgwojkIYfdgeyBYT
pEJeVKKe299v/Dngr9H0H0l5yYYhI8SLD4hmUe877Ls/ZHeVHSI39KQJcmYUshVh
UUwX1yaagUrb+w7XuvFkgD8Whd2n5rX90vNos/sYHtotvpvqgZ88ahdHVbJzjzM3
0jK9hrNZa5qpCIRUKDuqqrCD5lduZ/3qYzWmI1XXELJSaEy+2n+EOnxl4I43xUTH
UppktO9eK1QcofGvN23rmKNZfUsef5Z6TAK1YqQEroiK89Bc4leXOvRealXTOTrx
NPA6gSA9hKLH5ietLX18QUDKtF50Gn4OXSRopBgexCEW25MA+FvescE+xVn7xptA
r/WWXiBKn4ufcJ4XIiL+Fe/v8KOPyAbzpke17yVX87Q8h2Sz7OWAYQA7xyxQcxQm
bLYa9ivf8xJXk13xFMQgrYww9aNgj8XClyPr6llduHdnd2wdZOqLkWGTtF4ShOeI
QQ8JEh1CHCYJNPm27qSFKQpnxEkt/ARnbP9o117NZJ+WPulC1ndZioZKNmHmRe/a
QGWl60LO+OiapbdhSMYPm4ch2/GKhcZbwsnbYfMUNpc8DpBOFVqNlQkLQObTUUPb
4l39zVGuc0mNDqvLyVTR+tMhnByRc1PrtuL8QPtUFzQiQnjaGuCo/8R0NFiElOn5
+DF8GfPsx8qkG6Qz8BzqnHB/2O1G2P5SbDy0sxUJfQthPsdEJRL1tjtVeUz6bWe/
AqMzGY+FPRREdyvGhAcQFKsbC78lq1P+z4RuISRn+j53NwVDDE6LZ52fZHyFMIGY
Jw6TsnnjnQUWy7QrKW40QbD+7fL1gwmayI66JIBzOeISibTJw6/HHmf+2davktWw
0EU2TVMt1k2ANKKQ52OuzQaVugL3gHObizMOuWjJ1VEAF48L9GhxCZeShMnZkXcM
xXSIpVaY8I46E8h/lIvQ+nXPTaqZr226PnsXfr0FdifU/RmzNr8W+d+uMt8vwJbV
7dZKOFEp2lXB2GrNnfRvIw9aqOZ+N9Uf1Uq1QAEJ+5mx43BrcULzpFH4xr69mZep
oF1uR4FAKylFbOC84mwb4nsFad+67WhP0t1nIyEFxvayoviGWZOZa2HKEcHLKOg0
cVTyVmYyPgyaavv3nirHIhWQkJmiwaa/fEGrjHIFcJW6zMHLgN+x4XkDOjiGqpLV
o77gS53YTVJtcQu6Sp3BDhDgeqR4XV6yRUNFLQwiuBSbIogVVK6Vtaie5sUlNXVP
5/fNBiFdmM7oQQmiJ4r1qZJg8wSv943cRQn6fj6METtup66bxEKGCmMtgK70T/NZ
Gvvn426smnylTOl2cdxFwojwnpH4dMAGK0mRe2VF3yF9Zub6yaYcrM7emVO2CTvB
C3Kp1RPZlAgVRqqvHeso996gGlFSRmXM9V5aqAKY7rvKPauGSyhHzm8QiA9HwWKc
tPRQxT0Rcxce8Urbi6bUizAFjh8/R+wVbqlZwgXsnn3Gmc0XKOa/Bs3Obhnk+cJt
Y9gxlsQw9q5b6XU2F8mJWNIY6B3p/nDNYqkhc6JKBE7yZNPDnTLicKghNNNSIgtf
6Lho973KR/RIN6whJ9z+pmMbmFD/sPm3HethMeqqlfoplzbZss8yoY65t8uM5oD9
wrYvycZc4X5+ZEUeDHe/7q9zaoV3/nAx8pOovwEqJouIB3QRIN/TfznPF/l2BxYR
UiVdIjPeiyBuNws/25UAXNk8VQf75bUGUjnOvPmnWHOahXQsnNWzadjQOR8IGmGn
et3xnmQIa4oHMTVU714UDGQ0/1FdLaA9Z1uwlDjhdTETk3QGUEvvTzN0r2ZP4i5L
/yjP8pQOf1W8PWu/IQbRN59LAznQNtM/G099AEIEi8dAAjATVLDVZTWY+rfy/mfZ
RM6S9J70PZ9c2tWOyNCWLaTxoza/BlfyRABNW+YOxN2qrOeiFRla/ZS6sSD5SQd1
0nIXqbgx23YPmJyjpe01vIK2f+vo3JzHv3e1LyBApWjZz5UsM9lMgwIZIlsw86AC
pZO+YKDfelEVm3bpeRmVqbAtgbUTijHQv1cukTKoY1V1kYBPbswO2MYVxnMOxAej
6yjVYh9QGvzNRP3ffRo2hGWER7/cBYpjPqosdhlUQPhTSH930Bry6qKHPZMc8u6/
oyx6x6UaXDG3yaq00JawFa4KMGf4xgEwzaHK5pCGAAOAr+Y+YpPrr9TuvPclrqdm
VgP9a0E60yTaWCqbuAblns2vDq6u+UhLmjldTcXaTLTEvHWm8HOv0k8hsNlWR1zy
cAWwP7Wl7y7wP5I+q7ixbol01c5h5njIGzrTho6P/lON4Z4m87TnLwrepsIh1pJ3
S+dkB7SLeGyJp3blHGtng7TLp3lC0kAaw09HtXMd9p9gGks9iezRqSbG2zISdpkR
7jY80OTqIKrr/m0lSYs4Ektocich7xuVXg0jLoLZ1uuKKEfTG0TfrMvDp+F7hVYh
pn5vR3CzpiV5ECre8zIRlA3jR/98MzJ0D/zW1T0VMCuVH+91tUKlTwIpz2zAZnrB
n/9M+enkvLCHulmrrdV0C/OVftJoAMYo2uGtXOQRTgwxihWjfuVv1I4V1B0a7rCe
GCDXV1LXnHENB0GQ7EEfjBOuFCrQzZi8dzmLvBoFpwea+Km53XxOgRAmIwoEuWpb
iC2FDDEZU425slsksc/loAEOvryVpM64M/1C6J+fJFQTwgk2kpWQDvsH/1KjYJ3d
uki1JgZaP3CwV+MbWOD/q2sT4q8s7P7Ub4J6GL3O0YCLUXma2cZ/IClZC9r/uuMg
YJJgtUa1Dmt6CYsws75vYj7an1Oi6JXnGBpZqVec/EyIsZqWnqKEBO34s/5O/yVA
lh9cBJPLMc8ycLh2K1J6T4s68P+NV/4JDiI7oab3Yrzpjg5tgu9cejY5u66SlHv2
bXTgbNktgZh7aXlqJXCw7dnKcmDKR0sCnbVrlgaCiED+8OIyJ0kAKDL+36XIOCio
QqV19VMpDKHGH4qGGq9M62lD9L/sCXCW16SKF+qpBX+lOtfTyw7BSlGVIRpOoYNI
usAl+DnBV5t0Afs/lZXeACm9CxkQIzaj2oxcnwBPe0VWyXgoWTk1S5gjnySvc3Da
Vh8ulsQK+LIyqrVsvkRd3uSRRrU2DjU2x7Lc8kT4sBmLTxYyjIofUQOtvQ+U/8gR
9ar/GrDhFftXZZtBGY5fLxsq76uQqjHUmtYo28rUpsqv7MAWEc1ICd6hiNqcq1PR
1yVDDfj4HLuYZU4e/SFSegabnR63DqPJKnMFB0NrOWzChpaNnVnN7wLfLgURObqG
WvAVP7gGQfbxNNMWi/lwghfxb4p+yqeLi83T8kK4IRVVL0VooALzCZDzStRbCTdp
A4URQf0SfP6VbJmeABDiUabRQEPEOkjPpZvsINID/ux07QMtwibgSB+/Y8t3BA60
MaQtaVuKTKNbr3Jr3toESWheciTSPjblWcrKkq8CDCcAXNucYExD8WIpPTkMjdBB
ILIX+yr4b/OUI3dZiFcU9ibMWbHQl+BnDXx5IBn5kHmY+EsmX9bkfop/lG2ZmcVL
PYb1Ve80p44sdbqyt0bia8yJkCWEyQq82/3/WPn/IoXkjKt2gkia9HH1rbiCjXIN
O6UFpNNBI1ulzeZQap4okDlfy2i35ywS0qTm1Nyse5GjNPtovyu/AliEoQUKYf2S
g+gTBUvq7HL3AAOFC3Ey3DJSV4jt9oBlstcWl9eTWuD+qOkpE5gVIpm72i3f1PIZ
rYdNLIaQ2ltwfjO8Roxw4kmLDv9wCWuEQLA4Hz2ZY/q+Hq63DcAz4wm18t8Em5m9
Os6ELOV6mx8efFpMbs+YKIYDWBz2LvO3hEsVs9tm0+qOpxl44UzcKahSuvFYEE/x
BGpisvmAdb1MlY/xoTglfeJAYxi2jbKyKLguvX474bKvPHVqe5E6kSqoN3z3gPaq
c6WehQBYefNgY7YWgCn4wu4GNQaAPHF7++g8/2aV80qaXHTEkp30nG2wXzuaNU3v
VhrtJAYNemEuE+GGwgMblWnFP0f28rJCnj2oz5tJFXoK99YtapmUelciwWevv1G/
9Hp+VwSPAHyzF6tRGnLivqKuSodEUD4KI9qfNQQ1+92VXk/RLsz8MgmoDRlJ3L8H
I8ihLnjIKJ6m5m+rYtqyApBSctMS+uEcJ0XY02YxvcNVm1cLJOpa1BKRFTixal7K
aprm/JwNMJPn466dpqq2oFgx505d2gIQN5vg7hTAVR3YG21jANlTRG7G9Y46r2Jl
+L7xfzOUvAgnI3Ch+HUOcQaGzck10u3jOyKyqs0wGVIWieTPgVdC1Z2/+A3T1Wlx
in5BVNU4gGb9Z5RtpjOM1WCXjdPajFP+/uOYN2l1dw737/QLG2Zrinw+vuFVI74p
mJ3+D8AM5SuUjlY/bubdJyv76y0VTXDjdspUyV7iULpBXLvnXTUCY4lNXSLDvaZf
Gpr3syeZSFj/8lw9CmqW1m18q+L9Ms1eLRZD50dtYITcjIYVta+PqIf9ObgorDEW
+FU+SFAgUc2Pci7tC1pQ7lj7iG6EAZCTG/S4W3Uy1B1otm7IDxzTSaO3HHDbO9hG
zSFS7kUux7CNbh5FmGjD4mESFTBx6i6KH82PI4YqXFyJfbuoqmIMKws00sYg8AZy
3qjudehoiYqCu6CTYXoJnT8C5DZOAplHUWa5r5hZZB59aB9wUZhzQ41U3C4xFhdX
AtCG/6lFvtF9EHOWJLGbKL8p40Et9UIxqgrx6jRV8zoHG87PQejADIzUitDMhJD0
U3Nrvx+lAykyRHIAVCeYX1IkRpBxMgnaDENBvMyf/uI0HZmUiiBzFf0p3SkKwtim
K2ZVZg9XabEvDNn3yrqy2otsmqaZ50soiwKVNq1QbV5synMFsNYXiTaH1UgN7xOP
1G0gJXM0HOjM13X1HIa3wKaSUtBrJAZO0vj4Lkx+KRTR+tIhldDf2MCB4rlMk7/U
Cyfh/QEko6RkwKhldFBVWnV/sCreUejHIrgFJwMsEjtH+SaQJA1Up7ahIuvpm68j
lFH06XNt3CmBYajrATPgacOQ8xKlI9LkBUKuOP/ueBAJsuQhnK8bIQnrBWuP6inS
5ZcUeHWuxRENEzp2SV4ZkGRpBEJIJArd3jaGyuA0NmiMl6jzECLAz6iWlcAC0J08
Z7RHbUJrbym5GBJP365VNfdgXNW5VVXi7Scfv7GCXJux9UVhONHWfDzw1JvB7Ad6
Oxxt4t9tF50BfUw4DO7Zyxk2P7i7DAgzRM4u1jCLOTqkUzwFPorlycCMKXB63DYc
mM5HujEodz+OI9IK9yM3a4+M/uxNnu+jS0H9upeacwbi08KhdXqNCz3cc3qPTbmO
aApgl3482OGmKYPYfFVihdI3hLgiltvA4dQGLR2xPPl3xneAYndWq0Klo61JnWMg
MySQq4pI506hvw6r9v6hmnrZ8TKWie3qYxR8xgSzJZ4EVtN/BCO4/5jyPAaEOuJx
E4gS96KtjHUI8VKFIZ/z8VICgsfEzYUWwYRz/u2luSDZ/A7cY7ZLzOgKMFZMndeh
KJPVOaF2U72poezcVL/VLR/XCO0PBXTf9O63PXyNHQe+ElOjdrZPpO51HHZ9o111
OigVBnwgAs27blaTvlapeCWqmxpS/IzmL0XuTg31uogI4uNjnW9+5FhFWZIl435W
3i/VeItBIsvmwCbGWdkwQyS/gIX7mgA4TREVIq+ASHdDuf72cr7810ZLi5uc0cs6
jVyNMUgwgoOiBH+gMaq+PJTWjni+RUdBTfAJPWTYBYCRavmpnJrvdC1l+4T+oYjF
qATsgmO8oddzrDee7YQ6A9/URIEXj6hn+X9brkGGtPOIWLh4DGb5z755vOrZmZEN
DO4+NkZsh5rawP3NKt7YyeVGjLMTvS3tGhMgrxzvSWyg91YzNsob5rkJSJagY3Zl
g9VDz7Vgel5UZOMQ4VRx8grF7Rgb4HBPT8JX3DdkXlxKgiXbfT8ZTIX3jywz9hGE
VMgLSwoVK4k1kuR2roiqhawRphkKlow90/xDb0apj1XVTJKEO+Af2fWftsoR4Q8M
x/+q7qgyfjfUxhHWyRjz+Zx7Tl+w+W6Opq2cPOl4f8yzZL6F0yz8yuh6oZi0y6tc
7wV8PCTNgXJGaBVGflNTJcMNsixBzfTyDP3BMwzAkI5tiV+U+99KNHKebzOdEKGw
+GMBZmGwgJgXLHj5Lj9Ic9S6rQRjE+6YIa8IxPABVLRo6TELlGO5rD03zgFASGii
rgMiUT3X3eCr80ux7TjXEdQ3xcDdTvtI4NlusAqMlX3C+a7ugfE9z+jAoZ0zU1lD
EcvM+H+Aih8nntJybjVQFemploq+bZqem62JaQA9qPd+8mu5bYKkskhyq+oFyzti
PU/25dyAW4npN49ZK7+mHcCuXN8MEhq4y6x0loM7e8diHOaqgNE4GpX25QKS0Fxt
47vKKkdviGawjg8YNlLUuKk6+cEqTybDk2SXshWsAnd+Ntajrzj0FphinTYYDwNj
lZcAVT+Z1jfwnX6D9GWesRooM+YLWwgagbz08RYGFPpFR07fOpdyDB90qzsdnIiI
Bw2OV+vlHtQLggzJNacmBUw4c1hXjOUUqEqC57jDglCu+j2KkZPGTJelR8hLHRVi
lUfR04gfN1ht8qdZQPKP9X6zi4gjSnmx93vllI6pMgwwqxD2XhwqhR2X/GJOjQjH
Hc8jbdT1eBxWeIlsnxyetg8hgzZ5Q62NYh5QMQRg0hcs2V483iDuXW2p/SqpTsNt
8OJ819kPqgTmHemVAtHuPxcyM/2lMVE4JtQjUSxDV9JODXHuskbiPbgaoPP4p4Lo
/l+Tu94yA0usAMsTvuP3Eion544pjk+ipIRMkStrHqE6ZTy4afcN1Kat7LuDa8GL
/RwS8xWNcWgZB0UU4SDS8d08om2Y5izN6Op9AP+/bc5qruj4+hJXF35ohTsNCS8E
rZ02ku9fiSpRTM2187eOAe9+xOV41+OzzNBnDhb0v0/hn7PmYYxrUtpB0/rNKf1l
WY2Ba7Y0VoID1cGLZr+2H6WNAln7kqhNsho+NO/IiqaJqL6gjKyTeK03HrNcbcMt
mcVRA/VgVSw95KpZehMuwsfmV2DCreu+7K8nA2PVRyb/gJ6+urTKbwTqjN5wciOQ
9xfgxLCSaPvKF9F5UlTf2JMtX425js+EjZB0fJE1YFOAQOcG+rjw8t0elxrs3fJE
eZ+BfbXE1II4y/nMfoWDCRBSZljeDwO6b4NcbJv9ovZ1Dw8FslBqFZquGUVbe7II
DYvgSie06pauVPYgkr/Yi9Yguws8fVNoYd/E0coRmyJ1MVNu/t2wCDj2GRuLgaeT
PoNFPy/qZ0LId8ITmFH3red1QmFqCWKPa0XpSz07EseEo1IMBzJVzC29XSP+0yGe
OlRjtq0JovAt+8mcxeP1+REFoF3FyDNex2ulgOrqfn3LZLMfYMJam6gX6qFWs8xF
iAZ/ENH1LAY3D3OELo33bCLWwgW/vDAVvTWYItg3ueZH0mzPjkE5brfinuNtRdjk
HMHQeUYVwz2NCBi9tWMmnNiHlODvQnEJ6WrLY1OxG8lkAdC5QNbSEsiTMPGSkTZM
axFC18BC1hU+PG5ABwWZdusjgk0KRK3UC62ACoxWiyW8XX65B3L+Zk15lhALMzBX
Ii9u3NgTXkVREHouOtVCrOESxsj3b9DBE8tAadtmgPB1N7cGaJ7EL4Bep6KmDBuU
fkvb15+YcTB0AIQggR2ARmb17i/JJ/TTKud9TpiA0qeWfgcnT9N+DAJFUIefF81X
IHGDBhCibBYYi2/JSgH19Yjz1ULswuVJLxFs7CSrEJBd5UOx3ShFovHEB/YxANwg
/sz3msbAL4C6LnfyOOljwr8XDY2O1JLUQSF+pJUYQ47bqxBn2RbAhF7njH8/VGjB
CBJ+C1CUfsNW1a42mKo7JUWLcHbhypZTbvyTqd5sFnNg/Oco0qk0R96zoHTD4NWA
GQruZaFPRisKiSyjW9SEc2iU3Tec9ka2HlfiAwcDYW7ongU4OkLA8e4lSvXdWeS5
jmRLbnepSKkdb9d/H1kccX4J/XIf+6o/ujA7e+n14vxjnyQ5+6yuGDJH0MQCtdNu
+Z1v7AxKoxObM2b3ZGrzmmApnzHjBX9rxkd9E3Qjn4M670gy8xrNdiFIMCmmtIwT
euPiyZ6dKRSNyUW0rw8FYY4DNZrZKO3Gxi1a7XxZGxkX31mVYcacapqJodDhN+EQ
s3kV8lXhnMwElNIgRzf3ZyHcXR6K8EmqoPMLazfRU6sGpjrJWvpubiOanahQE0uL
VfL2HYGbMaDpIc9NjPPvvILSyAFrWYp5H3whcaOUY1PxLBFQbI5oBjIrW7eIUYDy
xcXY62qtk3XFittiroRq67eDxHv3RLYabTxW2Z4sifY/kgi2fKy+yvwGdc5jNmo6
xjsO6G447QaACf+ghhURYV3n2SpR3/EsSIgHu1YIN8MyGLwp3pAmThdz2Y7AsDel
GW1o9XmxLwe3/0llacy4uswsAfqpDngw+GMSGXvlCKR76/ZgIb+4AL2dLxLm/AdR
5ABFjb9TumEu5yEYBe7BIH1lXYhPjK2kmoL5dVlldB0/7yM8NS4B935AGgYCvPju
AwCdNZFnQP7NyGlPtPdQ3kNYCBEK42YBYBlmmL5v62t9XU0SWdLcfB86PTXt2/mT
nQ6eAj1XWJTE8iP8uyyECFTOUX00NjOW3Uw8HrxPkMKT6pPRcvCKi7Hu+Z/h0ltR
MYpzEUNNA86OS8jWphIrOCRpxvjPcUPHpQvBlpXi+gre5AJ05UqKERISeDVmkGBZ
wIX0c8ET/gZT6wi/ZDXtbxhD1QtTHfu4G5dUhVkgKFCBJMBvn5GDQr8qqqlUPCi1
SiHJwEtx47+Am2L8Kp+lhlCSR9OnDJB31Gowl5YHlvxzQhU5LCailc/3MUINZYt7
3WGnFBMMZ2xTPjGL6PBbyQxClJxfRyGbq9I+qgUWt3P7FPaR+WgMpcTrDExn3mVl
fHJWUDO88q1vHAQrJ+eziVVKls73WDD039wycGc+kST/nRIsuaDrxO1mwPCe5a9G
VKHfN/Du51qUn6JdKumk2yHKTVPAnztcz18CFhZvvxa9nM/N5Ci94zxLWW2Qa71V
aZJpnWEs3bB1Vre6SZ5nmDFtNA0GhtNPa5J/mQkf99WkJROD/mHtngqSAfFbv0v/
jK2yVEyTD65y1IXKxk0SAk5kU5bUMn4ox99m8Bu/tOeN7TkTdYQYlBG6YuL3KYOq
fDAjg/2mzzGlzVSRDH0NcPUQ7/IuCY/4p7VEdHhX9TGeHS97hnvlGkwqEhxheQ+a
0UUDh+aOR/yhCHRVQTh0lFkiHyfTGOl54pKoiY621bd6vSYzPkTcOxXC54/ltx8E
sewI++l80nxoj6vGvtaKE+JNlBWmtBE6ZcgixNchh+3iIwb5xPkZ4FFlTtEtyZHu
Jx9TyjJe27/7TjOlDu6Q3LHDMgCR5VAQ6TDPOQPVithQ3Pbr2+fZvKpRUyWJk5eQ
t9L2qSLVRpnKIEdNYY95Q8dL95jUQEAA9mm0+298Wao9C8jfGjLZP5lxv+zTIkN/
2WHSjg4oAg6GeYOix6E8j1cgChCGX80w7pjSxKuPpX5PzLarwq0vTiQSsvG+/JVL
HL+AMprNst/naLqL/Pytw+SHZCtu+LV+Tx6K1195dMYEapDQJAKhffEU42BJdphT
jK39KzUUSopaRisf6XukP7RaJW548Y4JXg6YoXJsHvqR394DfnMARhCvoJ6+MtlT
Z3W0NSUBdeedHzAVd2oDU9B1aqjUNFdTAm+QWdy5h7NE0jUC0Q7VopO2V2EJCZP6
xwELOiVttlm7Q7QwhMFvLKcJdMsgPk4Lkgf5sH+93xF9vBcssWT1359aKzIIhuF5
w7PURaXW/3XXHGuUzgGL7k3HEMRdsPKjdvTD+h9828cGXwTHINzTUoGcCjsZg7bi
Jv8RrbrKZbq5r7I6C4pEe2x5hYE+GA8kHwlCRDVRbYdxO7TTCEJVqozxqHcbpoYF
0LbPwaOtv5hpaPeu3dGpG10VF2kB1kluMpp7h96kEtr6AN4+ZVHPJz16xkoU7tKR
jjUGng4TcsjDuNcjuUdPi++U18I7iilIcqFVVsTyV7HtHb4WiwEYqowQaIOU7BQk
wFr9rEkB6OIX7ddexPm4X9TFG5JYRKsqO1b51V+6KUOIGSBu2zZSIOeUYiVL/U9y
l3KvTWWiMXj+oplmfNkT7Aft3n306PB+ay3wN3nAs3m6aANu/OjbfOa3mib8h8XP
G6O9zXoKa83Gy8c67oeth6dGVjO4WxVo7s3QkRUnpiMMWY9bUyEWRtn4NfrvE/UR
mM8KhjeWDvNYdKkrxWuTUyfY8ve+C3L4Rfg0D5IhQYVSVzMI2MEa9omX7++SbGu9
wj2Ewn88p3CBo6RTOjXk8RCzoNzfsoch9z1MaQKt56WaHii1FipzriaiAr/bAW7s
siKzfbrlbjLEfZwx+MRyNGX0ATxgZLsY3t/oHID/OJbVmJAsbOOajdngEHZxBsnO
IYAqoWAh2kjqBJhAOUeu9vbeATZqdvlwnh4Mk2MNAx2cOGRnGs/9W5WoQtBOPEJr
Q21fy4Ky7XOpopPHRAsjc8HCQrB42/UoB/jgbJiKzFjoqlAYFlOkKh0ISVNkq10l
2g9wS1vz4JEc5cllTQt0ygaZ/AkklCTLOIDMcoaNbuXrMA19GkvPOOdWTd3+VOK5
mUUqjUay6/NijTGMdhDgHN0voY1a0MiWtIHkN3t689x0Va6UXc+iTeswCx21W3NE
42FavrAS0UP2CGdsT0W0puVEVTcQygFLIhZnG0CfvWzNHnG0xvNBYDC5JmX7YSSj
YXrBuRNDCCZ2fJfE2APvLZtkK1Z59JgcJsXORgrHIGXVTXsdYrKcKIX6lD9Y3cht
30cZ2v8XHPs0EHMkCR4nRH0fk5Mha62k6aDwaNt9Jx7t6eU+m4d3RrWFz0aGhzTN
bFY5HCndT2dqHhb+8KGyflcEQOzIDkkovWs+c/5O4YPE5Wn0I4vTSgq4L6rQxJT2
M7s07ZmPeOxIouQ3Vb4By3ZC3bNLPLiAXhuv9aLGvDO9AEYq3KnUchOIku6b+CXX
OgTLZWaKmuTr1rDxE3+ZzqSUaUGN1AWSEhitjTSS+1Gg+tvfncp2hkC9WXoE0GX+
6RGBOUQAFbku6mC8Zy2wgIQREgpxxfvIoXdlYWYS8+N+ac91y2yVk2hC34F+n2+N
wOTlsxijoEQA0iWS2Vq0m86IHLJMJQrULiFeP9tLA0+ShyU/jMsnxTo815s24Iuz
jFRPtyE6AKrW4QP5o6M218E1mNBmj0PPD5l+rV6xidLXYR/SQ/UFjn+ZoPnw7viG
ERSiGVSR5kux4655rPS0VvuTlD2BW+5o1q+Pq7+gcx8BJsupwc1jyFw5e5G/9XoU
+A1n3D7qOIOjhkb6uphotBCYMhDmsSrjBYWmOqpyJNONCYJNo8/5/i9xMIlq793/
cqTiPFb8OY5x2cfO93kpKpKTjyJvWR5o1DpSQD+Y24aK3UJWRhlQW+HmId0uOWzN
mDTbSs2/DIQAMY6FbvPtAyYn29q7BY0BESVBNmxxsmt6c+FAqKFfx90tAmZ9sHCp
ygoBCALBQhdBhLtD6vvoKsB6JPZVIv1PylRKy9del59TQM/nkvXI/mUa36Cz5A+6
5WrW9CQSlNJpQBhNo/t3ueVaV8YjVqWWEjYhvprmYNLCopirsiDpvNhyt4mE0dWd
MuWHcpxEWvLFCiHXJBSafPCUFMOiNgobjaZoiPO2dICAIe3T8ERZAs5H+hzTdGsO
eWYXYT/lkhc3HjXXd6QWAtpWTk3aaBvCrYFYy7ZGb8CdL6+SP8cWxaaW3XzdM0+o
a3S/YiMKDs1wd3hiql8j8IEAKvM+e5wFqEH3OJqN0Owu7O1nP8Fl4JuAu8Jg0NUG
EEsHWeQKrTCJyDLpy5nTa4+ijh+E2ADTKMDOddI0UAXb71PQBd8wgCZa1hQz6Om+
YV8ObQBj2IAXLiwKvvCzf+uh1A0yNACmzbEMXreIxGmsc6kYp+SM9iZwGaSpb3vi
l4diohzNKoLFf9t9AYhzLbmQpgMRbFBiraSI8tC8N/c0tiA0amJpEUUGQBVeKmyO
nPZ6waCRYzfCrl9ouEEY8DCDNnav+bI6TZ5uOQh/Aytws9CC7CVU4N3V45lHn6ES
1uyp4XXbCHlpzUp9b2ZOC2fjNwZad6tT812R3EtO1doaB/0VynOji/GpizjnY2aM
4c9AlvwwcE3fkspKbmeNzxrKrFxZKdnpjqwtz0DefaA5ebgKIIqFIpPZ1xGGa+Vo
CaqD/O520obZbsbCJ3rX7kOPQwndPF2udv5taVfWkRgjwx3GFqy+4i0g7OLpjo5n
7CDdlAbsDmdFkp112xtDvkdB9nP+Dj3nhkVVirVOeGDjbA6MVWIdd1OrUOEcUquh
Wr+JhuLwHJt6YWAXVt2t5YWwentUnmZ49tcnzY5rRi2EqQuoWsGf8K4lqWwhWb2f
IF78IqZMO+GlRnBL5dMidVSN37oDRFLxL2EMhbAizjpoJJ1GUml96UiwAJD8+3u9
kJ7/j/Rsv7tz2xFIuEKhK0fmFJgP86uyQQUxByWKUPmSBuLzpCA1UVIzPMVdGps+
S2+4gz0GXKZV58CjfHUEyad71a1yRgFiCNPUFafadEyAfiKn8zy6sR7nJZlhte8U
8iZyja4P9Gv91gK1e4gP4ITS6oHgicUxvFzLBgaA85L1/zDWUigkjt/ByoGmy5+X
5xdj6E+r0/C4ud9CNMvaiyOqe9ozIFOvLXLrfH1jKJxmlNGPuhRJi5FjcYvpcRkJ
GePDJap5XtQim8M0WINy4WhDx3CZkCZ167h8Nm1arQTjp2am2PdO3r212io1bjBt
Yewl5XNFoLo91FqMQZD4mXeP5FCmp3Qk3S/1I3gDLopX2qRZbjk4e3OVxD3PgNKe
PF/ys4NXJ5zbCFtvWzJRRgWuzWeSd901yXsxbYBU0PXJN60Ht7dvrxInY2ikmTZZ
wgWYsD3OKy0X5RWx/bBqj7s49K9Cy4MKddPAoJtMiwdWTKr9aAdRlqJYcazISfTo
npzVLr6g2J8aMRJ5u9F6Xw1kEbU4+3wd9ZIwadm0i8v7bM/YT5QE/i+YDl0Km/6M
WBcHJfbl444Sz4gfDlj339LY+5930hUm2UZC84T8Sv85irILixWlwMU0SfzU3zod
iKgDhvx7EWPppiFa23mH7SNj9xg/9OJ6nSn2Hr37vxlLuVv1pXDunTx7YJCH0898
5B8x1MmE4cs7vAiquJHc8OQ8cOtgPaEuhVofa0NWHVAsaAogJiZ4rflNpQ+0cyXV
XIubrjQzkgvYFKy1H5Ya/z9lPZPtlRazx1MWtiKaTqx7k/4nk62IuPN4zzq5c27P
l6MH+77QQRqCtUu+ShDjqUe4hsf+0aJ1l0kuDCFTRdXRO9vQGZpeBftiGxYzJfgf
naYxUHb2RTqxyMZIKyN9f9POIGJxduW7SLHAsAIHp4MuUZEZKR18at0e6n8ZgY+W
fK3fNZJk0ftg7HeOIVz7Nb9gP1CZf9oI6MB7NJ9TWRIT9Zwb+TrTR3wZBLTkG9df
OtQyiilI+YUt+K4OR4hcZHuhcvvH4n2vIIrgq/1mVllpyvVunUKGKdEUaiMN+XOY
87JbIK+whLF7eM2zzyRwsri9+L1AjU0xKjMjC89214O2nP3PfTLr4JSuVKl9Oplt
i7dDuPSXEUhF+6E+RrfRMIgTA6y+violAwm/VGIqcrecfIruh6hAZvfZfGznO2I8
Qh03BjvJQAGC0SRW2vZjtkkmKK/3IdxKN+K41TWBodKS6VpRWD4QZnMXy/B11zuz
6cxLIEpRPcdo+sSfPBx/LL6oiyq6cLyDo8v3iLWBJaGPlHaV7bZgSmgspimLSVf8
rCkMjuIp8QF4pQq3qsJTsPh6eEq8YQnng5Wpjuy7SHcnznvzOe4WXsXE0yVyubAH
aiuQCqin5xaWKaCB6BvPeOT5a+NeKuf5M8PgtnA8wzHH1tRPCpb+YNh2IPcCsMzA
CroBcy6ELAFyqu9E07H2DbHwXZpk7yd+j8iUKpEWq7/6VmbxOKi/jWmcjGUtpQwW
RZqYA6fjBgFjloMepIu0dOicyHNbgJdTtzuROBt9u4kgF8KAoveTRJc/1NpPTQwB
EgZ8zYt7Vgtio46BXswbhzsm8BeTAZJR1QRhnge4Uhrr8gzoMbQ7XlHT9jbbRyDZ
mZNqnbiIuFc/kA+n/+K7cIyikAwG+bLIjgJoGwivtA3FhC4FCHYS2j237rud3GNG
+17z7Z0K+OVNHe1mtcPlsGGT08Ng5BygPUsxnjunDdgSOcVrKjJrI29nvFS33Nvz
SmH0iH/bxGTIsDjYycU4imOQmzDQfWPlwPj5BlXNL5X47oAtBoCCUg93IO2n06bB
ZFuAqIb7URZqO+edHEb/7wUxCOoR/DP+Uo0w0MI64lTA2W6Co1SFT2sJaVlyO5Hb
qlTJEkHevzs9WpxXVD/HJliQFaiOFxlmfk7CB/kVr0NFs/lS40QlcTqHr4CfaBtL
TM6W3zcUVmppeGonY1G43G1SKyEEm37xGhGRDerS6BkpCLtinKU5NNqfrJlaZ9Xn
hLzpd2lCgTl/6VtT9tutNna4x40Rz32QjKXGtKRETs8PtbkN9czlEtn9OdNigyOn
on75o99NJ6y0/aAs6V2YCCdT2IfeFgGBhpqduj7lg88wAIEeaBCu6RmXjH4S2RBO
9QDBxYX5qxl+tkAQHixTrkebnZiu7abckHa8svSpgUU92dZT3gQBC8q7KjlMmCJa
hlqnSFwrC37moeVAyDd6yD/CxhjjeK19bz5iwOGlcy85spopexnluSzNr0bC8m55
/kW6mtWKN19ph1SlYf0UM3k85wyiejHSLxC/1UiQ3WmAzlEkcm0VB+bER2nEWqWR
uQdtNDlJdb+3/+tPV3As98Zd0S66MWUKYVeKXxfl/yOc1r/m3vWwdMyREvpbzOph
iDikY5lDXfZbFi4ZxdqSKoVPcwHgajh7h8cUjezHGzAJ19jiq8140Unbzq7sp61M
CVxlV15buI5dUyva/EFLzWuMuk5p78W+l2lGiu77T91S38ia+XrTvLEYN32spM4e
lHWEumMhjkgumnzEG39+kn/6+3ClzY/JIjaPH1tHKS1PXJYjFEP/5A/EERxJCtG6
9smfpEUuYtdU0tEYV2fFDlhyJEH5E68thNXN3U3do5iHghWXVQV7MHtLz2Hk8uSE
FdUQC4ksMVFVQ4LK8ZkF6nogrj9+dWsikPvDi5eR7SshzofLNrcG/SF+p1ZYNH4N
Soxapmcfeai78njejUpkcvw5OptI+QrrR/H1s/Vtl4ftp8pRPefBEUONTmtPpMET
Fttr4pkO/kunazStxpYtD2SYeWn7zXB+xoGaSSGugKIKfvNcwYaw6oNOvxnnr8Pk
2mTshFT6DKdVzja2JvQEZ7tbCdjSlYmfFs57FwjbMUK1vamOzBB1R7rIJGLvlghj
khg7tHYkBe4wvAGJAjXZ16T1c2KesFYiW12qIoygUtXtiMQKZspgXV6UIDf4Bb72
ou+OxVhcykijMmhXsIBKGGSRtDVOvywPlUMWwNxizQfq9Kfs+ZaMeQ1WMNK7SqzO
eQ6Ousf7oLfu2T9kD4actdZg0pDTLE2N+2cz40BjNdXYQv/J23+kxGD+h5BFn3P7
sL9749Lfhk5m/A25ZFATviLFj3khhi4dOnbWoC+y5Wq5cMyDvi333pisjZS/osHS
H49omopiT8/sdDt9TaVNjmYhCQ+UzGAzn07vpLKv5DF8/gMwXBdW24+nTZ/dv4JY
jXtlG5m6+SB11j2cZDAAbnITv7NaSbbyKw1u0C8nSmvXwy2TN2RiqS8eVysChP7K
+uH99Ho+UJqN998B6SFKJawX+MZelqRoGgwJrkSra5G+SQy7/sFwx2QMUUnMYq8P
U/seCgXO1I0HZjs6EaBafPcz1v6/quy3GzQHsjupLIngNA6GXCD8MosS5yX93Vpc
JFOzYUixIO5I1dhDNTdavOKktWkhegskSkpl5Quq/XRve4JXQU1OK1+tB7GUeGrX
8dmkYzLiZ+N+vEzffv0+a/rNCFcj4CqNM/T6mzkfl3Vmgw3c583Jig05EFjlLP+h
6+vDBJiT7tHEvG4QiH2aeDsBfEqMsKrlrxzqeZVrBmCoC09NY9RrBFkgGFKWPwgD
tSaHfKQZg0PzMFtWTV8yMtdxU3lCiEFewQRoGFaWPxZBNSY5sgLOCT0Dvf1yOB9j
PKbePyzS8SYAVGXXS6AgQBSQxmoZCbUXLfmegkq3YSo2a3iMVwOUnNXJEZb5REHD
kwweTauabE3KnDy4B9ATmV8dFN6f0PwlQ2BJnswUlhMZ3gnhk+MpLqlANrivSJtM
U15ii4j0cSYwwhxXEdzk9BFj/jvXgyXGSouWzKAZ1nA5+mhh9r9YCaHwv+JfgcVp
t/kP89ee77aPUl66C7ErXkIe2GUoF99xOXXJS1hMlE1u43/1xfq2Vonc+C4A7Nfm
fCOpMlihPIz0rLKH1s1ysToivGqAHyAfZXYMBAP2AKkRh1FEYjcXhqryuqhcWtmV
/aq7EyLoiMjq+jz363I/BPcmbM+Eenq9os0c780aqmNuAVTIwvLsNe8ZcglFuIuo
w+3NkceqS9/9k2kZ9xkA6Upbv261iyD7M+gWIL8gRwpWUZ7XNcLnlLX6LYHHoTbq
Q29eVwhYm15mHHlf/VmApcnAIjb/ioJwXjdxviozSLwNkJueA5wzo/d5K4vvT74F
5K21Hp1tlMQp5V4jc9n6y/80AVib7LPGK3OsjunIIXSYJJrHy82v8U7mscr3bbkF
6FdUgfX/IRf8Lt68s75JGyNObnlx64eHZjvl/0sN8xPhEJa63XyLjF6/HFCWvvXG
Ma9IKlVCwV66wRRmNJE7sD3u5cTizeCq/MGbro8Ea2odHaeCd/zBn7ztk40NUREd
fJ2biDHY4XdJy8EuhotyBNTfi3Rln0STd36YLU5WGX4lTRbIRP3N/66k+Tf0x69i
Bdi4ppZF5VZElmnJM6oOTPcvHIkCH/iQVUMHcz0EjBrYDi0BnAz0hLJnyZc+6/hd
tmQfcgAiqqNUHhfx43EFrky/fRhNGV+ea/5j6mqZ3RQCDE9aUL8l7doxS9wFxE4G
nYmR19oRnv+oCDZUqzLzYpeXQAw8OW+6V72f8p+wOwFpKfrV05Wqr8RKgjTLu8w9
`protect end_protected