`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
gfpsjEbW6UfSchdl9yxrheIGuOiOB4kllpRw2Cv7FpwyRpGZ5e3tE8rnbbfhWRLK
CBLNdQM3LmJb35raq8zCkwJtDyIRysHQPlnyDHVzVIgRQYbS2VnNNVKCqIMoZi8n
BwMgNh0c72a14fyKGi75nzmAOr8o40Y02X+35yjyPPybIHOog6Yq8GxNU7WfSuSl
aFv/D8+EsGHpDP0Bdbo6tyzmAfejZXTKReFkvce1DpHNFiVMCdryIK+TuOzc6wNo
8N9Bb4ay/VnLWxtqAOprXDqkvCDkKPIimKR+/UcslzWKSgve6JF9T1pDxBGyrGNH
qoV0J93sKKUwjauViSXmRAW63jO/dDCTH0512MxstefR12iWszvQmrwvTJRlCpYn
SYcaxGkQrSYjN9QrKPCdj3KHZVRRHI1orTGGjfnUX6yRYxas6i9vInCq8HENW/x7
6N2L9KItY2BwU57RM3Be0QqHFurq4LhKYtsXtvcYk7xKnaUhZVFjlcqPxbAqThcf
KGas0lznRJfGZzjou4bmJb6pKqyyuysfJwinHS6ErbdR9WuiOXbzatr9+UqHxuEw
S4+moqMhxm6U0LjJwc0tzUnoISkO2X/YsaqCIPqRprZUQyd7lVTBSPeDBAiuY38l
YzSd3SrPml9FamApXmuABEmCqL62Iq7NE4l+22NFv3Nw2Zokv15BUtsx8ExdyKr/
3K/7VjDnlQvvce/hYr1bnT39lHbmtnRWP9dmRxLnA+YwRIqxeLof0jegjb/L2jvR
7NRcCTAh49opOP1UxnOoxwRSpqe+tDqXuyBc//faIa/WoWRIHpjq4almyFeXTOlC
prEROVnKdWEW8nVcaFmiJEvTihReOAAziw1aes6aXEP/yGOF8xlGPJHuTshl7c50
1KFHbaH6WMyeY3Zdysv3d6wDsoUCNwByn59ueVFyW9UP12NPU2vFXxfHUHbJZF7f
S4dnOaHkjgBLK/wXFU8Up8/wMoFG7eK/bZ9QdNMFv4wjCF/kthz3Gg6QD6onuTbs
ersVB9xivAYFBb2khLY3nwOJkP6q7RYE2mKp9mt98nmqjgxuJcVmAPcm9ahopSHv
k1VDQkBma2moZRWArEbBVQh7Sep8ed9SpnFNOBGQvXlnb+Og/2sU1hqh9hvdnBac
iLUTsym9aZt4VeEMaKsCtZ8pH13oXxLhcGzsL5LKq3XcldUZl9YGAz/rONUfB1Mz
iRmdO259qL5yjxj03aRYGrU/4pvoDtxCXHjsiIktwC9f3WYg3qdGV5eGMZjm9Pac
MIZ73mnQ8/ZxygC32Epz03E8BL6hRo/JAvpcez88GPiXouAOPH8KWNsx0swVMPWc
rY0CZkdq9bm1G5UVZMvgPdfL6KFWuOUcUvM7O74KPP0L7JySchgS+QMQdBS6dcLx
9srjEFsuOxoAUWzExQHQyPvqH+ZwABXSa4ZEpuTjUOEA1cPfjaVVc9Eq1QHeJyAi
wQ5q+jkI8jl454u6paRlBUsHlZQEwiSy186jxpd1wbVa0gX8Z+udsUwGJh87qqyo
EPNus5MXzzTZ4XtvGzgjbSd2/MNEaQgrbJBp0a67knXUfnhwmwdLVwXPAFkOhm4F
jL7QjPra1kLIlhjyixfYzqrl+3I7cqGzzgU+IKNfV9SrgYonlbJPmBv/v0q3gsIh
7s49v9utDa2/oB899zfVzBfBHD7THstN0jUheTA/3jC8c2+2P938MIRm+Q4By0d0
W76UCeRi22sb7PzpNylw4rbfG8nLL6AdKcAWkNdq3p2l1g319kHqej3aQMwmxUdx
maYMG1tkPQG4quo/UqYACP5yLUkoDyIPhKda7/9NNiNIQifOzy1NpLv5R06OTNkC
0RyAhmD4rQ31dyQL+PKh8tIgNp3svS5Xf105QfoOE8GHe3VdUrZPOVBG+XubMp5M
J5AbPP8UbQjdvm+PBY+I6mEbl7ZsP0Wq5wpZ8H4ZrqPKwQntlFvPcri9Zisyq56f
cS35vUoxVxB8jmBBH6HCPtm2KXHHeFRPBaiJnJpkTapbkfE04fHwtxJgc0x4W0f+
aQ0zdFgp1IiH+4aL49Sm8AmQNWZYgXjTU9OHhJse03wCKB+YuOEQz+RbdufqTueZ
UDybqASWVQ3GiVuxOlF1clUBE9ZRmqBVzbj7PY7trmMkHYpiVRVTyzVN6v06P3KI
cXW+kdyOozZyUvscVN9J9SsLsosZRUzPx+4ZCVWgM6Bv0ed13X2Kx500E2fVBbN7
8CJrnNEW+zJ1W4djHZUh23AK5sEfwdLQP9ELDQj03LT+nyZVpPXmdNcwkAueQLYR
jWmPtd+kAqHJds/WC056lteLdgDdGo/O7+ZD9aSdm2ydcQ0iMNcyepZ/QrtjNEEV
O6jlMR2wJn/RfDWGVeGNSlVpalr22FfVZx5TBFkBAOAsIutJ5EXR9bylO0PxX0SG
sqKKBuMkQJF95Ub6UgtbCJKjuFUD1ZCT4hP8T+mPkON8+cxIRaAwKkPFIaLkZ32V
ld04pV09sReGt/iZhUDe1opQIvuwSfUVnqpA2vwhza966LCLwsgVuPta4EKXZdab
84c889Eue8EGjNTCOQxChfpUbeCKLsMBcds9clwMBFcMvNNmIh6xWt2W+FlUlsSe
gIOz6o9AbYYol25ngu7IE1vUvqIndO8w4ZVHKrC8XZbj4Q6AYEZ80fIgz65nuQ6z
89vP/spJhV6eCvz9d0lW94crx6ZdW9yN0W2FAWNmhPin5+v04wTwGmpQpTIIp583
lk9Lyhm0keojdyj+rpTZ8a1VpJTArFuY1j6xrAX4puoyrjzYzvwj3/7eY2s51tei
Z6WDQRpNpbaafATpzlCAYvPq0x5l6G2qLYd74w0m7VSDRiWN/aQuDtGPidBtC95V
2NCjyNAQSlaE2sXxo5f88LmuQwi8OuEkKe67414NMoFifl6cWfKoWaCD9ekypUi2
9L5MzTc1Vmux6CGj7vAvDp3FacEatxouDkdas5cDgz0AjchSYB5+IiTIgd7Ylkj1
M33e11IXh8qGfogdTJZCHyH8rnlf5ixyMcsThX3ioiqoP+ZbCVx2yP8toC0LoQN9
h6COqG3517fRVpEWJZpCqBaGD4yub3g6kLd8mG9xC3vte6voBfghO9Z9ED6cwPtk
gWN+MY4e32bS058oqCsmxYpTY7teu1L6TMH64lQ1lWTi8eCuxe9TeDDzS5J44egn
7DVAzrmkQdOC47vh27LZ6K63Fc/Up3MZDLON1lCDjXcP4eUN1uVR4EkBvAd0Pdyl
WDBN91FaPHuuZo10EmE4Ge8rJ+2l2SpF0aAVso6pvHXL0bhjivySD7inZZDfh/h3
D9knGkgk6+3M1HGvNwedBoxNaPT3w7NkrGbJaVKoT2DtLdi1ucM3CspaZxlgUkK6
S5dsG3WiVJKKeK/pWPXmMnCKZt9t1AooXsoUd2yspts2ZgfKfa73132wQz/3/Njz
`protect end_protected