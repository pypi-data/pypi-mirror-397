`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzT5omKdoi9lai+a0H+VrzCT3nhHPu8olGfM1d1MXlYbe
4Q6hi+Y8RwX4Th8rS3pg+L/OuGB/u2M/NC0CYWqnZ+eoE278s+mZFBXDZXYUThph
91p9YPUHlsCYmGJlpjoEdf/0mKh8V1XuMkKnLFZ5/X5yxmG/36v6GP5hfvfDu+Sq
TQ6rJJWyFFI2VDngkxCcuM0NHg6hjvrKEpEJ+6O4iSqJY/17T8rp+6C3nQLMvEIQ
JC3mKwSgRDOVQO81aKbEX0ILtruUcASF7IDHi6vmHF2jw3/zxY+cmNigt1r8mZzg
pXwRMcVIH/2lYJp9SyuEAxP2ZlOR1qmdDfwr9rpF0QzQC67jFZWKPq+lD4xWB93I
PvPyQF2IstLUyLfalc+MJGqAfci/TTu+FpUSX48ApTrOC0aKDTovrkeasSfP30yG
JlMxCHn2NubcslVfmUNbo3h6BXfoFNX09xsTzWaF7Vc/CtW58d/ewYrQQ/qGb8J5
4rdFasoaT2A6fh2H0oKMAA3CbTZKpNZsEwPpDCXOKB/HZi4ePcOjBWwuC4Jhq1aB
XKjKQwIIXf55Q8EXO6CXDRr0Vy8CMVDRLhQCjleW3TIlQw4tCOEYu9u5Lph+1/MW
geUm34aqmg9dey1JIkzZ4HDcOweGKSXxjHX1+czvlivOW3zOwAz3c/uV1KQ+0mtS
c7Rr3cuXI+Ma5IMe5NVzmQTTyjpD+pWzZzjNoLJUCpVJtRgbDW2UMwAoSgPCACnr
v9iQQvoxIsRlHGcahfpxegpmGez3GS04mGqSatT8tJTziBySG1hPeGedYCajqKdC
t+GjGLdOJqrrA2KAqToRyRFTesqeuyxQvZ8wUULiiwpcDqafuQPpDkkC5ApKz+Yv
c3fsQZ9Z6qKrpKXx5FgNMmALchDfqp5VevQkAHrDa4KvEb95XA8WiE1cQS90NrXb
Y4ONBtGcJR3GuaA4X5+mJKXa2Gz4nOPBOGJJdFdi7zpiu6MzrBZIM1V2Alf0MQ4f
biR5kg8VvHLuHa3p0eINqWxLCsij+52AnCzV4s2MyBKYA4B0qnRgruKXDg/RO+pl
X9Se20oX8IdHv/yvLr7uM5wSuDEhl+uphh1VDI6ThumxNGiq4PdQ9izvjiSOhwmS
bV8DYTEGgtVUBHDfqhtVOalhtDbqmjcrT4ZN9HsI+j2ujKlzbgy3aEqecOBirMv6
vTfE4ZcXov6aEcAvtZUeSy6eeXB+ZGVlebXLHbVD9kf8Dib+lH5UVCIIXGA3AGu/
1mWtMOwHORX4UQUqCwmpAuFDyF0xd/cxno4ORIFmeytVaVRQndFNQ2cFve1CeH/G
tQG+Q9hrtlsnNlSdF8A2pTP7xf6biVZU4y63Nwa47Bx8dGevcdUTX01hjnOmv4k7
Zr5Y09ho/RmmWWJCvozDEve83HubQJhyPVslj1k4wxkL/EoHbynS39QNHbk8v93s
ls1f0tZp/m9pvK3MmCQTgi8sdK3+inpqvwueX45EmfY9XL7dd51WZOYFGw80VsMY
uDh/EAZev3wYrd226TvsKVtDI0cdGk3C63hV0Ef6C2/NpMJqeYAaZaxzbazyUUE4
CunbBRZ25VQ41LkWRpOzPnL3p4j62eI6b+TcNG9zwpK1t/t6n8nYOPJo1NI6HR0L
wBMoJFCnk9whueGiExTtG/2j8wOlC2vkHTpI0uZbMpAOLbx0prIWb9fiY+esVyL0
rJE8OLNm/evcr2ruu6b2Q2yPIqMpLV/4KTsgGrPBULMKIN7jidOUs3AjT8m1kFZb
Z4WNVZ/ildNf/mOhDsRcdA8FsS848DGLgaJmMARjw1UI+IvO9Rgvf+Wi5R3sy8fn
LaJJS0emVBFWu9ch2RVtjpX7KNrCEtfri7jrlIi9JDVLStCNH7snlWbzNk/8ij45
ANFgG2T6monD2k6TVu0a+7oAb8BTdJhhvK5hD0LmPE8UTGB33xoxuXSEHlQQ0U2u
4QBgnS+g7atnvn1SEIQrbzZOGPfw9TDVIuJijQ8YmRzH4teP2zMX6DVXBGoNZoBZ
pLUCxpBia+SE9GGnSRIbDcPsJ7OWgZUb24bDciWpYPYevEHE4e7XNh954NLTO2b6
s3X/wIbMLMa8HmsWVwosq2GHbgFJdZ75MwIyJ2396ra8hLMxLQxb7xh3U4j2r8M/
OUEkdtj7U0XbDYLf7fr0TYGFLWvRT0YFJNBFeVudVpK5/IbQOng9GvNy7hnKNsMw
jiKKH7tZasbcRSemGesAWmXNIqZBzz9g0ujSlbjKjEdTDPeRac6u5hDACYxZzjp2
/6bnLMCMJjG1AVJnhd+4cqgBVGTdYcSE3BM0vL/kIqH5a4SO5WcKmHNZ5aRqijUD
lHy4SFGHvrbzrCQBPOnXHpuAqJo5HcQeO0GFlHb0hVmFLbfq7dtpjmMwjziBgnzl
578XRuM6VcFCNphMecamrf+2jrDcf4MUCVOtOlDcQ7XFH1OGP9Q/KI8UT0VEJtIq
Z9MfIEM6ZeK2HivlhOQj0sHujCPGaVyZauJ846Mc4NxIXwgqE/38HlD/FU018BqQ
B6SfidOpFHoc/dgdEXw6Q3Atz1uTekGOuAix0SueiFxhxW/JEtZtnNa+rKMKZLsu
jGl7ct+A+ZdMobo1wAtJGLbMYQUPviEJuI0QpYqzwRvuu2OSsrR5EAYr7CEF8LsS
p8pOR7Hjd7S5xgHhLdXZVr4cUTj30vfLcoc0xiTezzzxTHAZuZZAbE6Ht+U8ukLZ
CtXscnlQ8jrHD0TX3hhM5t5luk7/U+DoNROTpXCTNHBbdJWEBBhf/zROy69bYUKG
Od1XZGrvf5CILTCF5PAwcJKR6fjsIgPHaKKgXOa2sHPSF8Xa2NM45Rj8AiWXDm9D
JgoAso3xmhpep9Cbkt/Mf1HSOvZP9z53TKvVZBW9XK0fNfBGPrSS4eVAG92b45f/
XOCJ2Ffjq76rYbZP1oKYgtMMFsF8roX9i/+OwnIEe7+lHaoKs+dcNLWHGhROiyWV
trOvONib0iivx5+50JoRjXrW1Viu2siKjSM2BweLTvgYGfPzF34Uhu/QEzuEXgqw
yOC701Xcl8fUBeO855ra3m3iJ/8wdVUQI6r8mCECkqT1P8OfZd5BiJpPmw+zQvv9
0hA8XvwlBgPmarip4n7r/p4ZAYRFq++YWBjXqNB3a/+L87zSW7lH2mpwYFZUTHWC
/n9daSBmeZ2s3TvJQxBtyjGGQGvO+KP9OtBLk8NVrMkXeuGJ+auJ4kBsHcL0DaL2
i7JsZXCcyEtZNfwrIMsJ4H306VtsyaeG0HEchLirOm0h4pnhB5rOiCD/NOdKZoR1
5TthfeQNclOaKcJZdiU1oKDklbO2HORfmLDu0NFNauN/QY2FeUewdCZJCgmOKYlZ
VNr/cpiHtsum3LWcYJ73t97TALyoNb4cU0XGQXmgLKoKl/tmAgpkslBc2z3rpp1y
duVdOeySB8pSQ8iS4LkwrPy2Ct3RxNRR/LWplLkAHWWK7101qkQTE+Z9E2IRHLc0
N8ITLSQkot/WqiM9hhhS+28mnSJcvdC08FXGVCKMX/tQiro8RK62NtgrRYMC2p+n
TQ7jVzjqxmmoxUN9nbZcbYzhanZemoMNrtXVD1nHPftZu1uKYns5IJxJ/pYgy0nt
/rihY2WiIXzVAoYgU6JdNGBL9LiWuMkV3v36/zi7CakwvCGGOjXkCHf26FyJX+y6
TY4VqWQUnLK4dzjFakawpflacD9M4HEihsW9hz3z6Y+v91Qfzkn33/6jBqfe0UYm
OQMrJ0Mf7peHWbCT65N32EpwcKnZifZ+Xmk5B04Fyqo+j1v4ltqrhARWTuYJMYQI
YHEI6BeMJrePQY09Sylgy8zxNwVp0Rfu2wn3Z40CtHRuGZefFbEYUJ6sy0VrKu++
KR60tRPkK9oVNYvxlGLzeX2VQQcOgNvuhA302qaMpHrzggayiE8+sRst02XLRdc3
8Qm22jg6gefbWDAqZi7amyc/3++VbktVZzqIiiM+W3rC2Yw4qJ8vtHqEkVEIQ+fM
TrSdEss093YIn9XyfbLMIidseDuFpIrknVAoYZyv1iI6HSAQHNJOD30q8Xx7yGe3
2zQe0wjNtjTacmPix/RknuYliQEh40ru8SMt7EMt0wxKtrZfmonYmM35QISB5Jv7
zBC2xSBGf51M10PXQ2/w65YO4qkHGbUsOo/1L1dsaOyflZS6CiuduOgucEKtHorg
z1Y8evj6vPkCY3v37XxuxfJpuN7wL98YkvtUp/BJ3BcatjBh+o7WSab+uKpajG2K
ILgrpA/N+RLRLZZqK5hMLzrR0y1RgJ8ae0yvxqFoLFhYCb3f+luNzoADSU8hyU4C
Jb3R3ll5uqy1IKm79ZeIDKTd/DhN6ZbBVmA/W5/mX0UkcuOhi4wlJPsl79TRghXQ
e9oSuGd+cy7dH9XpfDYHYdlF0vsCK8zbV+NwNoCFHnhDfUUMVy+GfRV/eVWnMHN2
eKrZSqtuHcyYjKlblBtUdoYvnS8RE69eQf7nZ4R76LKlIGynszNrovhU/rKy+Iz1
+n4ijXcoj/QmdJz1dfDxGKZqPXgrzWDy7PUX5b7Rvw53PnbHm/oygZFTrS0SVFKW
PtE5XZ3vgtFLzrJDJ2urQR5p52Rr4sVjrax8iwHYwPF4u0Nbo7OR287DTjZJjQMx
kqjZrl6k8kmDA7VW0usrlcK/2vgVbL2YPljoM3hj6GsJRGUdsVJHk0DYDpSpp9ds
3pqqvwd1jr098A8uMEeiCmKtOExbtZ7FQmxSHLmcTHpehZtDYxRGTJzutHW46EKZ
W70t4lazqgB9IFAwNY2gYzZ/ExNUJmGKOo1zvGn2AQ+aCCV4uLrGezsSHns0wYBu
BNi1HlCCxJo75k82cdU2cmmLGuTLzQdDPEahO1CTeVGNbBvM5e46T3+waZFgbwpx
5S9K+DCJSqMEyzgA8rAwdHeqIqNooVxhW1PK6zMA5RYFgX/BFy21UsWMXEd599+S
4FSsnHIh2e/d6B0eDqlgJpJh1E7CVXIuAspE9+RPhBPI5pq5AMMy2+Uv8q7/D5I2
KWYUyXennpPmR0uf4q6vk5kWEkKrEfLFpS9XZ6fpoDsZcmeOqcUwoaONx3h5H94u
6FiCkBB+jcM3B2SMvmeNRpTO15jd+fI/ctMluNxTSsUYpuHaRVLNQC9K2L18o6l3
igXmcHDrAuyoUKn3bbNRNG6LP5Gl0mjkNQsvue5ERj3wtiy4BoP90r9BMAssW2sG
rbImZAiw02KID9KMcwc9IMn/+ZMm+690ZryUr0zgQC1FE1+u7Hg7M6DZ/yPwiXkh
JwJWocpATlcgP/uWMK5obCl3Xw/BKZk3MZ51o0c2jb6ditxU40IqqQRy+raOXL8E
5iytXHjok0ZfUxzuhO7JQz8T30JyR35msavnx+7ZtTlbd+luz0cBYlYA7bTgCG7Z
hVnm7eKzqsMkpUZuaCPo2f0DCw+B3mpmcsG/r8g71XfvlbsrZP1sC8q/RqJ9vKAs
i4+gP3qqZxvqcD+YAyFA2u3FrL8Zho7kJTlJD6N60cslK4MPp9rBsiZugHnd6pWy
kqBZBy2tTkNT7hUWlk48MIuq7tThFDaotU1StmfA/GoQHawTdatnrqMpiKWLtUCM
acT3osIEn9V4UHJB8vRIs7e0CKnIwI4uttcnkTZIaH3iszT9TpQj7qV9Z1WpUhpi
L90W2iOpBDQn7VkTCrUdRW4cLI44nUeqF2b0h5iU0nbW0PXnp8GJufKMvXLvFXi1
nlQqbfd5GikheTmkoTDRC6nQ2lAmHR1mv0cgsb4lr3O3ePgd4C9wbLXx/fYfBosh
gLfatxF3VvenVAExBpt8b8cah6keLqTkGxmPWphIYuLn5AXCh6Kj8pPBOUX3Z4Se
ty1YxrAjIXJgmWOXBxiMBY133wrqhCgBr4miLw4gh4FP1Cls92HImc+tFRkH18Af
JGn0dbOmwykgsQdYilXf8OXv7SEb4sX/rswA52gRKwBwBp8LmKSQmMeTlDiEwfLK
2kR/P7oJ+U+aVG7UMtXKIzBhxjPOR1acqozKZeYJbRNyYZp6PuDk2CG0L2tPqIZW
dZUF/QCytFnyqzwOuoCccFh1v9qe9txCLy+Vudb1uTWs59jg8GGnCfREewwHvZo8
NxzbR3XDbhhqFqqIrnuMT1tjxmCNoifKPxbaYXCzUccrmPH6vIHxM/lAqpyTM2jp
F84uikZxjFIUp/yI2i1ee93D+/YqU7yzH8DIMk2k6mPsaBXs3qYFQEvNPBMPvKT4
+w/YATWm5UXAjqgabv2S1ARGkp/BOK+iU/7/OWdOyzlkCJQSgaK8Oh4IXe8BS9JH
qWnHhU94CNzKmIIa64T2foTbZ+FzfBQctQCCFA/h8h/AFp/Casqra7ZSBbE5fqSC
bBBWV4Ptlv0jcT/qaDf6Rn3ZXreSGx51bpOz7vjFbwgyh+AOYK7JAsqAyDp2gvg6
nV6aVoYU5lzfLRT9sYp/8I2P1MWhiSJH6dKTPongBQ3CbJKZxUS7Eg7AVU0fEfqg
bDRQdmRCE2wldPvGIsKZUf8DX17iYPVitUUiObi+H87+8rJ/SoUSoyMU0ZeE9uM3
bcYBEkQSGPEZingF6wCgBieWa794C/vCjnzCBQmTrShYW0ar6LAAPwFyRl1Z2yFg
XiRNIWhBB++QXnR/yB1rS2/p6PVb438O5Zf8f5ZdlGnNqiOCpL/ufj4k6DYyWFnY
Z+GqjeSYqZolBX0lRUF9n2LhPbvHo+5oqybbxNahruh0qLxEzBgOw+5MF1VOMyTr
FxkWl2OGaBDne4JgOu88qucDKdTrtHRCwbDg5mpVXqg0mVptyPBrjhPiAJqhHQLw
yJsFnYsiD/3xNVk0LIcHzSWYkbfotq0ZPhlhlqQeY4Cokysc0U+T5zqELJBHwR+M
PT6YTzzjLRu7s4BnGTptDRjN4y32OZwBSMg6ytl1LriUgmyZrTpcbjMvuJV+fAt4
NN1RfIC1EPWRVtLi2Igwz7bl549ttvFcSuZvFqgCwDrQMDE8LEEelf8OnhRG8J/9
hANpKElVuAGmhgfkmBEqGLyyYGvsH/HZtqRhozi+x++d3bZPZ4AYVZYZM40+DkxZ
WzXrkIzN7a/Fxj6C6rs8a7Vg6fnDcFUZEC8ZzF7hJ+bexhIHnrOyPu8NXj5sdKyV
kZD6KTn0x13SvNN2qz+ea75VCd1p0a55ZJ3ToU9x/6e2Mj6q1EY+qj9uoDZ5sDRr
+PX0hNnUqlfshQFqqQmGTnrmq8wm4QV/X9Dk3epjbcnwufOEJrMFor7O5NSrIpNj
DrgJ6EseB/qZ110O9NmVYgJsuwlL9zKo5S/ANEfL3W3+tEsPz/FAwGvzSt0Jnc9s
iR/fy8M3xYL/EaeyVVvnmWk1x2oM0LRIFxhgd9yZY1F3lbRBxQJzrzRjSwbK/7Xv
sGVmpW22uNw/noheqwFS2BsGEQf3QN0nRm10XQ5owIQjEnzu82T8NrEwvhOVZ4Ng
Bsvug1FIZZ9cBvpmzzTeDDJI954w8Ik0s3IuBLzHAva6BuYfhCI9tzsqjXt4DuiW
xa/l2lqiag+Iqa5DVnUAg2j9xsZSBzGzWud2hDp7cqSicmpTzVWkrz3kYugQVzi+
0pCdAqk4pyQtZKAYH/wE5b/UlMTNgWzZAVuAtHdss6vq3DRBPQSlpBWo1Qm64ODb
tCPqFMMdCZggz1iv0L5wGNyX/O3JZhJlIq1zdlLsOkG3++TYQiyXYxSrU5cImGyO
VV6ue2WPLDNT7gbuF/gv0KHOPrJKEsfjd2HCvmnD3EOTlJZKU9JuIRszwutxVgfH
utCqvXshBba6mW2bPCXPHwYpGFEg0zA/CCFH+sbGZKSxyNGCZbNvqGk34FACMTLF
3PVdGOetPwIE/ABppVbsuDe9arDtjN+qj6kJTFZ8e3rsg0te7aa8iazSkf61SzI3
M7KhSKHRW/ugqcn+HGTQrJRrR8N4WRGVfYhdpfaCvh5koVG53zOkLgsliPiW6oXC
530RsXfd5ZZ4zKhg3Pa2JHMb2utV17YSRVX2Rn2TsGRGzndJ2yJJNZXqNDrl+36t
JKgucdTrLmePD5sVdCaDlWkog8N9rJLRTZHLJqCJZXYmke5oyaWwfxBSQ+DchBZO
PhynBTLHHawSeR/RZNzyWNkS6npmDJFI8KogFIxd/ol2XwlQoRG5xW0S65n9KkOo
IgNok7xjXS2VWkXEuTV+SfFpmL0JBpsjVvTSvYGbLjOo00ZuAUfGKvY3m74LJYEx
k22XW5lPNXELKDr5pBb2FeUd160yshHUYGMhcIz3GXZB8gtKmZ/cuV1d7yTxaoLX
dRG1A0/Qo6Qq2Dbg6K/T6ZrOKoZFdYgjB6XniwndVpAkYWVteHJ4K0S13QTq79zv
intDWCvc4IEw2IeOvG1vd13EZwIcFAZz4LXfHipbdMgfeiL+7aLpIqm+QCPfTAxH
L01hqLDY0aJIEMVCCoozUKaIe16ZfEuFr146PUSs0Mohb+yHQIBFE7SUKCgG137T
0fdPJ/Ot7qDdtXrOQsFYflYRYPKj9S3Xqh7qABvFB0eyhlF8x0V7HdFCsOjEy1f4
8s872IVxn9aOjl9ZoKl+bPbj/zx4/X5DpJyJk2eJGSQoE/pDqKx5JF2W+Uwy63SD
6p/lLaQ3v21RQkLZ3/FVT3/xBuL5/r6jJBpMwI1z2YNWqUdnlohF6iHeTqR2+7SA
8iy6asF2Vv++xloYij3dTFUA/vJNVJ+poC4QF0kNrO1kGZK6nd4SKy4gKcY2D7Vg
p9I4OPaDOqZQSHIgRzxUAEtOTIwV3FfgJWv/Jz2PEgWlFF55vJtzrckCFRISkn9x
ucDPskXo4tfSe7K0loLDab3OctCTd41jQudf0fqs/c2mJy25HjexFDQTv38KLKFT
iGwKnsrOURLKhlLddC0b30uNFqbWHQaqaVytrcwxpGZQlIk3AIZ4onajVPsWPw5V
R9yQzi9aDpzBAEnearX41fCeukHgur7Hdk832tUXncIclrrxU6c9oSrhCWRWmRSd
xVq+QaG9IykXVUAGhT9HJQQ0wj9n/cJJLmE7oskc8BJ89E6e5+xf9PohBLH87Koo
IlUbjHxxvvEniwcxy1+DwNACaR9SBQkbk+MVDop4NLevItkdWwTDSAmPe7xqbjXn
xRguTzrADCgM2PSqKRs1gh5wajHxGPLKaqh0w6IPI8TMFYMGLsyfDUGUkm+nATRv
O5rIV8BDXIUCQkxQiIJDtfsI7B3gYyMMmLwLsD7hItSRXrOnucV7/BK1Hs/jCBMu
YuQfpzCCAgq3PZuOoh5N1xWtIlPHb/wqjZ5VXlARr0Vh3w6Jsvx2S/d8DZAqbFAc
qF1AFVPRi5jc4Dxr1Roa7FQFumwyxWXA8bxGERAmgd9jJaA+q37xnfCD/pH9kL5O
TYEuEkDFgXK0OOmFJmj+qyaPfH+UqMe0JRcdCDLKXPoOuQ29NKGYvALHHnfsBWvL
uI2XcE2Yjh0Y1jO0hYaQl6P/w8FB0I4ojvGADzVqOYincXSzRt9UvjRCrWsIcf4l
bFbM/6zMG+ek1sN9Ac0OHy6zx2DL8lUHTW8s5DWny9BZyalT4tVup31JUk//BIlv
KZq37/Bzl9yso+i3yJLkolKwLlyBzcQKmqdJLcXkkGqn8rGQhElUEsOv+pQbWGjn
SpKyrHyk1Po3e4ru64LZWoAqkV1rVsNd4hGG6y3BTnlRaHu+noKsv/FT03uoh5+2
/SHbsMTIZeKQq6FOKJHaPy1kUPW1j04sS75IeRGkoxTXCci/IhlKwntYCFWGLrjI
bCyFWyvRVTDq/wIx3XExECJgZhrNsKziORQNzmnwUApy0bm5yHI+PubE66tB/MzY
7TTSIt7sfT25lmazRrS4y6kTNl0SN8kUHMxkQ30E4eqz7/zDgTNNnTzMXYq4By+W
jaBWprf+6cKI/T3YZIGkomyNysdRXOFB0zJ33DXPDeGnJ8Pd4axNobcITGzf2ux3
bFLTWNHtDMFLy7ZdRfpkQMQfvD9HJPTw0bGOticyUJp1raWv706J9Yb3SctbcMBz
yxlGs/5PLaeEM8/BxDFJBV4GLellmK6dswgcvvEujk8ynALxTpk8dYeCnvWth63q
Wy+KujbEZz88BsrG6NJqv82Npmpp/hSRN/fOL/44lYH4lsz1AKfIlJsSgUvB23PJ
oYq+IEeGVuqNhSE+ZWCrhBXTq6QBjGI/4gV6LF4zVYw845I6zYi3rgr6OTLv1HCJ
gO+XXN5fxaP8OS5MVvG+yscU5vIu4Rgey1Aimpq9o1ANoPgn8a06hTG9pBWDH8Di
3z8bDpp2acVOLYgcOuuW9djGQHUlNyjDayKOCCVHh3VwVeDRwbxsfXxSTMdfS+WP
9ytLJbZ4znOKbvHfBvPzUbwUWqlOK55cZ9Xf0bAQCOc1XLXDhL82iiDyTeas5Y2a
KuhM6gJT+oh+CIy6RR5iFoRuBQZpxLbvmMNEehNkCHo9wVUqXbk2rHfCI64lxG/d
fWZRwl7gy+qQR2Pk/Pq+rx8dSLSjZmg8lBjao87bS32tQjipAqQ0di9meTqHmpxk
j/KFiiqMhk5cYy6naqRsCnZSOVzMNP4hmNIP+1UAlCjr2FEkh5GpwIzPNK6F1oMl
OkOggBGJfoUJi6I72o5GognxFHW2sR0BIQ4cuVoROdXU0Zqcn5iG9FBoo6KStTac
94klH6A1qeW5SbSETGYslr23nWvZiJqofei+t1zzCtWIbIwMrKPtdbarYwG+415O
7BwrZlPxffblqwchvwWEktWsL0Ur/8t1IOBNm4WSQ8HZRvuz4FEN2xDAsmtCZfLG
kwTYykhJ2+rKqEgQDNdv/UOtktpv6yfd5LHTN9/E4quXmtt7pizs9cknqHd1gWMx
q5SXum5EW9L0HacL9SsXfiLFmw/UlCmSTihw9Pidh3H9hJLWpw+LEsuZqtg0w/e6
axWoWu/G9up1LH8P2eu/6URWwhAsT243vh7RXF4RPgIlJfTw5hMqCUa4akWTt3yf
FpLG6VxN57ARv0S5S43Z8oKNhMzBn8YkaLV73BnXVdDxDol3krR0kzRwPImYbZi9
7Iqb6VfQjilXNYuvZIj48ZLbSIxQOZozmu6FHxTi3U2DaAZ3vD2AN9Krx1yqfAh1
5a/frF0xRtoMZmpisT99uPOJ5XHxKNVWGussno4rV1ho9KEBWmbpKam3U0bWLun5
Ij4ORGJ8Et28cd/ehylA1zweAt4aKtztqxwsoiMruTnpmrwmiQ5LmNcxL1chNgrG
Pv0Qh4WViEU8+GOk89QxqW6yrR4+yge0mfiv61D7XnVP2/OPQb4G+eVtjnh/U8kH
h3tRA2hK+MpDrl2JCtBH9zr3bIWHlRF0dN5QetAuajQgJ7kIEdh19XAYB0pmz/R0
AkjEraOWBPcbcPcy27FG8mTwkF6ODOroQzjjjb4HRKmgdt6FmRLkIurEc6WZjSdB
xc92drWI/F5pzLNViKptIm9ui9Pc5IapjcN6kw0Js/Qr/2HXEOapvNwtsvUgoX69
eUWlJQP04Hnb9p2lrb9cou4Oa0YaGKls5SWrO90uEStu9I4t34A5sUAiToQCRizR
AFNIzHjwTAdUvdGAMGHJ01elp6jbWUI6Mlw864fWg+1gXMJK7fZZrFVl6kSIIfGX
wqZ96TDXPa2zw2wOkjeujB8Nvl7AKTxB0W3zw7dd5PVRAnJKMsOZBg5a9B6HjdQK
LN7zzlmeHzj7fRwX6EaHDr5QyEWs8+QaP6Eg/hI0/WnhAsLiKesLXb4VuUWxbsw9
tOFm5dmhLiuFXYe3CzM866uf6Hs3KKO2A3XJNqcbJt+rUSxKYQyZ/3LjG6eEFIu6
OdtahkPhozq+MsFb0ShMzymFM/iGhzDpS6yy5BEFtCEVzW+qj1C7OhlWyWhTYl/X
daFja41qbugnbqYK77/ytzaXQuq7LFoWFwcv5bHzEnDnBeuVB+G4kdGLv6S0SxMb
ese0NmlGXO0tFyq2KHmr79UC++9X1XKUObDu8Z6+hX0F6TqZlZ/1UIJsfV1v9lp+
7zARs4Zj5RFtaPb1vNBsRsbbYt946Km++UClaLDQQchX7k3lbujZ9zzK84hFZrrC
wOwNPH7LQ4ysUHdQqhU6WMdhwkYObGr1cECTTozmVkYFZJ6AKgCGbPQ8boQ4OHq2
ibnqMvo7VVQwURkIroM0DDOMBgbgVSrXD1l1jrTORu1DyGIWlS3QM38JHMkc8KZ+
zTvUdXeFBdSRB5KZ6hFLCOwqLiT98g0fVKcRDbnTF4kFan/o6GRUJEY0UOlDMh4G
iudAmO3ZbCceL0AbW8Avl6jj1KBCqm7Dg7obxWrEFJL0Q/k3kvh153e+MU6Wdzw2
lu56tjd/ZABNDxf+D+agWR9I+zlR3PwL/4CWQnf0PhaeLT1lKLmzqYUTtaItkAOs
7lDG+UT/mAPa+KRTpWhswJT4T5zfy+4YDJJby9vb13pwkW3fOTAImZuQ/XcEPiXE
htVD1KbAYqnadq6euuCJZ16H7jux3AzanDhiv/T7TXF2A15w02MZZFyhzxhLc1WT
YRLYBFany9g+O433Rooe5DG73tsrtiWgWUs+yfThpWQHd8t84F+rzvB+HDaXUl5s
rF9Ap3cRMSjeEuuS1KX6McsYoT0VyrS00Do2Ql9DxOGsUhplsQ4xWpnRE6RTyWqE
Y8avI1iLaosRVm2Q+B0d0FEiR61eqBRpuHSNcXGfCWw2aP8mpWSfw5DVusPEYj9u
w21XM6YMBVwv5LQ+oOphwBqWFyHgvTLoQOgIdrlokpCrLaTdV8Zw+Jule3saWPCJ
g3AbiNKkTLgxAEQ/4kBL4osCcnaIaZWPdJxRjjhFzBIDAlDDwwlTKUt8RsLOz9R0
7VDVKIpg5r7R1Nuo5oP1I8gJgl69PTX7TdWzGoWxzCcHTxkll2DjIyWwvxllQidC
n3j00jqEBB5S3aHuYp7kgXCHNc2QdPfzhKuZBrCQbZVYuaxTGew2F8I1iUFg3kQ6
GExSNNz7NSqYWhDIVc/gAnS4rZ9K9F/ao1TQyA4Ny0ztdj/KGV/K4OfCDGi+mO48
g59XtKxRMF+B5T4/3h9eAuCE5QkDYplgmsq3tbiqbVL+BBKWKoPcD1G6+t9/ygnI
ao9svJ940mOtXX7E0yGY+Kfgpva7VPjB4OpC9A9CAgTb++d0O/TwS9fSVklEUI1Z
csMVgIuPehFazBMJ7XX91y8uaP+zQxx41pVorHtlCx/SRC+NOcJo9qP04rRmvPHZ
eXotCFBzhxIpo+yycwd82iMKIr4GQHWeDiKFH+Tb9Fas9DHNdbwW6vcV+F4B8rmr
J+bGX7bt+r7Enl78sWtYdXziwbMaWZ3NlDygkv1CyXpeYONDlgfhRZVN3eXHmUyp
z7Qd8ulvlVBHGcHO/TYY8xDuqwUwxoeILHmi+pHIMvnPtgj0nUVkGC9XeYZoXT/P
l7KBzxD2TUz5XCLWHqvWZ4MCJaXsEKNy8HUZCPQ24ZgyeLf1q5oaSHfxTVRs79KY
Egc6KqcI0Ts51G5hw0bKrQubHNEA+nlFHV2AXbXnvUoffqKGdiG6ttmLVKI1RA8N
H7glzZB1qJA/ZzbeggrHyd++mUoAlIElZnjhyHKzN9PsAGyRgVCzRVbx+d2VdNYB
B1VtVU6ZrAeKNBfJH7SGqiEmswrtcup7OBNRpwRaEjyTBAyKQImI1GbuMPxhKZQi
07QfSnuus5Vhs2xldm0e0rN6nuPQ9SnJi7nJ2xzFOsTz/HOFoZJegcAn66fBCsie
4CssaeatxvK9bh8kKSOx2nhNvkdCtMgjw0IPRHprWu17/eq2yX4LPKS2mu/+11rZ
LGuKGcCniOjyZVab1t6zh2yJp0M1Gm+3b3V54AHgCKu2vdwE40KtR61fZLz/1/4e
FbvlSzWPkh2bghw7RQ9yDtKgG2PSLrNSSxGEqD3x5e8t8KSOoxdjG1aTipkxjXzV
iNLxoi3U2AuSvG2KLJTCTam05zgWbJ1MMwep+9WKUkHMytUDCB+//R41dKcXfmQY
bUo+0pilhjk+G6BHfkh/AlbdTK6Dts0P3g47F1/w0PFf7QZPwxvu0NWBRBA+v76E
H9qNDkr898hJk/0AESfyvBqVYDGYXEAFS4b55L0e2It0UVQipMHHEpQuTCGvdmy+
2dPmONkqA/78GNvqRyPvtOU0cFtghBOnItuGu3Z+4BpYVkYRemWDrw3D9KHJKsBH
SQbxJqvQzYfKqX4WXsi3W3KE0YUz+E8gJkaH9qJr3hJEyt5WvymTq7E1zbZu4+sn
ENaZZmz1YhbIVtxracm7F/6VEuKuUQ2c1HeQJyAvT8teQs17kiAfxyV1eBG3ZmQs
X83dd7A6DEuD/lZvaEEC5+eBBtpqBqWAzIu5tW5MhZCF1z8dNT7KThZJQbBXjnBd
aKE7Iq2IJnxLQHhat+Zr54POILPTY2ce+2eC6uk83+tkflVEKJoydHE4PXCD7ejW
c0twcTQdaZcHZCNeARPVfgQ57g2JG6WHt7guRPK/xN8rne+hyU8ysuY4wiFNnOkY
aXIqCfG1dTt4wlVo5KJFCFpAG2moTsMNvzsLfw0qxY3L3jOIJYqeAjJDdeZ4lLam
KnmesyfgPRezzI37YW5wBhchJJRbL4Bx8/hYxlAizfnBcA8tjcDOFRoHJXdtYu8p
5dg4lnz0TD0aLNr/sREYpRPMbfAlmlW87bqMRv/wc0ND3eXq2Chtr6W3i9l7ReWv
2USygh/h0PKHRimq1O0lrrdK2TMH9ZBigvU9jKCzjyggSqa8Tiq3SnUb/2eWbQVR
DTo75sW+nCZ5qmZlXAPWUywPx3eAyehycU6td1pLXObTxKFe10soEO2vNEn6ybZm
DPFFf5thN7bA+T7WpJ7WW0GG7jK9SaruCb82C0DgxWdAkKhtB8IzzZIafvIg/Imx
jrNuq1Mf3srKbVlrrM+s+LWayWJNac8EaEsXL3zdw4v7kvuwFKhE2MB8YsQfDuNx
J+YVYQhvRRCKYUxWMA5hSCnUYwipfx8Oy5+gbI+xSSeQXVvU84gyu4LyX0hzSK57
QuJY/WcF/MCmurjYJ1aeT+BM62b+1PP3Arm8EzAEf+gy5X24Xx2J9Y4QLwbY/hCE
58OmUQ70pJwsekSoUPnmmuDcLTgI8lcKk4j9s3ZF4BZ8knEt1h0hb5rp+PJmGoGC
8v6H2P/BhK0oe4NX8PKMHQlc5fnftS+7BTppE7vOt+iQ7fHW9prMibANeJRG+aGj
dcPBCUD/SHDYNsrAHfi9Jc4CbvusnPoy8intGBTlX0sJhWW763YNLTnrzOlFvT+9
5tdGGQ8HySIH91yES3qUI27rewVh5IgvizIbIg/MUH2mleUBVX2+hSTqIz/RPauf
XKWhfAFxYMWKxk4pUHmZ8MXSyYQaDX2tBGyF2t7KwRCcY6ga+NWC925URpWKVZ1j
JgRv1dV6U/lUkRkdfLbTKt24L+ZobNNycr49OBVIgPisSmUQ8BBHB30BC+C214mC
hAhdwET40W7V1QFHHjut+WN09SfFQSO6EZdyXLxHTTNLBcqPdA4+fkYeQwWVMeOc
w9cJUC2XgAtiTguL/iYM7m6ms3voiClqcsu0NHikY8UtvDreOrr6Y43IVJ9DEYSe
zAAZPrzNsE01RwrLZunF5OmXKcqwEtO8qFOOxI9mJuiQnMT7IGDKmKeAH6F6Fc2a
9v+RXq35iYUmejbFuCbMiOwqLsANdxQJDrnlmdyI224SXBfbwPow+DCZJ5lenj2t
FgmoMZxdY1kTTobpQjHNWiUIQfbCzlssHouUia1aG3ghdGUuVFy9uCHwB9An/mib
zPEiVxr5j4GOEe9DwmeTFrnOhY7kG5JftcH0KV33CMewXjnVkKWbnZZn3vpydO7/
ncVN655IA6bf1OW8+jgrvZspKiZLLb4h1pSSj/gTb2egXZ+r/OcJTn5Wo5brrmpG
pr0gHOsvJgIVRiqxtn55RgU8dVF7xxbHGMIZl5l0FjjAeeH6Q1OWbl4ku0qb8Zry
XL79zVS1KHzKkqdEimYHout0ojLquGoLdHvBD52g82I6dpD1Kkoaed2dezG1ssF2
6JnnI7CMBZUIhWzkA6chVyzftSkkCAW9h2GW8XOpqHgEOybp+uIwCmTMbdTGasgw
aozO7rB48jouU3qXAJ7/ZesVtxsQwS6w1z00d//TwiLzMjTGiA8Gae/bEMT57QlW
6+y6frefCmUBOrjgWnEfedi8KGzbt5irMdDlh4OC771MckdgFhP/IzFtXtBxUIf2
StTrigszMKvvlGL8ZsZNnY0oepks/I5PLECdiy6WFbbX4FnemClebewhgxQBHpHx
RjYnMPX++Mu/WtHZpdZ5Oqhc8ZYZPSt/VcITncmmL8ubuF++dcoYGnARNO2Qu1+O
HqnmeXuT+lvZVmfMOEFHGS/DxfTiJqTntJyDd+3pAu+OShk3ff5En+ta/yBCaVGT
zGo4S3j8QjT+fl4pW8guCGdXKZke2IP+JFV5zbHXZaO8EAfS+tO6U5dcNrEeq2M2
BO3yGooNBseBs4mi68e2h/5yNOgLWxIaf6ttNDS2g3VyZZulprBvgQizD0RSfLWt
ttmdGHw6MA+V2p+1FKHdY4ADWpdQC4muY/QdYxTSGYhoIxKar4hDaeXHh67MCS4S
JeM0Gl78pHbPgTBPhEYGDTIUXaMC/e3vpBGREnaUBq98nsYykfSJZUGohvLd7xk3
8zsh8bvCPJcHWkq5f9NTPX7ieib7wMbDBw8t+hMGyg+GperUSFnVH2Y/pdihoOV5
nmuPFtXcEti7m/RfNoDWX13cBD2mR1XAXqr92l9690zcQEgaYM6AYLQabBhewOni
eVqWnJd58kRMq8WEYSSoSV31WxSIcpAQ7qYUApjgQI57Cm2VTppJhZnLiNyZ38lc
r3BnhT02AKVG0q/51OeN9F00A+eENJ47BhFMXY5nt2WqLXupAvSsI7ylFJv5R8hv
FgGcSstA23RRZLbm5EHAZdiDyd5AccKuI0wfcRkQExaEoVfuRMf6oxIoT5tPHd+c
QCra3dx74rZbr2Re6M5om+DeP9ope96lTDXbgWnibxAQjCHDivoMfLwXPAhHApqT
ZjOroL9A9T8wQDCMxZm1xwWdHmG6FTGn41w74EoMBhhlhjbsHz9mW5VIxKu7230W
fZ5IvimWZbKR8ipJ4iti2FupXGlcRyxSuJu2SMo9kKHBlOZglNcuOggdzc6xEeAr
t/u3edZ88UmGS11nf2QvNCeBBvW3Nb5oIS/0AAZ+fUKaNZyVU1x/34AYdOTTvBpp
gNzmm/5hOSLLpsqiswXQttYJCkBY9wPOg7+OpdYeB9xrZkB/BfXzNEWwp0g8VlSz
vFWwukZGj4L+lCbG+Gd0dVM3MmQN+betUtqo50kXSJ7K6QDkHR8phTNm/0PqIn1j
ggyOYsMKB0b03mVvrru685cnd5JwnG1V0urB7nGiDygS+3oOK7FmJZj80vnLPrVS
6AioKIOLFBHN+GcFQTu4P52eLv584vTOogWrWMwAKL8hXtikHLNLtBYoX7x7NHnj
uLTZ0hg/Aa7P+yBM0hk4P216dYtQXSCvrvwz5EfWfuMM1kIeO+MDYH3OT21K96zT
vRzPpurazATPeCsqxAyK40TPqjbpigx4XzPpM/ayrucVU0ABvINAd2/a6GMU+dIj
9856BRf/orCL9hLvqK9ffJ50jAyr/M5B2bYphdwIYf9nTxm26FWOPuzQeiYay4VO
P63uE1yBgYptNg2b4miA+Gidnotcm+FnD0O/h/8et06zEDwqWkqwoUKKcYJD/Q5T
Yr7YR0EfzuZCnL0pJVqmgw/HWU9y2K5Q7mT7IVS+9ywtKQkB6KTOZxD2b/VHj6YY
MQHJzZkvLyJSw5SFA6md3ljY78vUs/xFrvs9/CUcFoFDlVO+7OLgp+uTdXXZxkOV
2nN+W84KaXaM1NTfk3hPpPEK0/U2JwXSttRU0j3nxL13pNxM8x+Wy6YjJUnzKeOS
v/R8yEejV8LFxO0xweRA7Z7PxKMymrbPBRpd26BOy/1m4xguf2XQzfdFGAn28foD
boxSyrVCCz2en6DmtHgyNKBuvOcDnL1trW0D7S3iHh/GhWmZ2Paw11+jFhunVY9t
L4OHj4JXsJMe0FnN4d4qJJmfkZL7hDVQ2pWZjzsFOxgOT5Y2o8GIKoL7umlsr9/8
INPh9aW9C+mmCSmyukX0fyKuvOsoxbSg7+3gYz8m0bXkUdfTQRgB2aH9blpC7ZZu
qSRfiSBq5vIFCPxBsa0cTJ8ZbjscXLAyEkfdgghjNXRIstbeLTafmJfWZn5HL5HA
hMOm+Wlv9d3XmgZgbMPrrsAayXF4HIBLLgkP+5KIk2B4a8jkF50HK6GzeoRmPmHy
hr/GKPdT9fom7N97goi6obhfk8S1q8eK6/LC1yODCZM3nT3uaI2RATHHaybmDvT1
rNCz+0qcbm8CNpIMRGr0kZye6fVMtP/6Q6nsxOfjorAo8g3ngeohtQ048wD3oxVp
9CPa4X2JnyIje0gNZXVf1d4Y0OKPSaam0th88dUuxYgB2aXV11+NvxTdzg920JxQ
XwAIizAe4MSawclgX4rQdLXEEm+A3coKKlKKIqfEfxQPMo/GkjdrQnuNEwWcvOf4
1RGE8XyO+ZvKRzpm0hOxa8yYPhk0Bnuq3y2ZmDH24sP42zkDD3roCJnlkjE9rRxa
1b9wFFPcEOXow7ghmgCYD/3IXCQZlm4ZYCVP3m/V+aGCeZFGM8gNZDcptc95jUsG
DjIvIGgpUa3Zcn/4hMrMZe3G9ILDXCb/4gdlzplFrr2MUPRWlO2Jb6A3D5Iop5pP
LiVzLoAsyZdPygUY4GaW6vzDCJ7NnZdd31pGIvByFg6kac9NgerMgn0yC/AFsT3T
321gJP4lX1xZAEFLTZUi2fXUWK6Nrxjc0mtCYHwHthD8daA/WAkbtJgTOlMCYEYa
olr9WaPDjLDn3EahPrNbMiKTyC3PCAaegAHRTH7WQetdcrRDijnFTWBSkgFKk0wB
30/2NdsOG3nzmj4n8ualQ3Rq6mg6qhc2BUDDRaCBE5KJ+Xt0egK+E6TFrpNISft1
to9fX9BiJath4iCJ6AodqNwQ5q8E3gEF6YcHwSCHaTYOkMx31GeAHWHKEByX2B2p
5JI9U3EkPz0ssVfAKJR7B1FcHYObDShv20GqXomk2SYkB4zFuJ+TQLQ3TLyQfPc2
4obks6oU9m+/bO2Ht+02k+y1u8tLMQCrOPFLNx6KlV8A0efb1FSlf+sz1RoirNTd
zeQsNrlCmKjzRJ5Ser/NLo5SYMAE/91+mtClFMfxqjtzK6Fxryu7/CxHMpH5R3x0
utY2nafYHcdg1D06L36VRJ74jb/Y2SMJ81gGLCaYyHMhzls8696KMHo9h2uw8iHt
bKuGo2JQG8Puewlt5xq4Y9z3IFSXO4mRIbaWhZX3DTuwnORSszJ2AeQaai09yzxQ
JhBUrr6y7nmBE1jgb135k7O8BBUeufXlee4yklhN9VfNRdu3Fz9oUUczMjduJjLq
Fl3biFpxSRri2LZgCy+HhPJuGEv70prpECw58Lk95P4M7L8eQUf1pCA8LnjHZHl/
bXXwKeKaBbseKrPDZ8voOzRelQmK8FpN4DPbmIXdTh+f/vCa5Qy7GQ8lX3Hwg1tJ
foz6790c1MCv73x7BHBRSzSWfO95hFtPIejhkVmjT86vVCelncrtcVkclvP+iJa1
aP1GU37uZuoQhaTu346JXoG54QZR42g5bMpJd5q/heHzuAmMKfNgSRD9qol60gnk
e60w7y2/gogT8ugAPLtKulDGuPXMdxiN/80V60tJegKvYRcaqCt8eIlrxB4COcyq
1/DXC5QNQ32HOL6jZgvjRI2pCYS+x+zrqMccqqGlz4YmS4KSm7H4kyhTjPZDaWsQ
9g413MVdc81/lngxlH7YgZwSCINGrhjvpgTOzUFVlBZ3Swl0xF/0G/rKrGnbD67S
MYTzJGK6LYRhZyRN1aVbysQXUzPlC+cCA7FGTCb8vVxcp+duh/FAC28r6lvLcUmV
1H/FUzniHJN/S4bpdhzCN764vUZWKRiOEDncGYNTgcKJCD4Jy9/E0nkO6x8VvX21
4Ih83N0Ecf60XMDh80fUFd1j9BY7djbgidh1wCTPfISmKEiFPJuPV7np+CrVQzgj
P5VklrYbTSmRb/3wMgepIuoRwnkSQ2G0a0EfO3i3av/FwUJiuTIWqmpKLSVHSAoi
5zGies+NqE1SSeOZFZ24hyDqQEbJmWECbBB5Pp4aY9PFJINy/QBSLMeUzpIt6N6T
Ceuv/oHqPa4vuFgjUg9UAwZq0vwqsrYQ/E7Tk5EywCtXNnDj2F6yqKwlMg8Dwls4
NvOODcvqnIaIEQ/TtAQY/EbWaFcgxHdrDbCIYygcgSBhDdG9MeZ3gjCM2iCP+ec0
TtXtgM7KSiaBdbRRcdP9ZTLL+MplIRol/0w9c6zyQfwOgSpqaS35J/ZdpZHJmcD3
tffl188yTKvResHHJkvrsvnkuelzHo2s8Yf/B8Kt+FJL8GkroJXRGEa2hEoGSgCQ
0RUxbsLjzRbAc3NgQX1g2WYZ+EbgGSgsUtwJdsyJl9Hy/6F1cD5xl/nFMexV3dWS
E3lOM2taoFdDAbiKvVCyx6NzvGv771EFQbZg34D+Ns5HHPOXvv1nc5h3cNr6sX/3
HaoDTYhDQwRUv9flDiNUFU7o3Ei+888BKCxozjkqm3fbj3NmDqJXcfSZU4N4CE9X
JngM43cooZWg42Y0qs3IuGYcWRm89DRYNZjqZCAos6lH0eOEIOxSDoSEk2gySbTa
BG+slWKznygkwMRjch1SAKbUTXVWps2UPOnGU61j8d0h+DbAGvBZowJ0gzFibDYC
8R8JTLSQ2U8ywjdYslCDUxzMzJqdebik12ug9S0K34gSlDx6RCI4zX4elO/UNWlT
R3lLlkfamzktNw3VoLZOLGDHrStQL1i1ePnczA0Y6oolc1qqzzlLXlfH4jOh/gV/
teyLANsYvlsS4Ic/d+HfYaviWoch4emqworcgtIB5x7Rf79tyhuEq532hIoPV8eA
WH7vvtstzdAkqVIAYfngVeg59e3/XEV0ucNIg6dkBBJVKfV79x/+nQpgZICz16ze
c7CzRv7jLLzce5OQm+1XyWRoljvPofxFKbvfs8rwT7LMm4IgiNeA7ffW0xe+PuM2
McxOwjRfzVMaybNMmJpAubRD5KIuU31ayQ7/+eunzry66BdT/ACU70s8rGlbKF9U
8AmvcN1TJZ7ITOWFDanq86mbBFyZ2ByGjiWqKsgAJ0ivy/AyOHvGekAOyNGz8Ga/
dv46pFwinPNFvrsnvkkLEWEa/iWvzoo/FkWEQ5Tt7rH27apZ/Dhd5mpKnw+ZgU9S
4GLLaGKSqzcXY6RreuH7KqQuIcD8p1LjvsPF2Se0JoLqqRFMpC/OmGFUhwN9TExg
IQdQsLyWD8ysAAKLznHrrfahxYJWAU7/FM+p6yQkZL9vT00b99P1TdcLwj1bYwSw
6wYiqy1vcn+S/wW6OlpfZHneTReNlc2pRsYTY82Yc3rvJ4l/VGVo1Uux2AzwMYif
HaK9XErLhzn7INzXYJ+cFdP5YXnKFNB2mJzbz0K3nArB9kH5PMgAhPfCPXFs3bzi
kPNUcl7inCRnEwsOvmXa99RUvSApe4KWdVAP9WmajWXNOyrr4pEC3aeexi4Q7feU
q6Jy1jWmWmNKh5uZVO8FLzxzRAqDOiN83tqQTVvxnnNgwFxf60JAfTQq5XctI66u
D0an1tIj+XuqKqiKegqWGTllV8J2blgb0gaYbn4m9teQ8rNqDyz66TtCHJs2cqEi
1Gn2HKMLdrH2g+x6j7hWz6oZsuC2fjVqSNn0DIn3uxpEDYaJEKNP6PlPEprbIgN1
oDUtPzcsQuMID45oWU+56pit05hkNk06KUudR4uVeKTwzwtoaZWvyncbYzwQWkPc
u8lwxCnMiyVA6pLF8GDwOFxw92FZOMgmu27pptN6P1rXziH/S+0qTT51PREgoPDG
UIX5P5p7kC/tZIYX8xreriVbP7ZIwLNxQwGmwSVZ9ndqpGEVx6hpPlcmja+4yNtA
UzTFYH91Zh05n/gAPvxtVuZGglWeeOht9w7jOWEadUUca0Qi2snZOjnbKqbaNbQm
0GFdKJGpruQPb34mhssRBA4s1ScuveXB9MMWxfy1aWwH8b1sx80rrPN1bgS3SA9o
QbueIAgF+/HQ5319ai75eN/ako2q2O/gt89cAL1WHS9u4GTXBQwNrphJ9d7Kks7R
bJrLdFxcRWRd+21G3o7XaAOT0dYgnnAL5+qQuYCKsAoahg9Rf60B8vUvFSZpNOwu
o6SAP6eptRDgWT1B9+TkrfaWOwybdGXO5MBB2K4byfgYgj1P7iDOUkT5HTPeZrMs
4S3xRkJ+dRdrekLb9w8DeQAamdtaz7szAzEFhCNmpT2ui5V/uH/fdeWqRu1ZckAH
5jEq6DUcH/tDkuzvpI26VVV/rs4rLqzCJkjDHd6BKKzkUFM2/NnIkGmO8NclSh21
pfgQPd2es9ohyf7AXpa1o4YpYKBrhLGEVJqQTsoBuMoG4O4rBFNUAgkZo6lqH7vl
ds3WRQoJpZB+Q8tiFt6C/KUqGmTQ3g/bBomBo6L0T+0OVk6ptv/kFANNo16jVBYt
TFt1uKl5ktkHefQS6QCElfDtWZyZuBD8IoAEPNBJ+DlQcC7jm8xwr3yqUk7VcWTR
8hDyAnHPdnfHRFfV8Zy73ifTIQ0r23QeFh47ZOemBGAGlS6A2JikXYGwbwDgBHLK
RRiqRaUUjxx2axLNCsIl4QZNEni+hbqkkbtaGzip7isrFcCLqRSx6m73lOi2IBon
wGupX6guwZGwDZLAWPJzoVNwhspoXHob00HyasZQTByUERyymjuBGntErqUEsxui
5lMncd36ibJkH08lqBhz/NaxN9rRNSRd4u9c4WgDeizihF1aAbNMqUGMZ4cTOMoW
1m/ocGPKsbUEqQsEIBlIuY+Xeks/bxc5svBT3kwgkw9y9xHzQm/6Qh0mAgah3bm4
D1kbskwd0UPInLqfG9Ct+rcrncVfYlMajDAIGDiaXkWwcS3PQMX+beDbNvRqnfwo
+P3ibZKAY+oPRBdE/+WTEv2phsvEQHJ+TgsPx62Jxzs+psbWs+6j06ISy69KqboY
8kGExILyA0nSa3XqzAy0WxBHmsq7P5hJ2bE03eWSmw00md2HgUCn9SrrtwyIIEKg
JMsPkgziTypk73FPt7dS5JKhjOvCTXDsZpS39KNrWTSEimzO4xCxTEcP2sjdh6X3
44hf/QY0qlYd8mr5WYTQej94XB33kgB1M/oruXG1I1cQsBq6S10u/HiuwWPLzdqB
mdbtv93mcLd8VwX1DRrl95WAitEFkZqU77NSnEK35U7woDtg01m8xomGCeqmocqZ
QNKyqZ5CQgNvbgb1FcciyJTS8P318UT5l2RZuIjaxXkuwqzYQ1+R8S7cwY5ABjMu
h9a5kGHpvM6qS9XAIn5zzz1jYKiodNwv8xfezYO+PnSMqKy66O0bX+CBOGi+HijS
+CQHye0CuO6XFvovPhV+QSEUEIpFpZVAB+FJ33EYTS/t1QJZAlXcTRK9LWPERjdy
QvfOypKuW7Bgeu23+u61sJ4wQBIFGlYfhat/MqjCPxRuOijiB+3573hyaoRL9rzQ
dea7bJn1rHY47zId5jCxtZqH8oReM6/PVZuTI5zab/wh4BGl9E8K7BD+4+ptUPg1
AVjAGjTrGZY34mKwpkBul3OgXetEwxmlBXNn8dF8X1IPucDkhdRFqpVLGHXL33FH
KTEwzHRUYyUQbBgL91/tcWWnirGHFIfCnecQKTxKDKLBUY9uvv20LaB15q91urVi
IJemIugaoMZZwI+XBnMGjgOlme8ps/8WnF2AvSfVDXr6cRTj3ntTiphoXo6nvP1n
cdOvJwfTybKPwulX/EwPLunnzT+reHdnvJqpYBauOsONwm14NCWP18L9iku7YbT9
5cHDMN534HR3xBPxK0eIhxU5x5mvTyeRb0CwOKXOxUINqvunylJypm9ygdtT4QU8
+SJg2gQ8zAA5SURk8eOBVwEMZH5TfKoN1MrLs+djXUao6JN1erCgSxa5IC2WwG2L
6RPIT8z3bidNCYn6s6TImJTQXlArD02/zapcL25hUD/yeHQ2VInp157O9GRTKEKV
ygj/ueDfZ8ia3akjdP0PPFhUvd9gOc6pU+dwR/nc4QahFRAMWNnqSHZoFlh/QJ50
fXMZoFmW+Yr8jaOcTDHj7qqFB1mDn4/g4zZ0YjzxvEhha5ATDfN51Th8b0LGGVt+
Cm5Fix2IbcObRcC666iqeWPMvCkFxv1tkt72o7TXBWJyjAFAnewJ0e5fibkQN3wp
7o/yrcbsl+mtClDly3bgUcIU9dyQW/CINJSJdTFi/1/MzsTDgVKiFHzWPftwvXHN
tnH7Q9GyzMYz3Uw6kyOxf+m1ZJTkNiiostdpGtZjC4hY6NGXHM7XfGpySflJTqwa
WqT8aDB4QygRZatVIhTcVBOc7jDu52XfVtu/MFNyRHOvn2fNMe7fAMo/AFFySiIU
JJWeqMOCgKuFL9VvdecVD0vqUVClI6ezb3bzTyog0AqpQY/4KxzJCqENE/lZ7rqD
UacpZ+6avleVf561YUx7foBi93dkUTeDeznZ1cOslG+RkwKTyW8xW39Q4OnaHewp
lCKXEteXff/sU+woTUFFu9iWdyZdFeKhwqNJEeNUSRStEsTaK1IMn/yxsH0xxQE7
huTcU51HKr7sV5beJcVvuLt7a/W+4uhV9mLVCa45AxeWzOKsp8xrfXj6AcMiXjQQ
bPzNoeIODPeKnZcKk6BWv52JD3cjhxPdP1xf9iZT4JWExpeyse0J6mi7sD1lMDLd
fzTJ5CrA3wHboeXVt9r7ZhonN1VY2bulNqrsfe14sI+Gh6870QKJ0WP0PydQ8UEF
hhYkWuP2RcqJrnXeY1s0Rs/1FUbBw+FgpGHO/RvWiRlet7f4IweUSVMZowjuR2uc
/Zep2F+ViQJwKvNwHo6mfLJLIymou9lf8twdVozSLGYEvj8SvwtULTkRl7N1kDuA
wrdUqpX+i9VFXJ3WV35vP/76j7u+UYJlxV2yQLvUUWSu2cw7XbUEFwZx9Ek2VBlN
0m464/0fezTqlZPPt+FP4RP9XPrv05ahxW8sPfqTT3FdQCrwSSFrpjS61nbuLa9c
Io9fdwBNPTLF8qi4/ZsO1SFU9MksuPGUOttC8fjDVxuw9juB5ZKgCsq5ERlrrc0f
NyBbXadSreHUOiyDSr4hF/HGZoe9rJUxMPNWs47uz3QhbMc26xdiWJynz/crivYH
TO3LDZhYusCQhzIhMFd+5OLFR4YIHjkls8zT1hhW/IEAwmutEAZNA8GfYxe1fvXq
mJeBn9Trca104a2+pmutlaiBI8deFWjntGB+Dq/cxVPq0wA1h6WfID6llCY/Kz+x
OJIDGLzCuJPTaGqriLD43VTAxqehDqU9UDIb1mP465V0rq2xOCo7SpsQbf6hOCgw
3Fxkw+98PS1Q2uHRPHRu2gCEVRYKw1vuYyDv61qRB9dfXFtBeMESaDx2s4Xe5II5
nS2apbR2BnzUdrIDzjwO68uQU5+MuePV4uA9viM4UlFBTegKAP043Bun/AHl1Mt9
SbkyptkomWMT6rUmaatYZIcUHzm9WqOqAu030TcVmaFWoHNBDvuesPXHBbl1a6FR
xSM4cnDH5V4sbQoyZEbmMH13PnoslR5vlNH9WrGbr5Cx+nhFlPKbnob0l09G+Mo4
4UqeyFTCdr0NNfr1+HN1bGl2Txb8EKfeudfVfVgGEQ3tDJGP+xNQ3xxA4yZ6Ahjg
OfOp+YIAdPYf3DZbxKmkQ5jqKFYHUXxgZZwSd6e4RAxQ2twPt3NJ7Zs8C+6P4oP9
UVpz//yWJQvu+D4pNQqOwBNBqO/B4Fi58Q30h1GYrsU9FJHiKRJleuo2kGktZlJ7
KA24G74APDa3c/O5hLZN05n1RPQ5JYFnVf9jXQ1/00r2iP9GkeTBFQ2SPy4tRoS3
oEoit+BqO5rZ5wzlbqKl6rUnn7H05VxqBxVqaPlwn2nJ1I53ZLPp5hu629V9O8uD
J+9VifXOL8ibxFk90qxo8GWs3azWVYGUvRvzGDdGon9zNAP5nXBoPq3An4Ay/okZ
seQfAigBDr0YVIljjEuydEn/Z93jr9dM21uAsYH/HZjlW++wt4YFEqoPgwtWdNRb
VFap3wpUMGRDWiOl1749doE0GGQKmhF9YSCoDJoIPBlc07gKnAlGwqlEVxq0JQUL
1tz7goktNDMr6VIPA+jMGKKuK3INAdKjkxzHqt6kPKiQo+ue+Andaqh6KYSwxShf
MnN+gqJiR/sA270mDfKvw7PWie0ima5iigRIPPULQQg2eFWhAWnw2Ld3k+YjBJRB
rO7yrb9Hz8CuV51GwZYhRAdzd29CoQBxl9+zDznlUhXYawpeHBrYIDwt2wSnRiZL
Dor7BHwUH+wqo4ksa/GE5xCjuRs3oDws/uksdD2ACAUZ8f9PAf5hrJK9GzJnfxWR
o7rDkxhSfnWT1RatksR7gqNeBc1JbubQS3TPtNE4mnQtTwm54k/iWE82Tlccq8jJ
8ijuLK3awFSDEm+zpzCq+mIJuOWWpdN2Qsuq9nOYvU+G/NVRKLy2qouVhSP50xDe
9PDem1iAivWqwuTOYPTf35d5udt1yfEHfOx5W1roKvzXqT65ol3fgoW9AxppjCcC
How45m5ItfLZF+WffnqHudef+0t7m/IyP0G7MyNMrhp6uVWDpbqK7ZIQLFLfJDRW
Mw4u27yRKtMybP9btINLsLYaIRGxbVonhCbrH9bYg/egHdq6+JplPow2ER0iESWE
Hruh0MnoxQ+hiHPzsgsIuEbWhz0E2ag2/TD35Gdvy9FSd/GPz8hAOdFL6KDcO6gz
WB88TClSZNZ2Zuy3mwHJHHu7U7EhI057dwJ7XYKvrjgLOf0Tg/wKAMIPenCigy3J
7+jI5vfhSikWiFh9hSO35pqLojRYfxYlHgZq4EN4gdvzyNNtSJVa8M8ry8fkKAik
X61m1iocGxmUEfUhgLDCO92mfCLg5xpvYq9QVo4vqfVdJqOfti6LB2mBwJSTWch8
wcPnZ6bUDuc/PTVjtQfgtjCQqd/em6gHsXxCHiMBhdubmbkuj25VRd8r32qGluzR
V9FVogZgRyDL8ZUUJolwEWE+UFAyi0jhtO0AOWAnyeVQQrpZQTvqaXGYYzu82FRq
MIVEg33UGvCo77ZeiCyjU4Uw8tlyohUZ6kLRqjIyo+dMn10rbXrr01KbQljjgtFu
+ZbVE1Zj9hKwD6MGNjGAglkTG0QwLedjzUD8L3RbZS7g/+d+EGPX+cSaFQo+689b
6A2ckFysDvfz27tZ8Kn06qIM3rEhHM3lEkcOe1Wx0TCGiFRjO+uEWqDTTg3Uax/W
52HvOlZgLB7IFVjLZk6d2aceft9fNSVoCTAPpdz9VePaEGFyon9sqWrOycDScv7x
TfgQbgsCXtwz6rOV0tepYGOoTqBcXHeVwA5Usi+Vp8AOgSIatF1VqDB+KqVAhPGA
iEW44oGNQxjsDofmbYBhMkDg0quCE5AdH7idqZfCWeY9FUsItNehvCZXUnx7qJt8
45rBrR5wa1nQFaXttF1RBqKNF8VHg+aJ8Hvw6GACxsZRN7+1CV5zKYNewBj/wKy7
hjiTwwR4KsdSGDJRjAKBhwCyoKbS3waXaAcESQHSjSt7ysBaeyj00rXjIdjblXDz
46HmtchCSmmzGY/qyrEnRATFvtQSE84t/DPzAZK5VRU5POZci/Y3Ravkt/QAtOQQ
QsjwgAhQwZPXWN09JhWam7IWrUByjHZx/DTX1qLjbFjA0NkMxW6dkJpJhKuy/c75
PX+62cl5mKX5XzesNgAI9EkJv+oRTuedJvo2b2O4j77Z8sWYOCqcVkYULong06fd
B+6yjG+n2gJzDCCsJbcaedRbIdtAGrfu1LmEzLa/BJ2TZXi1005goG6OvItTY0I6
DM5Zg3l+Jxk47UfP8RAJB7mf3rZqp1FUOieOKWnLJofOIKuzvQg+a91I6UIepArT
0NtXWpmpMQIlHUMhSzi7hng9Irx6Zgow5wTFyY9c7gV77Ne7m28cVPga2ymW4uzN
xkXjAJYbi6IUEIBkV3GdKcAi0NbaQyl4y8e+9e/gMTgWC7BLrOVf2dW90fNxCLGQ
aOpgs0myXH6+cNCfBKpnPjhm6SVzM+QC3sfRExCnIPTM6iuXqshipv3tD5++HJ1N
fHyYEud45AWGzB46jlqlFJu6PAWLneeQYxHENRpF3RVSQPQDP3dph8vaoA6oaVfs
y/5Jxk8rzU6uZ77TBAWCVaHb2Fk+JTOv3rV78CK78CN7L5XmAf5yba/cfKejToUt
ieXmftGDBYTUhDmsCIhYEJWc5uta56qg0kFWsh6VbugPivgOs/6jC5RbcPux2ueM
NcsZYqFr7UUCEsOA0f3zI4baTITdKP4LY+UCs5ZT5zklkuhEKh/mLUcy7F5i81xb
jzL5XrUHCZFKSCBjZkqaM80WsXNRbobo/Xx2pkgo6ExrDrAajE7CZJBLIDj9RJxN
ZmkEwsD+i7pVBTVCujJhkOiVG3TPTeNkNoVgAv7ATyfwMh/z5TYIyHebzqXOkz3l
pQZN/Pv7FITCCjalikamEYuBX6gpbiYgirJ6KRM9RRDgBAAP3z5QDt1byWnQJXUZ
RLck8Dg/VkVWoNth2lXm9/TnNrRM1SleI1w5aEkD6YgQZ2qDHWLYp/K+kQI98upA
G8QyFGqO3Q2YFqFnBAx5neinGALzDYAMlMv9ojYHpCPGVyQ8kuuemHZiIs5qcIfd
o+rsPzgyWhCxSpny0pkIHyhtFvc6xiOEVzhibjhL7PiXf04j/LaB5wYnbPCI58jX
k/xM48LOpTC4o9DmY3n9CCvJrrA528tU6nOkTCkr9Ji9dZSZth2JjPHXWXYZ/KIm
BjbiqEMDTDgP+4q6a4CyNsyR9p6/kJvOCNwBZteGcXvfv7cilDl25laLvCFXBlUw
vmC6c9J9NSMM/P/Rm643gXNuHRh5u7pTv/R6ppG4S8Wx8JU1lGMAvXLzA1voya03
FsnVvdP6SBqquicB77yi117R8eR1VyZb/bKdlVxS7xdinWJMF+0yCHzTiijfqvvs
WfNgxSt6DJ0lQ8QTqfWIzqoVAgISYqHmj9/KPuFFgO8=
`protect end_protected