`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzbxWtePNA4xLKWL+TYXD9yg7MHdW1ZcoSDFbKYqmZEkC
M0yd8rR7zJynZXBcuyvv04m553ncgieVP3KCdvMkqAiZplayi+QBnJAEP2F7+8NG
Tn17Z2JD0pFFMgElx9fQtfU/ASmFYu2UOXXeZmVMmRQpCHEyfI+nodoxCXc8DSID
Hk4zmf3jzysDJ1XK96lmfBNRQ3AVjlLdXMPwSc/3OiYNeO0UJyv2GBNiM8Iw7y26
JWY5mEToZWGDfhntN6g3IJi5jgeZmCQlJ8fklMNTuZqqQeyEy0bqw6fD7ZxdCxRy
BeI6nyqgODL/Kd5JzMKCnBTf3Az887jIDfAzreIiHpe6jBi+K7xMVZc4Jt1bgy2n
uoIruqs9tvHDpOg65E1w1uNnMoqq+QCJ3HQKulPlGNNMYw5FeAAizVPsBtDYwjdz
7jU61ztHzp8+JI0jyO2qmi0yjpx1sffNSPNXBM58aEXI+zwlKO6nWhom/BirWxLN
8bATQigWvJKVaMe9wzvBPOEWlg2oB/rKRFQx81L7KKF/H5EWtqZ1Z27YwH1ajrQt
Qo8H+zXQyZh2jsuFriFdc2WEOzNw1ztBf1+LfM1HsOZUkE68LhIkb0XwKVHD0Ugv
pHpsDT/Y7i2A1CowjkcEhRD30PBkWZpq0dRm1zhr5ZuYHu3xYa0yGWrzBQ46MwUL
VF+GQtTX3c71UQsN2GEcpjKmTfMQ9oZyYDpzW0pC+kBJVyJ/TyQwXtY4t7+BAVYY
ff5EGmVSMHaccgro997xWk/SLRuJuAjVhjg0+vPFf2FaFPyXVNDrAmXsB9VDpuwG
k4fd10BlnC9rnLuTd+GQPwfBOOXWGx69t7jI6vC/GHy2fGrQfAw/ALWK2MXdroc3
ovN6mGhaUYKujcQpOn2tqa7pKa6jhMCSyWJ98UWYZ/U+17hvNyYgWsrPh0oSn1h7
kSLYqXMNJLjZOKEBwxXzet7Kd5YxEzAW8mHrxQiy/d/f6OIwUZrt+ob48LbGuDH/
N9WmVEhqCmF8JPMlxDhh9ESo7+SqJSivWInj1fPsPX3uFUeTqd8CVPSqEoMZbndr
C592MnyfMQ2Ued6BohK94ZsdH9HDhEdjbdR6ABK30iFKt6Pkh+vILhpYnGRVeoqi
uOv6c2YY1qJW/MGdcPRGY8RQJvif3wP/KFjNyk1A4qN2bsvi3xUFMA/ngYwGLnqf
k8brdZBYNNkrxUncA8fPaffBB02JogeeqfZrS5a5RUiqzV4OQhaSa7pLaoXv9RRg
SGN+RnmbzI1lpyV6yfITBoot4NH60u4DVVtMQYC8s5HJ7wCZDp3pH44q9D2sWPS4
bm/qQX9ze3nVoNQjzrfu5MPdD+2QxVkbaCk6Zw9ebKt7UcGz+XSgKFXSin9WSLAJ
4Qkz3HZl77bWMiqsInQrttjIhV36/JlqpqFv0VAOHz4vFp/a0GRCtvJIf/GOA69g
3O2lf9G8u9J3LTSU2nMdib6sInNYa4AUsuLDy95uEEYLUXZVR8xcBiyiamYlum3Q
/dOs3Xs6MAQ26gl1OzNdXS+G+23nTjC0lxYB4zpPSSZOl7ilGJq54LbrjfiO267I
zYOW7JPTKHkiOqtxO6FhmQEvqbUikeVMeLWKLeVngIkic/CoTFXrTc0lfKaFNYiQ
R7KmnqI/bkP0Hp9FwlYhiz2cg/3vPwNN9M9hIYVB+Rtxo+ZsRFsBXZJRuy91o9nz
MeqfJKl1fMaP/xhOvRq/uB4WlkYNypjAlim+tz0Gj//N0ZvGMaV1TWQQXTPMX3a0
ADOP6Vow7hVaXUcTtOkbvzfrXR+nRItx7dNvf2Vfrc3SlrxMqlZaCGwW0vZRtEuQ
jq1QXIW3OvkPpX5zfgXvYrqh1Zc3RJQ7wd4RhjqRxpK7H+H6+S4BVtz2o29WNC6Q
q0l516Ghvh6eYrkSgsuNXhUJLKYLfyTZRRodwSyxvnjCNJlqZa4LfwOOX9zbSPsi
F4YnU6S7mjWNQaJ95k+q+6kullgYwAAaK5OhTOduYFM1hIveCra8aLkstCQqwVUS
AjGbicW84WVHtGgsVqZY3n/htewC1QjQQMEAUiiMg8Hu32KY1i5C0rD2+GxNpw2C
avtuLB4fJjcGYiYQ/LRL8WSEOS00qi1cgoby7ljd0mvLqsJHgYMwSsxaUN++X+fc
C7V0AtZcT/QnyncCR6HKBEk96HbskHJLDqxZmUWaixD4t7k9V8+Rjgn8LuK8lVDo
jiMbLQRHoWPC7wKDEj/FhIo1Po6RuB5u5qBJ+9tAC/Zdr1I9CNdamZT5yvxCcYf1
+WarKuFOGI26D73cxy8TvGJ6NSm7nGKKBre34uYvrgr8cCkWvJzeBxe0wX+DQ9o7
lOnJghNr7p/VUAerMAKkWQm38grlr9GgT7S49pwUaEIwJh+7KYnZfLjKy+ZG6wbb
b6t5ZYQlb4cIcyqSBiOtbAnIHZ1LK7h7PkfS+WJP6iWG3OB1E26rbBZruGSmYH+c
HcRmI84RoVY15rp6tbzTYlnLI6glonvO9cL0Yh6oRgbyALpZ/DEcoVa2W1b8BgTf
yhzhEtklw6wwPMlJC5Z0ZubVEqLiMeWTcYk436pQJ8jFyTQtoG4UXa2eFqwQ03b7
lvS5u0kEfbI+rF2OLHkHk+v2FJG8abdEyZIrHfU7lZjVENFktMy456bZi/MbIJ0+
lpZOclu3Ksga8XVDSEnlWke971O1PkbTrr3CXFlbV/kjBpvp8gWWKL5wvHO7bI31
pB1ji31/fbjbDm58bgKEduLpdnZDe6ag81KJqj6ZtRejjHGWxCC8ldT9phjJvEmG
XPTOm7tdZcUajlsPAQGo4sQY3FPlgToXIU67AEtkGOnzujXQKNHJt5G6KXlofoju
mNIky6zUloijr9A/zfq7LMgKXzbZC6EXLwlxzrhvUyAYK6M6cXnmE7p9gb69cVrC
+CrnS+9BixE8aoWRvffUAQ0yUzFDRXzJcTqO8gboxJixn95IiO3qQc9mcMiwDXBd
5i9YAodexX3tGV1zrDZyEf0bqMnzACNYmsEpqFxbPLp4JMEeUcB+AdfAd1E2psUB
5mq8zU/drRmEfX7Siv4MQebBTLcquTeyd2aZTG1Az3R4atOfohOmVzsiYKtiluba
4LX6vhPqmpmNGTfLYfeeN2q0TovcMTDmCEYl1fCAPzsyKkP4NMXKFJBI+Cp6lP41
qa6QIrUyX9NpwBNU6pqeBPoTu5iQOzyPFI/Qt8N8auIUb8N34CKyr5yPEy+s5D+h
iKd3on0h9s8gqHGLK8a8GyMpBbxzGNsMJjBE2OTJS6QtivkKzN/s9pzWMbtyYvcX
mnGC0RmSln+cAUX6W3uHdIqYrFrbqAeQnX9dvpKai4oq1uJYqUKQTeAf0nQC+gXj
0hKVRiTdhS0rchyc0A4O/mIFYzr5FsGj8r+S5Jqgg+YIxXfxd96lWzex4/WV69oH
rlqNaPJXN77nMXPoOUvFIbk0gjphwRGCYTWdFx/ZYUnucdhKwfFe+1z+j6MoawX/
gfsQxhgnZPw0XAwMrXffZeuJp+cdfX/EVvydadHPcVqDDPkMy7T5WSXHvkLOO/+f
ORpwcunOai8TbcTYVo2Ws5pSZZksUnd+6o2X1HHZum+fQrxhwrgxUMf9/KJ4xMsN
OGB8MJ+0HlEHOxf90WP8UnPgLB3yD+IBu6V/1Gwiu4xR0gz3bJ+QXu7o22jcNG8z
bJd9cmC38wDjxy2OuAMD6j8LZq0huK5QIFP2VKyizlLCZ1C9EpKtNB+4MukIhrsa
cMGnRsdAV5BlDLMgVB0DZzorLCMjjDJ+reoMmhVwz1CB6i9GZIaYKCYIYYZdbHJZ
XM8MU+jouYJ9LD+FzIf1Bq46KtVK86/2OPJsWTHxmY0C6pj8vbvrjH3UEVSG0EhO
1OjKdn0M302dKfi75FAgGDyXUypMkGohU/BHwktfHQ8HPqtoKSwWsMRTmwygEI20
G/u1YFisWb8PR1/1skDzS0jjFFpz2umrBFiGCKYy1Zu8YwMlDcM8uAj+52WpXk6O
eTq6gJotHm/WU8nmjLeDzBpukYV9WxF9cm8XbQCICwPer1Ysh5SghaJ94CMPiApt
lX70NolE9KfU4/+WxMgDu5iZaT1TKkXjQeYZafNR1Fv/+tj0Vgp0BTCcRbcIDuxT
eHBloe/ShwlySYBkqIxv9odm14FT+CXVVXY/OBnTNbfr4sZMBzyDAgwwxy0EUGFw
Z0R8Maa7mcFgUuuNHoMYyq4yjbAXv+Hwqg99gbrH64Qt2f2wEjgxIvMagNbphzFk
dDLsU95EtJscx+gUX6yHxNwUuRj3cxM/fvTMTb/XQxvkAI2NJ9n3jU88Xx5Gk35m
2No0KmopdspyxfA4trw+0n0qyjYlAXgwzihFZSFSYgj2lhGvuZqdOPt/mjIcQ/7n
l/stqIDZYV6KDhUsejKSsA6/uCOdHRWskxce4phTfMTFUz+uY4l882S0iMctbgzp
5tej7nnPJYLINFfbFqDiyVALzb+z5tJu/nIB044DxDnzddSwKzuFKVOmIbn2ryVa
XH8698OWre5qSGXD18AeZdEFYkbvm8GDInKcch+rAo0yY+07Z8NoiojcsSL0uIiK
O6CgzW+8J0HpLpfjTwO+Ph3w9kRzpZCusl24uBVnXxX42WsSB6Fg/IBLnZq2NiCY
tuDxMohLclaxg0oVo29qEB/D5vb/w3swl/OtbQQ5ENmd0eGo8yKBZGaC2cSXKRok
1fZyynb7Y6IykbEaL8oWWJt5lPsF5AO+l5LZAuEGf75NNjPMuUzfhhm42ud2UISd
LP8/w8SdgN+CDCXnEnvfJPy3XKmYejCzvtrduc8+0m+eChWv7BJfhZYKz38pN92V
+E6avSdjqinUi3kTD6zh++f7zQLtXGxdOs+REY/NVrgyXaMHrDFmUgLfz/d4L4E/
UMA/+lMUeq0DuDWnEyFUsxhzoDnz+3gNrghjYOiHJr922tm8jJ0h3OkS0V3zEPxh
ok+CcqBfa33jWVho59vHou9Zs7Bl4LN+XtGqYH1+wqU1O/4GouitODNmLUB4QNSa
mbpRad3JOyU3J32/b0NSgrvLEuF8Avb5lbnFKwAT0/GvImSnxQbsUdcAZ/yX62xh
m6dDB/XJWsbiqFBXoOWhfHrZNokxCA/hFO8unQ1YZNZ9gcX2ZhysqEtLOAqtsBI/
9XaM28z2WLJzjDgZb7rr18O/XMumsoNPWEXLChTaAK1MT/aI4tQHAOud8xECEr0a
JH/czkmngBymWSWDJ2E8DbyIuJSIYpnGmmO9bbW4mzGkIwuJKCQvm76saA7WjjYd
W7nfAkogFW+LaR9bZgbL02TcSbFwzFtJt9WxQTxJHd9E39wfNme+WYyPpDG3r7s8
0SXRLuUu+WnxVWi2MhlyUeSFZEGei4q9ZPMaTfEWKye66VRd5hRzIp/juDNub9Xr
f8+W60R03xm+zgwDL4VYe6g8ZTY4l3Wpm+IBE6zi24+sm1G5adKJximBPsxgx5JM
2blrJrqH4mn1E+Gf1YIHFcBCnCy/RAoXqjzS8MRjh/nMy6ogbad4A1aQC4SBjXKG
tVA/OxlKMVQExrFB6gJz1aCok7POzzlKto3SYgty11K9G42iqOaXsQ2atyuvFPOH
Uoi8G+AyiDHESzG+2t+3D9zOkiR2pPQuJQ3kWv2aKtOlhU3JGCbMnvaMHDWPM2AC
oMru/bmZ6ZdoLXbB8xCiw1eI3KeJ/O2qQvWCWlsQcx9rNYvaKpUT01THpg1NuycG
iKdTWHzReoFAsdyZImPOhfyAaLQlmT7j+nG1bp6nUlSv2+6inj8dE6M/q23UIe0S
n0q9hERRqTdx99SuJDhET4THd347TWGsqgSrF9Ybk2SWqm+qZW9XLfoUDPrf15E+
h8YX9PZZESmtDcZaWJzJUvA53adzDaXrPB9HrlVavcXQLYUX3Tqz79HY2lJt1Fux
EXj4Vvdf0uuCvHyAIQ3JsXtMqgdVlo9CBh8oLrTEF4ApomJlrbbRpwd7cmEpenUK
iMswa3BUjLN8q7+cePtwRGX5mJZ71IjCDck6sqV+gN44AKMxlQJfSWCQrdtO0hVX
o2N6rDtKNCkPBPL1tPAtzzitYKDGPrDj0iX27dC5kD1zZFt7NdCJjlmJmhnZtdgl
1Ki05ILwi0JIP7SCNExdxOfaYFsKE6YoEHR/fnz/Mds3V4ZjihsPnljuuQKLxHJw
Vk4IKpZn8pN3f//UKU9s6MHBAZpEsM5gysv1xS1G2nhvE4xYaxTDZ1Nezcmry+US
abgVvISAAx1Hn6Y5clRBPpnWIAv664O2cyAbyXzn90RJZzw6CVoCkCtgFqvPSvO4
tPChlZeXEHSfuXYNnFKo9ybfHTknQ2cYLsJvWBj5xg4+qV57RCjtV3d1gntW09vm
P9XrNRYXBmk06tQI7kMqSSl/AaYc4uEPm0BHKyl2q8jA/+G3b15L9jDwKZnEaBdH
zjHwUFnqZsZux8C8QKAPeYka4gx6/h7zkdtm0MZkktXXfEcpd1zIlui/GrRsqrx0
H4sWHK0PqvJ6wUMdAoa8dMfsJulKXKaouYAJJ6rQu3sekuNtqvjSDLrfo4mkvFPy
X+xf1WexxoQSRY9hQjgMXi3xRqj0zjuanXle7WxXnyE3GO3CfNs8KXtdB54/v3/H
CLKceRobrCM+54AHGkG7FzxY1H9MyABme55+RI0ek9SWCgVAV4dDURXNjutAl/pk
C6v3J9NIg87aYQIa9eGRNuYUXbxgWW/j7TZnUQ9Qv1i6Vga9pg3bNvx150Bsm/Hk
gkwnO418FAMtO1aL13c4N1UD5L1KYxDd7rg57fvmRuNODUbdNNJpA5xhloc/H0Aq
pdl+MCwhFK2Y1sKF2zqYAGMqe1rYJV72/bOMwA4XQyjLgTN2nvcogIR9AfWhED3p
JdLaSnRyX7C4QUpzisiQUIbEFpUxBWjNkrKmLo2ftjUziIVGErCfoLObeqF9QQ09
IoFzHM47foVMQLp9nNwlgJz7yrppyFz0IdDzLc4J5WG3GuPn5yzMONsZFwhz2j4t
OhEb/kIo2+BDdwyk9CW8Rz8trVKCz5Gu6wthmCwXb1oo4ljIndFz6OJPXaGXCdb6
pA6LuLxBgoh7Fw8nk5JCHga/kFC4I9Nb/59nbM3IKhhsImea7o+gcmJFfnhU0emC
BdT0fm40RG3UHYFb9R+FQhFUf5NRZKfRUbM3au+n5YkS79ooU5KhuXmXJ69XodV9
Xetej9mfRsf4GgytC+Hr4Ud4wun6NwAsE67bwFUkAuxtXK62JTJOJ7yh1CO5SeRn
Dfw6bJNUmFdYHbq3WqQnmvB2Ga1nmFxZGrIImVr7L+rAswy+h1+iZ9Rf75daIyVA
EiXPdkOI2Z6NALWGM8pZOoCBabpVE7wVMaUqpqAcvdJCK2+j/pQecVWmDt9ZEnP0
bvwQZG8EhcoJKwzpqQ38ax34Nmo7gVuConWmfhdPRHeHCQCfULc2pBYYHxY9srsy
BwjgjAAgRL3pW6gXHRl7/TmPlBasnzDrUauAWjdzMQe7/OCEGiWN76sfPVzDUZNV
/z2xq3oVCukd+vZHzAmxY101RPU4PHwnxUiSF4N1Cayw6MuN4B7LSF4o+ZocN0Wc
Lw6g2m3D8x9qsbs1FwcVuO8NFXQY4ohNibCJUixMbKSK67zVhhE1yWpR4IVSxCeX
iPXzFN9JT+jlAqJcouAEHLEM5/y2ISOXR6BlJ8JSrgGmYx0w9GSVI3aJnwlN9j1W
YJBl2GTh0ZgJK4r+DcWWMqAZeDfXJGGaGwITEhFSuvFO2RPqw9MiksJNwDncyDe1
Csf0vHr+JT24i5rdnoQwiIZk6SkuO2fhPr6jA/23unl22HUIMfnqfhapNvU/z4t1
MIH+zNZLPx1edwE1S8TUPU0CoegD+XW95c4xJqtIXH2bgmUJkYXClK0X+D0W6CnQ
IaJJo8rYgcsvqiYl5BSvFb6TKevN8I4lEPmaJSm1V8k/jp5toSiFZ4BHJkttvdNh
RgD3cfdSNvWMGhE0pwYOLIXpffY2RvfCtHvqGPWDhtIzjZV5ta7XjiNorX+EvxwL
E2MRzHDuT/rfm2i+zYZS/Zi9FrNN3SQhq8WQYGJNdS3lSGHUYBDgogTsSOgiWEBx
PUonxi1xBypoPNHELsscbUQssupFu/1vMV7rR/HDh01VT1pIVvrTbzVG7GlKafiS
6gunvVTAmH9fCu2CjFWBnfIPEjSwAvgWy4lk6FHg98+OMwgDaU+9LLfe7HedDMd0
gzR5oLjV7cmQ2Nk8iEc/AqHrethSAsBXeyS6G0PIWOqASO/NtAD2ZxlQ1x+JyAn9
1Tk6FQHom+RWBjr1z2X+MuIUphKLq0vi6ijVjg9HK6hX/l5G0Z730QGumIFUWOv1
9e6PwDHqZcC7QILAyoFgK2IdWoWeP58vso1RVOes15RRXG+HaP66vEf7QWc8dkOw
rWKyDzNndoBFTQALeKUHN44N/zYoVYaE8DVbXp3lKCXMUeeVYPblGWmVmiddps/u
uUIMDoFly9ifqbg9dxsx2wBF4iphAxyRZUKA0lwaQv08KzeFJIjQjDkiJPmM1iOI
P1CMjWdbmDmTu9CdRCF9Ugpp9aTVhfzNFb9p1lSjiQ3xBTp2dQhIDvPfSnW1k151
EgpJJsuY7ERhsbcnQzQUrjP0xSjMSiofxPnD7MmekaQmOp0NSQzDI+qKpb1JcpDY
+iM9NRvhj8zOVO+um00CSwC2lNsBfWIqp9XGxt01TjUcdg4T+rdH5jl3fTHS1cl2
JkWH/F010LpK4ox69rIYrd9eBf6Etw0/rLJjlzMz1CBOLlcNNcNihJHEH7oNKnqR
5nlB7TRLYMjDxkW4bv//tt8MMkgIPJ1hIiWCSE3wLfRxf9JA0CQ1mTNWTbjmuKRO
xny9pCy+TBCZQ4rg+Hd3hBtkxhSNvW6bp/OOJRPaWKJnfAUTk14w8bC9NZebDhhJ
N0rVtpZROcgwdcU6na9DVrhJ2TH9ltebX3qHvWD9xQ3xGoQoRGLtgiUHHfhVQySS
+2quKyCBMvfMhOahUtkB/Vw6DTQZRcv3MqkF0wF8vcK/2avvU0fUfROpI0eu8/5f
cYXKAajc3/h5hZ8/sO3Yy30iZ2zcJlBYsUocIO+YXReiWLqgsiSGzfcSE8b5cAhi
nWVydURJXUOs6s5MC/svdtzz7euVzUvRX3nXkZkMCV1koPBbiflpe77/8yPKFB4S
eepjEeY99b8PLHM6Rkh7DNmOFb2wytEXJZqo2rADnODmQtJtQz+fOKkesGRjJREp
uW5YV01G7aQ33yyOmwzshK2819OFjsAQPIA/0E20VCXhf5bVnelw+rxTSwQCOGMQ
KD5rTjQQkRwbuVibYZ7VOlH2Zl0b4yaO2Ji8vnUTi/GMc0XDIrwiZ4+9wBVys/+4
CkZT6xnierhMMFzgRMWamK7tYNqJdF/te6dmeLLAD5YRCU4DGwxrXQvN9NSnC8bh
JHP4cq5gf2OOAvJWCTo3OlBuXf95ICE/jjugnlcur0z5NsmyasxKGoE23TrEqb7w
AAYNf8tdHFwfcRRgZS11RkzyrEYR4LK06aOWd7Vql8e8ho/DT5rISfS051QIzFyn
OjjtUpUGQSTiG67/A4Lmlix21/0tu4PiU2Hgqqvd8VwsNTG1S66xlA+HU493QVgE
9QeM1zPAAJTBnpxHnt+5KAQYbb30VffHNPDOBGgpMT/T+FF1Bb1d25vSuPSeqP00
9plSugiiuRCHvuW3GDQRiQkqtm9w0QNYPrjSq/s7pkjyWhSt0oZ6kMb8OaVOtykI
QLWP+8Qvpjtz+d3pc1G1tXiji+PWel+sz+6kBToGhHHkuTGUpMXSe9ocPrkX+bHL
qo3a4QMkXxJROAlYs6rSsRuIecurRgHT8yKpCmwNCIQNrSqEKx62PGe8/EXZS5Q0
eBroBdB65qUrc8qcEKFX6TZy9tGE2irSeQVY4xUQw84FE6EEJ/AvgyETNT8ITOd+
y/2n4n2z7r4VjluYTLkcKPmUxrWXT9XjfRZIIPnSkyxU/u//9nPzj76JuAyC+THu
VHoIWrLGCgaXq6CM4XXVi8J53IYRNu+0dvYHXNIYOYTeNd1osVF3s9grIhqiHWoy
TVdklsHiTvSM3XIVvAWiACdwYmxtyHy4mnY1+MCb8GcgCsfmfFYAHLRHinznHbsm
0r0dyN8mnK/BZPx9eHhP5sYe476ejoun1kYutv3+OH8Oo7nM0+8m4XOcXL0mzUtH
4wxjj1Tj3fWlM7GKhPxnN6sYO4bie/l/oIiNJknzfC8gb6q8UOrz+vldHzULi/m7
l4VAyTNmHQmXck2WPTG1bPtYPdANsqfQ6g3uhe2ODBDhYLoL+ekKeApH2Rr2O94o
shnEcl9QCZlaFuwN82jqnWbbHwZErKsfckHNavLBqQUg4/lTBAz3p85tpE7XFKwa
XFSZEzfxSGSKev9kBeEdv+b2j3TvFPsJqCUQaikoYF6hK/F3l7mxElEEQeeGjsgl
yNFeIVyvS1r8qFNZZWUe4HKqbhq7Wj5Fu5kko2jMW8olk0/Qon1aioJwl1pq1jWw
11xkNiQiMAyBUqTkU8Va0eeqY1RluLCP2RdeVR40em5iarRA9Z6Ta9GcVyW5K0MH
o/qwTf8ajTXPFXcPig++g2FRJGZNlzGawYKOHcS2W2P8Da8vcb5Jwe8CIpRvWgli
M3TRqoXkdv5jndxfZONGZ970Z/LbG06oyqx385kG2qqRzZSOxLKCUrHPHEzEzB5v
7njWoA6F8SdaZQ7JJHF3i6NX7H2x0+ftfWHsqaP9ot4n9Hd0KqZfWqOfxWyXMHcc
UG0PmkC6m7O19Ou+MWMKBhGJdisN9PlYX12q8kmDMLh/HMS34Wwh9qdDpM0f7M0b
/KxwHQyDkTZhymlXZwTUSQ5e7AwugwXbuothCmUXhb9Y+mRKVTzTpIahaIZgfP4n
W66zS5ER5stg56ZVtT0tx4nukiaqy3V8Avc7pDENJqfacsfazOB+RmBtBXtAua2y
g3nLRHQCZIyvyuhXZJZ70iMkcPydQBVv2ywp6Iy4VzilIcuc8A/fAiRPYrQH64Ia
0CD47Aitegn+vaHczUwTob12CRuZI7yGaeW3zukv1ro92kZiSkAKlS1bWqf6dB3o
X1PyUAKh6/Gts5Bzjk4rzynDZc7o9ar8R2rFKt/ywgLfeUlwo52kf/44Moiz6XCY
Qvv8DLG5HSUVLSuP9sJl0fLdpRMf++IzNGQfXutmzNxv1AaHXzuf3IxaZf2/76oC
NqZCgdhMME5eF5H9c2k+FjbVa+qnJZk1xOI4d6SStuvN7qt//f4bRJ+iaiB0ENbm
WOqKNjI2sbYv+Zc8u9po/bMDaPkAzXlt+iDJnRZHrUBXlF6+i+s5BCTqO1kMLiWV
WbYMrc8uQF1dLS7neMmDdocFNZ/7fqmTyDPqJDYore9C78TQkPWqhHbtrTkYuPU4
q9cpsibGWHSzw3alu3X7xqLJBPNcxgPgVSLV7ePikM/Iwwp3Pu/Nr1GhCCdXl8am
ct15ma2OBT7xllwT6oNeUvyJNDuAhpDdIywCGz6/A9JOFXBXs52daJRJiJr58qA0
CcZLHkwQXZYNxRQo/Qu/Iss6Ytwj/Bs4CUSePkTAaAtdy3wgUHKirmId13wi8+xb
0EPvJl+855DNZVKpreea4MciyEwFIubrbKGlO44xDMfLpRcj4ri2q/qZ1w/8JZbj
19nIXs2FXVIp4FUv0PzSmHz9FzZM2MkcdSMwCFcaxX9mZAtDyJT4GR/paxPaCpQg
2uP6N+fxdbnuBKqnggFV3jJ7DEOPrz/XutrVRDoi3xTmdeBU4b/TvgweNMH+tq/r
emexxCQJAAj9R9Qx+fd+oPL/i56bZwKY9RtxHBJHzgnHO+3xjwRyZ2uSyh65wdlk
IUbW5tiMqagt5SWDI+qXRfhlfQNN09aBUw7lehMH/8kavsf2GHnQIq3/FvzN7QvV
ADpowQ3pbGoPEUEKpxGQUv6qAIR0NhGG9/DM0EDFpDu85bJRE4EF9pNZvnE/a8lu
BhYyIc+fe/fsRbWYu4mrTj4+M7dv87LJpSJ06VQ8mhkuNLc3qlq8IcbiAu4hsmnH
7hjysq9+xANFK4CpEvtlBh8CRoGvNvmRouTMOBdep1yclSDzINzaR12Ey+WAEp4H
gn0nz7IWap3oretUpnbpV3oKq8aruTaJ/2GCcNe+vYxdxBVxZmsltqaoz+xSj1kB
Ri1GnDGstjGrOlY4+nwGvATAtIZQYq1x4clIU9dgyID3wlL+ZRVjQD7TgXJDraJF
T8dGhuotlKAlXDM6HhLaAJ50os0x9V4Mu6PX32xA6DoQGCTETui/zeBQEWAgCsma
lkrIie4jvwodKAB/JS/auizwCqxhrF1GQADGZ21aoL0FDmkMCbMHFrnYeCNxDKvK
JwAnNWwsyhiuGTesIwamjd1y877CSjdUL924QJHxX9+AlvJkX6kKEnCfWDTEvgQ0
7ie7x+/fZCSrOcYmRX5dBn3xPgC9s0fQbj33cdVieR3xOzmkQfipZanlLR5VhwZ0
l3dI/aZO8RzLkOr1Q/LKTuL7mXJdWrTt/QM/xskgBH675O4DY66QzLytE3h0DQLm
L+aKw2Lr0ETPB96xAde2ljUjP8S2FvsSu475nPCEdu/XXMJ5UTNZhvToc4N5PPt8
xOZf2EAtbCDZe9O5tyTM36ifdvP8gLxmqokSKImtEWMYLgXNrPBFx2x9N9OwuxwQ
2kHpnT56at1OaWZXYmbrmzXJ3v35xL/zH5Bu5bkupPp/8NMCyGIDxU1+jEgE0G4/
Rt2vp342m7BwNpmLDUwGH/rARTIbKz7+LwKl8Q5i1MbKp/gHUkvZ7BLyEyBTRms6
E/9mAi8nuJPX78/r+pL4fpHGzEoaqCZbLBt97VLE5NwV3OITt/MLewshsefEbGWg
c/fKHseOdPcI0DFrVkVg/6ygjiRHld34GvU+m64i6SeO807stTvyaLdD1h40sag+
a3dmlj6yfrZWppB7BtI+pQqASP+Uau6HWMvCFqgk7p52wDeFJhRBT5/gSVpY2aI+
2mf23JfJELTsfM3IQu5z+mMS79c3mDpGWnbo3tOQKPtn6DKPu2YVLKz3S3l6AVlV
pHUcBdAWssQ0/AKvBhkoREomLYB1az02FNWBy9qrppcnLJvpfvQvO7nKM2EEv8NY
gHl3GkTOJuUVtUH6HWDIbLaraWm127boxFxN3nEIiE3TKWmicb2Ff97RoIO9Otf5
eR27tvCwoMvmsN9q74Awn5H1UjqgVsAIBjZA6V6hm6Lp+qTOp1ef2sSM/s16JNOb
kgx1i600Y+4VQPSEmAJb6rxq6MKYVP7SiTBa2/dldUxg7BpjT4HLfQY2qAxA4DeS
IcHs7t3axUeQ8pvglKN6xzgFmfkj86Q3qBEh39KTRKIeAN9wL2DMNYT3kqs5FalJ
oumio4JyTWsLL5coLpfyvAX5Y2CsBRzVQOT8azzc78Snp1VXhk1GSTKOLMJXHNpQ
K2rcRBy8QI51LR/lyW93A8K3TMAA3/sPJihwrAXrRDYjLNa2Amfx3Eu37bTLtb9M
TAQkGAgOL2K57oPzp9d7lN2ffIHthUJWxBsCcueHO0NdXsv05zCoIZ4T82KU1H3s
7n9KDx9fplk/aZQWFKOhxkte67eu4U4b7kUkzZuVenq6x5+n4uef2aJOclYY5p/Z
oPBBBNQAaezBtl80WxtvA/eZxV7BTrz6khkoX0awjKosaKttJkVJW7W58OOnCCR3
K7uA3A1SsFtcLr9tqYPE+5S6K4a1h3XefxhRJY74Lac5gGjce6kbWLeTmZ/+pZ9g
9UBuxGwYOb79aJwaYfNihl/PIKR+RX05dqp6C6zkT3JHjY0aWm/afqQIDd4/Oaie
+3wk98IcqenReYcPxdYGW5409RQpBmLV2T0UwBzf00ca/iB+vBLGpjX8WPASACyl
4XEVXDAJuhbboHEaHel2z4pDWcZw+CnCMlFqkBilHllTJQOW3QJQ4RdANSLcbXG1
V0gR5LiMmTrjA/4TYtgVL05taQ9JUUK9JKnroh+xIb9/+NT3pKG54E3c0V+GnCpX
SwC4DrAkon73B9KLjOZX6ccd20uTU107uR5ew8IRrIn6w28vy4M/8LGQNe67SvUl
MaI/Oa0QbYJT8JvFA9MfiKIJay1BlcyhVVJ3NXjr22truVPfFw/JMnjAnSL/SJLy
0RFNE3KPfeSXv/qfi+4s6j1FoZRCZoq0X8hnO+3soNT9rn8DGtbyU15NjTz5/v6V
6BfELgTjKGNveaptBvDk8DOSilkEu9q+YgnIqfCuPvooZsphgcqCBRz6OfygjeKw
RVSAPn/6cVExdCSe+bN9Jx+n2z2S9cIzX3dooFRa9Pj1pc6P4Y0jRsMuhVPJOMbK
2S+CiyNJO7sBNKO/gxMrk1HLwadQV9SdTZq8tqyGPU0BECshfcewggvJ6pZ6b94N
BlSD8QKuD/DpVq9jwANuoFWirVJsjO9GDHftqcA+UEnL7V7iH4HZ1V6qTKd9lP35
QOW0nRU35in2+WzJJ/xPx0Wjf8gQrtTI8FeqSuFBzfXWjfQk0W6z2mQA3Ax+g0sK
SaBxRzKumxUtV/T3Fod1Vv46TZWOVI/ENuqQ/eeL0oMYPazj0JnE4QEn5hWwB6yT
bsNFzb9GjPzYxUkdn4gfWXvff7gUQNWbS4LLOwMkq/9fpkMtdfAMG8QVlNvVoDy5
U1E76o4wam9p3xGL6QZDsxPNLbouKH/kFgmPSi8xFLHUP0oQekQ4nPTIF8rVrAts
U19A32PWHQ8QMNMu3oNPICxGFQaY1NhbR5vop17GQ9e70wA7NAX6RrvP3JCVUTk1
B/j2Fjhls1EfoU49/6wt120lTtjTNdG9OGPcAJUvCHD/0zr0Kkqosv6nRM4miMId
sER/XFC/nOrVxFah8EKoJMNncnOKua6xQXWjCxPr1ub3M8lluM2ULAel0FnRnfrz
U16IOx4gpoquH1Aq2VvE7irrMO1YMEHDMPI+t4CafiwbH1NbrSa0QhiVHln3GDWI
r2DesxMvqY5jtE233Y5it4eq19QfyHf1gHTdQDHllgrGJFSknsP8dIJHttMvY1/f
fKFGntZ8NHMDD7aCiP2cQ8odHuCszFP8MfdSL1/1qOWkTypZVw+9hsOBVCbUSlvf
mP8UfTnCB1dqTZXSN4FNCChTcRMSlID9FJPw2NdhwaPzsg8UWBGblXMgI8tWj1bl
G6nveFSR6TpETkwA9cjKrVDlFh43FUPOonvn1yx2ST5f0pt+A0SHLl9PD+iCaEha
+4od5T8/ZxItI8PYc90285oZx3VFmvHjfpE7FdTs0MWg5MnY/yajsQ/fiwC6lUp8
cpZ5V1njKhUZK6QZ9WmJjV96lZ3ZK7X0gIOcWzZkoL/XduYZMvELUZLi3utlsHaU
dV9FXWOcCmgm8UqB1Rmy969K0xdVOw4FVL8PUAKpG0lQwRqPLXGn5uuULD8YXe4t
Ioxd4IA4uEptO9SMduZuLob5SHgcpQP0ZUnMkNSkBSlVKQjQ24hJUU+IkUK/E1bU
Bea7vZ7iz05oPQghg5UppYyw/6WuYbOHKlyujU+kBAjQZr2fn29BGux2J+F0FxYd
iVhZhc1pAIHL8+vXc07hd/UFaT1izCOLVy0aeiedOs3StQPQl5WoDWbzUcuQHCMt
5F/HFtPtcgCe4tR9suctoTD/0kdgVFCYvIdLNwQtl/dUHO+o+DbQ46S4T4HpV2ho
Yiv2ZHoZ0iPKEtNCxDQYZdxAptFXyewpRK7Hpg9qUIM/BIb94O7qNfiFOae91Xt2
zm84qaeAShd4WnDg+bYDF7ipb0XPtFJa23pc6NW+LcL7I/vysKcNOmoijiids8Vk
ayrVC/P4BKa96vdEVtVJVFYAJf4eLNrubECjXG2VA4p0ew9DXXxD2UlkvNIb+0MP
URCMRSQSButgTneKqftTAGbvup07dmR99jLVCthSDXi2Pu/WFj3JQQjWY7NcJicl
lET5tSrXP1ahxgPZXLvGvv7ylq10Nf8lW3NIICdGJl7+ZDVSp0AtAhWBnkYQsheG
uAeFkSW6pRSFj3V/kuc1jfyXYFUYkxwWgwIATmHnP5F+7Q05Lce6hgBhDtwgY3WO
EKKrjUSpq/u2Bt3SS3zWzFm4iiy0rDCFmMeMVbzalWW6ZvwPHc4Uc1WYQuC2I3G/
wWt4s6WnfupL4knG5rxlwd6YY/ow0zsGdBAttDt2YdvpdrIhNOKsA7ypnJqY5ON/
ImiR4PrZPmEcdyHjSLX1ZaO77LUsssC8x0UlfvBex1dTI/kxkXizvVN/PVp4TShg
aX/mYgM6z4mK5lY96gxcT8iUD1jBUR4CPiDjFAf6R2xThCx4PA/BqpM2BpQMcJIe
Dl24k/N/TTzg3vbkRMEJkewRxKL/nLwu8aVjs7G1hAUAnkNoaZ1CHiliL5MhrzdN
Eik9IQZn2bBxdMxIs8LJCd1MuZ0d2ujmeN7tBTPNPSmFWszEayP8ABS/CDDWZF4V
MyKSe2K2hRXxbXwSK0UznSUzHpaYXtsIUrNhMOy0ezhttimVk/p2/u0Jf1ux0dnr
T7aIDZDmGfBkULOIHtIpl7UUiVWURqDQBP+g4I255lgKgSQFwTPZ4P+t5aUhcplG
WD9gGN1BUUzCjv0CZSMFaRwNASVEbDtj2RUEHvbTShaCaHPuCAq0xUCNWWV/XnOo
F3m5IRY2Hfl4quebgPmwVEfY18jldqR519eu+Np9Yvv0GM1wSrreRPDemu/n7OQV
c415z1zOrdBfY+4ve4MoQb+5NSYIoydZvOXJIVPsgHkjbNU2a52GPHomDn0aygRx
BYLT0kgwHnfnd9P9fJmcIcwp0p9gfdNnryGRMAJ/c84DSkhIsbX8qFYyYgtn4SJa
nE/d3dScVWZLkHjf7mjEet2yko82p9I3LRbwyaCBqQKWMFYULYYE6PZZJNcNYeIi
z0/ZuheN5l6ZDXF78ygDgh269usXHApUhVyQoAhrVzKFVfp4u583/fnhh10lk7WV
ElHhU/ZOQjv1WSzCXsTtaqHX7lccohOGWoxPHGkwN8O92inw0CYg5jLM/6SLSRn8
ZjPM4CVYZM00UcwwqSQWu3NQMyx5svmcq5WeVU96KS+YVGKAacpVZ4ZF8L13FIV7
gxPCULdVh+mB1ZficeavTKYsoYX/9Pa2gjA28LFukWLy47EuUbjKFVnk5+Sa2hCo
X7xUpCH/gn5zWtbO9zu2P7iQsJiGDE1WSG1cudDPiDoq5lMmB6TiIcsjycrDCtUZ
8ZvtdPifEnxjOntmgCuGvYiIIlm/5PEbum3e3TEKMY0qn1wt/AqEs6YVlYpSoo3J
/CL4hT8XZ7qlIz+kzqIssPvybhvD+lzxZgkSVhZanHm0eq8avlqwtBjc47eiDJqg
yARcDjMdWzhyBODNKf1J6Beb9+UXZ0FKca6CmWitcjDq0R0U7q1JGqlrdzIOmdQS
wHEcT9GulJ6+5eCWzTi5H79futQtkguQ4ZZyDkhDWXpQoNBo2xSj62+3gfn1u2dT
5EACjOmzEUXTHsi7qXLqSoP1dM/ukxys4J6XnPiHf7Vq65aHuhzdSjaZ21nd9LL9
p9qLDkN5PyFtgSq+rMtqP3+1H9XFOOIEkRnQjssOQEXxW8ZUEQicuo8Ngk3AwuSf
1JstfZZPMIHrCyiFqXwW7Ed4zZ4WlTOQROLfZmsOzY/Ak2UjtHh3qYev8ywQkR8+
pzU0JhPe0RzSpe0UyBK/y9A593BPyzGAGRfXEiq5zruVjxXGzO+EYHSuoFIWkBau
z2/vzVNzfRFa5pHffyIyjOEKvZ3YcV5oHK18A4kz92FZS/RgKj5A9nucVvr8aG6d
SB0YVtTnChQXj5kXujSoPymKgL1mB7hTgqT069zOm6ZOgbeDtWMwll/9kLSk+x7m
QPxtDAW8RN27AzKmLRUDqIPYNj3203dVrOAO/v5fWq0oHIZi8yzYzauWZOo+rEQ/
D18eWidn9swWTcHGZ99SLZsULboo/+zMpU7m8BboxyTah5uJ28P6Jlj9dgDgVfYL
8VEOfYdFV5keeNdTzlh/jA1WRZqP/fCNNmrTRuDpFcgbI+Od0n+HYTDFjIDWZsK0
IJiroPZVsjm9taYIaXzd+I4LmuRCxFdo0w61nK8Ba38C6vCIWnre/izsHNrIFRFd
1dFElrdBIONFiWls2CsQ6M8mQN6HsUM2LXKV9/OXzRchZht8dAqFBaqipQ2XcNMR
xe8w9oaVonP6ZDatLxMxnqIYnf/BdFLVf6YoRq7zVHj3Keb2QC7DD9c3DMyc909e
ONy4m7acdruoB/jHbwUDKBc0HfGXzzcsFIEdINTu8oOwJetmmk9g3+EHgrhH1Y+2
BNgLfe2fiqn+4ThRFyPqsrNbLUSVzk8dRY4QKVYFRdNVVDCffH234k59TOvZ0TwH
A1oqMcZSmDPJtyAdcz9Qj8RH9E5kGvRJsqGsSgAidg5W0FtR6d9E+slJ/lF9pyzO
kEhJ4Ud5HYKfHU3/9JaOmdEkVKG2Q0xxtI+fC+e2PXA9An40pcyhylSjMgk+/irv
PCvK3S6cE8ioM+7BNW9YL+E1WkWKb6Cy0s0debnydrB73hKtXdvh5C7ZOLiSL/th
E39Qv7Y6yhg5Vd5XK5GBxMQFjizDYZbp6VAQA49EOn9ZQicxRXTu7joScdTXGM/P
ZnWdkEGdG3KV4USLjwJMsdJNIyosA0mvtWImApD35LptYv9jtAc9W2AbTK+VNNKP
Jsy8oso42oYRJDavH5dYTmEzUW42ZDC2FTbJW0mQqIiF5FgKW7NQhPK9+4qOl1j0
x8FEziEzEPwFfgcvkgIoLPitZBWXMPsm2K8xEqlJXXFl7noXE6zbt9kfIWx/24bX
gfObSaF5uUOIiuoVyqCUS2V25y5vsnPt8L8P1ktbUgm57aNGfdFEuBmEF3fVoMVI
hXApjRHgVLdWD0Q6aCPY7g61LAlRzgg3B7RQRlERtB/xwahRFtGK5cF1iW6ynIr3
QmMAJD/RVmgr45S38g5tFTiUS2OoA5N4WBDmgWgzoOlyhqzYZlLwEeFqOxeovHje
NOfQwOoxhsaI4hbBGkfZVnMTcgkjK7+xaHaDPeep1MUbu84oPFL7HQ45SZGq9JEr
9CgcEzkpGTEz8zzBKKWV/OU3XQ0k/9tAfpsqWVJKpp71CBqlY4eOyrNSBpxGSrx6
wAw3HUiNy/qFzfwsA+8+m9pCWhnhG6n221hjxnwv5iOtob83XIjMMSOGs6SDDF8O
YnT+hTqd3cXmmvzM351/KAg8f1iLTc7rZZV9lW+wEQKi4QbJTSlI04I0+VJ4kiZX
5daKFfHow+g+wRa3th4+dWtxBgmRwe+qbCy4rY7JaHSSlJxXeMGVB2G2VzQMr6yO
QaiI3UBkDFRpWwj7q4LDw+TAcXbZzPy8soeBPGt2IaekmPRobqdjJFYmPgFFFfkr
07fzSmDRAJiqAmNEqeTnA/Qp4mMbSjfdWxZowZRoGaETviUEo+nQ3V3L0eI9XAoS
z0M2x6AAA+Rpey8LNZl+pLnt8PLJsFB1s3WZCMRGYmqbLDVR6Kvkej8pNuMvjl6D
RpMd2IVVKip5lwFx6fpIylR01DCy+lqr/8M/8NvLeB+z/uYRf/IUvEEWZJTlyBcM
xbqEjfwIuDlTgTcKctibB3b9jVNX2YO1mlCpCnhM5nuTntRy+6fmZ8x0FwcrjwTi
8efuGxE19+dlW8Alk8le41sIhKffDGw7ymxP4mYZxng9TsME03AuPt/0Pnmt/uRw
OGxpUA+Fx5DYfTSBKY+WRsl+8LoosNl7LlDUx0crqZXLgU5hq4Yvel9wS/UDV2dL
17pBHPNSuxeAEF6yRkhykDctlUuxmWfItt+SodSMaAAVYkVeePWtwDhd2oJUNma6
JGxruL1D2HaYJxrQ23xqrRZ8veqcwp3NOEJr8twIKqhL2zP7pikV7+1UMn5CAJWE
YmBQwTc7QlXjtHVxjejaq63eUtPJkKRCofA+c3Ucwfjlnh4UtL7c1FCwNczYS3QY
M/cxsXVp7i4v2eQZruq4bbq/rNxUS2ezyJenBhyxZksjNqGYGjFHkw3Fpl/a0PGm
Qf4NsnA/0grQbNaJFk2MYGoHw/ptixrCHooHmCKDh8ikztyLecVgLfgwvwKmNjXH
DMMUMeDSke5gJVRvvt0vUA3+8cz1R3HFD17uIOsyFYk4rkwaahTtkK1iQ/JAI9pQ
Vc74cQQ7Ij+PC6ncWMww9yCQQUWzsys5jiLvSOMPZitggHFM/BVHIPXUGRaqCmxq
7L/rXh2bsVB1SY7lJnP/shtefVXuOYkmUdhj2k2O9IR7K+A4l7CRQCN6cDg4xVDA
V/VPcaL+kH0YlMEZNCh6i6iCtT4xV33Tk+GscPJWhMb2kVNqM9ny3jcjrl1TYaGg
5gjvcw/o79B6cuFxQ9OF1ETW9FZ4kOakDZ7TnwtyOT9MVfKeVsFfsVZ1HkbIpmxo
bk0/AvVhzOrHYVZo2u2a9UXZLH+8HYnZ8WALoTLj/gcpTEkTbkFQofQH2Qdn0sVy
Z2kfWkAeT1ZV8g9PoXB2tBdtjS1/jzrYrL6PaW7O5I0OoeCb5eYGDWxxVW4E3p5d
lXMzvbmWtX+1vtSdGReIks4gnCROnRyGjHYwYHXX9CKgxXAkIbhcVczAGSxSsGnc
dN8eaRTetGNlN5HFdZCF69sXLL+M5c3mK6nC/BTcUTZ+PN6rkyZB/A53mR0YVuBP
CP+CEhWdtNHY2Y0r1trS1dm2RFIaojCfZ2IbuCpJRkouGVC97kGfCMIYrx3RYE20
PbWFtdXLgSptiIOWtHEJBIGi/JMLNOuzT8Ij5kXrR+pKX5dxta8hNI0nhGQQJcgW
E7PCxCRIxH5F+gr6lSViUYScNGCPPXs/dlgEz+/xE/upkuP5qwPPaaB6Gw0y3oDc
WpeeOnxJqMs7NjEkkYx41i7F9uqGe4Fw/tZJ8oYS5PHgdjat/pORNMVdb4fdlZVm
vLQNXu553Zdc0zEoUB3Dnk49t7JabuWYjRHLJoIJism4Yargs+xr+rBG6DtTcZy3
jTKTM77g3p691I7OxU4Lz/J9g39KQjoH7944M+kWTS3wXIM6BwitI7UJ6wNP672s
TjyhDDYAWSRLvKYAyfT2A5gt/KNVDE6agRyxiP8YGpls9C7rsZBa4qR2GJUsQF+B
/dFfrbpaYQRtyQrhG8S/vtNO4btGHLqdSEAksaClI4TkKc7p8fqRsWmVpCsx79QU
6I2epMtpnrQknRg8fQkMaqyFd4KYsbG8G1jTejzs2R8xbA4RhaaXh1iQgue6AyxV
kap1HwLXgWn3E39+j5zkLFXaPRcokeyGPAAFwVG8azXyrKM6v6YcYndfrxPKZTR5
DqyXxE587k4778Nz8opYtY66hhQ3H2PDBtDypdICaykuRmH+u3FTvn3Xp6Zi8iHK
8meRV6xKkQe8EupZsMrpYwaikkRLZ2bq9hNxCcpF9ts8YBctoDjZFevt7cF5wV3R
lhfKt2xDPkSfSviPCoVNzvITaDjc0rJqvw9MJutu7fjUv+FVfxD+PFy6MDgt2A9M
ulufabL7qCq2cNotcifF+v2bvaaRA907DqRg0aXdc/Txzm/45jILZDUuAvD4M2aV
yBQkmRWeywYzhBZn9iYTWmZQFlCbhzhKHNnIc+B8PLVkr65wMPg8vQBeG6qn2SUX
00u1kCRHF0EDaT37xeek6ItPuvyXJJYoqGDbCYJZ2AFV7zV1jvX0No8r8JSFDAoe
LzIRyCAv6AgB/veFvQc+TIErhcoX2H/N3jJZ3VOJV0sDmpOzZfFQg1vAVSoaQVSa
fvpqyIn1exaq5b1T1rDdWkZJMJFwgrBVAdJA9xbXdpBlIoPojktwx4rlLV9hAtW5
qzetz47O5RtgbbIY9pTMxB9NyyeAgPxnxrlOdWTKRxx3xzs6OXzqARlXX7Lrb61i
FLgsWrWzErd2y5dBvrtVDoJ60yV+25fPihuIjtQ6TW4RRvS3A7wvyRIRDDxWFUz6
VzXGxbAoz1sPoMgIjyyDjrre3W90dSZ6EEP85gDwmdRhtCov58m30LkkEnof6boS
tbhEEy4YLwHU/RFLGtr8Nd6v9OVijzTOCli9I24lg5FfZpPP53Z6QHYrvaUWVGgO
H+0tkLy15GdLmZzqmX3ELeiegTJBfrjWbgVnfJESKLjuah0g97U32IrL1OZ8bUyt
MPo+lu7IyiUPgcmdpgAZCzDgCaXeD+SXtvDc5c8mTgEoSArDSeuXIaJfIO0sx3uD
9lLCBDDmjx4cCZz1s66U8A51YhcyToij/UQd5+krqxRCRx+Y2xXXmSPkGjFwNOyb
qj5ZYuDXxc3YMQhHXq3cXjKQrmcVKv6BeYYNJY8A9+rqzdIg5KsfqzBmXaLOs7n1
qqZAuru+Ap+VFjngbsIJL9ZE+4rULgjc+5h0HxUdWFW47b5XY0eJeNj+rZ5OeUAu
g/wA227ys63LgvUtuXXj2EYXwadNLhkHrcUwRbiCH300lY/e+mM98BItO7eEaLp1
vxF0mSg8RWtf+t8EywAM+eUdy7pbRKjAQRMF4d54xQ6Ds0sBix3xkPrTJ1S5W8Nj
bcEuVLS/Z0zfQgN+m7iKT5MM2fiDF68tA0IiY3S7Ky+9/Y28qbPTuL6JRw1+qEA1
MoRPlgoVLye2wS/6bPqUrIFpXumHVOJDNtZNIep6p59Qk/++tkRghAnJlHeZOg9k
PnNECk+zK6sCPiUY3jRRzZGL5iLPGJm0uz8JtMPkrhZfg0H3Lh8c9YoPFxvyx4qq
LEwuo4H87XB2lOxGXe0l/bKlX2c364og3KDbCIOFFoU3N64BXfRHspcRMpwiR46i
300bqZbw6Abt2EgXRxUnafLHHdOgz7qsnH+8/Ky6QR3+ny9HDH5VJ+GMtsEt14rQ
2Z33dm+zZMyF+kwe5KRyjUidMnXUEyEKSuFsLd2k9q/6VNGp44VpbCC2oE7cugGz
7B3vBCQP54SiYZ1U8T1c9JiPyYc/EhSgopJXKEa+f2p4qXBfXUazbVT4G58zDtar
+ECQo0kxoGfRr310lEBqazizTdOVmklSVQMo7MkG6L/z3Y3Jq8eJkM34RTOjfhCF
BdElmXlnWVT8ZNp53Lc3+40XNFcaZsmcGm4VlUD+RARSbG6CweyfZvacnF6gvK/B
oOoytKVW4C1BrAMGF5/Wxr85C2fHE44CdmSzlepp8FdiKVgd7BIP6uHUWP6QzMI1
Yh6TA+8YNINCVw9huwvZQ0+7zE0n4pPPZTP8W+x/IU86fh6+MzvCVTsHeIV47Htp
gUsJhdZ+pAwfGKuz/uhJD4hek7WOtWKF//DFt/woAkbPwoE6WLVvA3g4qS+ULWKq
Z5U+Sx1OHk2++T1fpOZCqpmrJvotk2lf6gibWy8S8mDbQWj0dMTuFltt5LY3d7eC
xmGBlLkpx6jiJF9mpDF+LuUStW7CfvJ7QP6zbu0Z+WiXGjNLEG86Tx1sL3l4vLHA
fFmY1ZzVxoM+DkOMWpZ1ZCLeCu2nm5KdnM/slTDfrB9HdDtRKK/qkzK6ue7+z1/K
LMJ+4fj8EyroeMK7LTL6agPOYEw1ZIHhwNwkknmT2J1INcR1ZKZZN1+x/KMtjAuY
TQqp5fDfl6Pdy/YdnONNRjPKbWlH2UjYKaN21Et5Bwnrwv8YhMksSJab0S/zjPVN
/LcFV5qCJvPuFOv0m2WjSm4VF+30uQBUVfjWTMN9OUQFp0DIMYxAnAovGVo/4Z5O
VIv2HvcJdFQjkFuNqx3dmTBxInIOMj/CM57NQQ0RsPvS5KS62NiqPmTRKtTdMwMm
mEnpECNThTKPg8U4plQshZyky+mduC3lAjEzzHBBlrXvEyfdCHA3xXVSROVldTa5
Zmx5P8nu0pba5bkevxEGt9z9hhi3ZrYofMQJLIqEv+r1kFFN36SZDh9ekNS8OpgS
Md8Tlr3420RizKxUl5zAY0aUEYgLJu/1X1hNck2LzrPdTdgAsGUhuI5FAEcgt/5+
ruOscsUB7PuttdOi2gZoIpYIZwOTU2lDLqlzGHdQePhAIhtA0pjbWwjwlQUlfk6S
otyoMPvWsv/jZvZpC2CaRUZjCXBCvjxJpEk65er9aY35lGCobhgj+dUBBtgC+6KP
xosEhHW/EFelHS14vsbjXx1c9pkT4oN13WttNhMnbf3SpBslwAuhS5r3438jKLm2
9mb/1MEFyNNVF0w/ivYxZaFKgoDuEn2H1FvSS1XGuaf5lR2c5+M2kG6hmJ4mKKCy
B3vEIczjesxmKQNRL0wtiE5zFWFBADRaU2YL3rSRJhQ3oRRORuamrS8vtkbcAcV3
m79zVrCLIdFQPqK9TRmqbLpmj61C3YO8TZUE/VxppmAfR3fEGQp1p13usoBhnHiA
EcUbLtwqFtdzYrL03LBf+QWtIZr/Swu9epMYyyXD5z/lcEFy0hWQCMgRxNBsSSyg
UCxN4LLsHIYxDqbVZ5QwrLi96jjQ2sHgpds8Iodn/DLHGBOmi5RpQ98bTwOocxkE
kLfrmVFChpS8ryKllTU5EO8PJZwTDX5DDar5Da41dMZSNKJU71t3rT7s7hsdOvKH
LGpVNbWxsd+wOlPwhL7I1KzA2341bnxk9jsR+HtKAlMCKallYwuZZf0cBExrELc/
mBthjvmVZFML0jatXDeG3D+SgEUxHLZEVfKZfc4tZ3E9vT6LWn+UEaOtjZEpbVtZ
nvxDD9W83nrE1JhEZHqbTJ0jbiP9wT6eYrM183Y+te7QzpfMrrcsNi2hOffEYnpq
oBl7US3i96r8ukss8ZYQQiRVI55o3Q0ol86tOUZU3cSbySKieUVfV/7RjR3UnSct
sBfnJ0kvQeQb+otJ7h24SEUjY2xzy3BhNieP2NqmfH929JmESUp4cTBv+t2mZLIM
WPqjM1+9RKBCEfAJpn4Xq8dhf43KMWk3CB2MdyxuZc7LWl9p7eBjlFGdi6hOFpxR
WgG02+KdYSiwag+vgSVTAUvf5JkxAQqXduL3AGn1s5i0gaTm7yOazwYN+8/ofGRW
7PCQJ5ixGtMtIydSN8KZpa5q6duV/gAZ5EEft61XZQw5Im/ZJE1mXEmBGwQiRKVD
W4OHkCzwF50IuZrXbcT4hcwyN2ikrxwbniEhozH5EIuq687UsVHZ7Ccrr9O+vKh7
o2TXKd1srUxpf52Bu6sqgrRBUgOUShsV5tqLwZfIy6dnpnPQzJQNDY0/UStLXeuY
BHOBS38QMwvfCD8jbPDMsiilpRzj1BasRcthaANPUWVk0V5mcaxSUeUfgRe3Fenq
zgXS9FXwNBc06phXCWvPnSfoJtXxTnKg/xDutkeVLFHISQn/uB8sXOnV6wBlDRF2
OCvzCH38GP/BW96hgsX95HlqVRU4zcINoBWw52sY8vt8UEdo7pjk43Maud7oYKaP
jnb+No5RfZAxxfyVwx6ZEhz67tWrMaSvDi9nMQdI97WIPRKsFNJmJgNA7zzeLRBt
Dv7H6GIFkGxLmq9MFnxJ0RIyZyuVN4CPb4v6O++Kl90OuymMZVLHwmnTSjPVAczZ
shltCiPEulnCLIv8IXjpQrB+g8QzpGWSjYYZsene1eDDh5Mu9Hic98KKes51zSZ8
+I0JNilJ1vZGTRrPMAkHj6xrIwIMJPVmdwiP/xRq/GlUvJLiqDjoRC1ofQl9XsBQ
Bs4JuTQk0lRv6pL/2lZIwH5M8Zla9yhcFDgIRkMRotz0wzL0UY1zlKdPwtzQlk3r
csZAXOB+4PLJRnNDnhBWePOhVl4pQzLqxQy2mRgKXMBwxWbP9jGaaGvFQkj1wEAG
qlhiOoY8j1NC1qtdjrgCuErBUkS2Vxg8cA8ekDhzPhfmHX+zW0ReDr/QF3fPHEU2
a0iSCnt4PvNBx42P3xcFj2YcaChVSDyVW6pnhTDwZ9digX+o0rrzIelEbM89HiaM
LPC2dfblyOtyk1+m3RLOLFoN7O5csaNQw6jThLkQKsi2W4crYsZmBAqHMK9f1ngN
11PvqLKgkNvnRGtcIlFEaZYi28fDd2IWWELtCE9zI6t7u9oY29XIw4zO25vDpWaB
8WWfRv9Xznm++1PAmPBN6B9kjsxd9vobOYaL6qIG51YhV4RsBqbPnLwN2l3kvYNp
beKF+dBq0qyV5/ei6ZVJS+oL1FPNXf1CkoMSD4HAmx7AhGm4zPH+gL4vbius1tgD
E8/B6eA+4BeNC6aJIC0x2Z6TqqvvyZpFUeJxlnu6PQKDWsCAxa27ogACAvOZc4km
/BpnQAU3JZTOsVscLebdMvfa2eTAYDgkuifOt9aEWgSnYMEUbnllFXBCmM8IC1kE
U0K466K5eyVh9QJ3ygWbD410mjnR6myTj7/B/015GV+OSY4MOtcobAjrFVQcIfe0
DawW61XJfXsH+UUqTf8LhDv+WF5rvt25T+9CB5Dqna6jbuurYj38ydPHgI2e8bp7
p+P6yAfmnXlgoxH6KP5+IfkT15c9FQsY5KEtkdyWhjrRpWXT7SlLjKT7xKYWRW/h
vCA4LWl3FBZjgnH7rpmj67TfRj/dvWJHmayqEvVvB1a4wuH3C54m7Tf2k6BbR8Pq
W0Se9gKbEwdhLEX2fbrMtFSbLwX1E0ChpHlr0/y6QWwZDMtPB3QPDsIp5u+MD8dg
QXc3HK7kQX4lkLrXBVW1Jg+4/+rlg2kDLaGXVAtWIM4L4VSkpg9ekDtEOuptGt34
v35Ldpj8aX90E2dUvUn9UzTv65fFVsy48VRoyMc10JVpxFWGUBt2KOT269h6i15R
MTqr2AQPnoR6STYzqo09wEpiFbscmVT9ypKxhuZhe5b8q0f7nzCXh2Xq3YR8Nhye
lKqteHgUFI6ZrGLS9jbOp9SXYk5/NyplTrC0xOK72nBSKMt7+hfHyBerhwEcIs8N
Qgmn23gCIY7BMwWkQl5QF6awxQwkp5yiHnvOnKvTVgeHcK5hK8NfHm1kh7Z0PUXK
OA3L0qFaDJbd4ZycOtWwAsb+/6dalLtgx4S1gqS9DWxUG5O4Z4KQBp1fDiUtG7h8
kGNYaHkUcL9Ex7uqghhKX3hg2pI3t5b6p+JTXb3SZAyUkGK3fbRFoUY+/pjglK+E
YxGe350RwnrAki93SuaTjrRdcn1gjDFwezDYJx99O8Pv9qDc9vlw+UQ/fXEmiJXu
BdhUdc9wzJFseqbKlK7JlXHnntWnCE+0pOXzbTbWPYLIz7GtSwMEQc9p16fhJRkz
69+L9WEZ530UAZ/liINLXyY9B8Eh9eMWKDKIHiJmqjRR8OKb72fLILbt3q7orla2
m+EgVoTkCT8TH5yXNq7oSgqA0jiDeP4knv/JXOP38xRrYzWkHPXQRfpJbu1yxEcs
xZyDydGxmfsFT09nqLSDEcRbzL3fIkR5kyafAG2CRGUDQs3fOKUF4DMZzsNZbAO3
GrUKsRFdAJgkQKoSU0hMfiCduJSb20oxz3ZK4/4Fq03WJMt0PDFyDuu6oY/olv+X
z7Hytvr4H2VqmCmOet2z3g==
`protect end_protected