`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
dYVY1GBMsK1ODCn3ZUp8SoAWP8Fvt20jOclKciHf7Ysn2OlvHpNHbXI7BFbSBeZ8
c0HSNxtSIQSCmTTcVbiOe5bNYdnShY74EmVDlUagwaODhK9Urx30VHPfg7K0Q8Dj
u4EuL8LzGtWyNpPuuYUPfH/EWWJz8j2B3GlAugKl7fR1RciktYEXyNArDzj2i2Lo
icoQhkynNgC7v9DkMLR1BxAwtrFrckccZalCrbzlnjwD/DOLPtfjLaczesJPkKoa
xZJUnnMJHmZHdGCWDxS1eicDF7kXXzsE1BA2jAX7HQtg/mw+vmEQXKqvkKy9tRtW
yhUEHOXSIVFkC6gJ+buK9Q==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="SgR4h9hEc61j3UcDg7JP89NUc7gPf41F4aolx7zbZ/Y="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
PcTZf+e633x3tw5Pd+98Hvg8K8pEx1TP/UFyHup9OvIvZyp7VdJ/eQ7Czw0TCb/d
NGL0fQmqipTyP1VBR/CwCDPv8pUq9mWdoIhPzGBVMq1ZfAiLygNMWUwFu0/xPfyw
rAKvJfKF1tLDCsja4oREz1+w00FDmJ2gsQcbY/9d4Lw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="fB5pBzxyhRsqq3gFtq6qZ5Drx26WwP+GzJuJsgJq2oo="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 105952 )
`protect data_block
Pw0LuTSwA3gmWF21w7rVYBcj97hqvAcf4dxm1w8M8xOO9V5Zp53fD6281Uk66by2
V+2le3pjRQ4JkfVvu0vvltrqFdWvBln4SM9xPIyOvOjskVz8MBZo3CILQk+Kjz/X
fnbKbjecJcaTOqZL38FoHQEwjnf5cGCAog8jMuecu/61sEAHFkDSYGXsRGXaFaUJ
AP4+QfemzgqAzrzU0EhBXQnv22XScH+NLm1iSSWlo0ITmggpAAyCcESYfR9/XJav
x7i07KCTZa7fH4FzbYfe54ZtpODFZWpLdJcfAMjPpxTK8+70BFxTWVRpIOLVPTbc
yROzQiV0IX1JxZTgZTPKATcCo2yJTovZp5PBANq13EKcmlE3c61s8QYMo/EvIW6i
ZJ/AjqD2TldLSETZRe2qk3kgnW10nhvU1b9NPuopkINV6mNTrb6U1VDIyayfLPF/
Ep/40/oRj6vVroeTjhBhCILjeQg3caFUaUBrbpcskVFQC0bfNLJiy2lX3ZnlXK0t
2xYsKaUof+Gm00IIzB92INQBLVu9BUW0S0Qi1D7yc6XVerfxzA++eCIUSi0DP2ur
OdVQSbD/w51JTo7/u29i2VYES8zIVt+/0HgSgevj8NiP90ykRhcLqqkdQgFc5qnX
5UBkE82Xei7fSazmYQfqgVN6T2YXDpgH8OA/TTcFuLrRCvSIiq61urjmRBXHq3gZ
g5YFthowr2r6NtGAJGD3/jUDEpIstIs80pgsnUHWg6Wqh8BIt3Di025TPNehsOmn
ywbhu/fy2ueSuOFK4o0vBSVIv3voTnEgec8QlVJ1aAILzPa/86poeqLG4WuiOqkm
fqM11JRC60YyD+lhYGy1F2eiPq064Xogf5aeXziwg06a4BnKzdfSfW9SQhDsYk67
7hxO/OZGDyAu8PM2cO6OlVz1zJRJTEd0HsjavTdvRtCE69xeZMDyvWk7uaYXFQrS
GKXSQ0e8SzMk7UsDquy1RFp9iayJwthmp/PP+WOOr+Hi2y+ocXxym2II1rTFYkHt
4wAqt4s20b1IYQ71Uu8QFOZEJe1K9X663Fo6JlnCbe7HIahO4d0hZctdlUAi6Kv0
xCKuzzCo8itqSf1ibuFij8y7K5RK5EeNbm3PGVlQlPSHttuDUPwZIZCS+tK9cYDt
qvW1AAdJvBZZY5DZbqVOxJitqxtlxLyOnB3uIctKfw5/uuNxHyr1k7IWk5cFTUFF
2SJvwkyrZmwqX7XrGkuQJgkeo1DJ4Pn1evyu+67mvy4ctUgytq9Wu1ZAo4+cBY5u
CVOVXLItDTkhQcL8kBsBi/YBKwH648YGxmtjBXYxZXb1znztCuTqQ2z+hprAYZRM
1YZ33xXxIqsPM0hspQ3RjvWuRODyTuuf9v2u69w6+rmPYxgqBSPEVrDD778mLjic
VWSdzYxvtmuTgBD+vOhd2/tYlR6ngW54H9Xphu+iOYSNvX+XfWhAmjDr667f/LSz
Cs/9P9RlWSBkE6ZWp0FMYrl1x8U5wNhyMTcJi51+2lNB+SGv3vfPGFXvhQB3meuM
HPaAKhnqQhqK6KtPgErKSvJhwDY4C1ET5htrwXUDtUxoD+SAnyynbF+Mys+Db+3r
UrmcsMB/v4nUpE2Al2PQYtB/jTr7JcKw8D/j05349KNxvVgGp3pDrPgWBQgzC6RU
IGWTJuB0NFIedyU/j7zCXzSclNRJ+yAyQOhrlXPZqPIgBuni6Ryus8a4QIu+X/8q
cWYJck1dwAYSwKT9S1pFYUFn+HTqdIArXkI/ozpt9PnITkYbnO1RqGo6nxy5rZxd
3UGC8bfyzVx8tGFk0qYTrkW3gLpKjHh2G+7/N/tIUV8FG6wGcWCrDl/rzNfIO/iS
g9dU8N1ha7zTixtihStWN5mBdKaJ0aFf7WxI80bLq4u0WSORU2w2ZfSCwcnfiX8g
HVHyaCUUFGPT1AdAZmXB++2FonLQMubN7oGw3DrRkXe3iKSffTkTfD/6NIEn0r6V
oemH6wOkZOXCCpwP7fy323i4gqqJey4ZVhqPsyK+feRpakLU9bKP3pYK9o0lheva
WrBFbwa3DyDa6ttlaXrrZKqnaxkcBU4qOBVHarG6tWCNIPoXQ/ejQzQmDrFgeG6t
C1KU7jbXcCxJqIwRIBdQyndSNQMAy8zzt8NrJgTKgcjNeDdb6xX8k2FW8vGZO05l
wSGLAtTdha0H3qWwoIlEI7vc7MpsI8rFztmau5p0WQ1Veu6OuDm7SMFPNCrLEYq6
et7Lh/hNlPNJB6K0iFjU613wpB6CMzNqLSb88zrfue4jzRuppershCs/sNkv3awx
srxaGzrpbBAWZ4QuGfx3yIzY2aKa7Ku+vTtE6I+47u4JEguEKf3oqcf4W9QpwW7i
Gl4cI6otdctqn0n+KIXs49cSmIZs6ZRXU3IyaDNOrEJt2s27o/GXe2iMmCBjUDZI
Xvr7RcHe7dQ/7ojtnCjXiT74FuMh3Sukjhv4MxdmcyNpSWc5KgCyVP8XnwZKZH48
8rgFNHQDqbifs0JjTZj5fR1Gy3inkOi8pkrXD2taDNBqFzVAvpjkN9rPto6SNMgz
E0VXb+gaUn61geR2PS6THhRDtP2yDBanomx6+K7hOoBZAKYlFzO2uTjW8TTMqAsn
XhZRa88jGJGXUrOZ2+onyBmu0KxpfaG/jQ5aSjMe7Hm6G/C7w/4sp98yKBzYPsl9
GhS88AHpvyW2bm/LCRoM6d5bmIGTOvDPHR7xj3BTuCdo5auRu9AbgFGtQ9M8m7KC
6h9BiPjnrteIAJSf4n3+qC+AAy1Y20vd5xtp3CLnf0yvW009dxT2wuSCa3oz0iq5
P24tagWHVkgKl/Kw8PHEM34ELpyykCc3HlWmH9YI0mSC5gn4AxlgD9nHXJc4eUuB
dGX6BhVKt763Sg9jIp1H8QeW+YdeDdmq6uxU4MeTBmGnRgR5YEWY93uD9Ua6zA+V
Rjp+pzR5Evx0i0JedVcErUD+LJ2gkdPDdiJptWqK1mbhXLMdt+ZsX4DaVJPOjExT
0OUQAMTKh/l1KY2NLWQp8VDfcrvjwQDaxJ4tkKSnvzSrtSfY0DkF7IhaRgznVXVo
QtekkVExdvKUwR1wdHYzJFF0CMOXIIaK9GzATJ6qXtw8sUPrWtiTevGtJZpmacVT
iW3YVvEiUtfW7zuOwdfFtI/Zr5QmIUTa3+tMQHOo3MDh1vQzlRU5+3uVNKLBZSjE
QqzHkWxmnPyWWdu2cYPlIQIT74tTOpkwHNOWrbT3+utc0PFjclDr1IoZCfeswLqZ
wFjfYS4ss37BmuVktrca3QNXkZ7NdciPZ5N+I+0+0EzspT/rQX9PSXN6Rb6twJe8
sUbxNSyjofiz6FX6jHoXvwO9wFBd5ABZIa2XVil8SdmWnB50DhsrTQ+ov/gGlP8r
9EnloTqPDc1IyLNSReQtKOyo+nvADGmQ6OiSjwQ0Lh01sa0MxTw9SgEDUrzmSzf4
E88p0dlybXVGYQtSb4zA49uxhn94bqpfvUgeqg8wqwG6S9h/t9Qsh83TWj3i0FQI
FnOyaJCIvb5jfwYQ2I/84we2YCbYg5WoouCTD4TMwVsBMGWTzu/efpVmAuypTrIO
XJy48U1bOrXv7aIVlPo6GNlUELxwuqpNKLhEN5GVt2sHeCVoNMSL9vNOhvcQDZMe
QNzv8+QUpIBRLG+vkztEZ7KFyQ4b7bQVSXDwIStbSXd18hxYXDNMxgfw5qiLkeaJ
Qckd+aJayDKfjrAP1HEtweTM4uD7GPEGzQ5uCjZ/wOKShT8yID0ovHRQur3195H7
6fRqCZ9s+gj5F67eemocKrIULNl6zxlR71JSaSwsebkl/qcbA4t4FHhH9NdDh9cU
4EHuArTQnDhjHf4loIUr1UGxH6ltA9ZiGkTCyyAqL0YCSmIrhfmdea5/OD/GV8iX
DNgtbAuZ2bQx0nhSNGWLjQet3FVD0VRrnKhbU/UOOJwOgJI6AkaN63v83eRlqGOD
/bmhaOjMTRgSJgIFq/hkANePq/Gz94VZ97nI3BiH82w6I2HCX2bOWmJBfM1EX/aL
TS1zAzJ5pIuqbRZjaI9+pDD+hnYMGLeNl/gsZ/WR7giL3gXuR2hlNCn6jqiMAn7W
GxHH7HznwxVlyLPnAWa0Z/bN5w6DSqF00Q9fintGuJ7XlzR2DDy41cz2fHcl84I7
I7cJt7ax4nqYLKzEBVj68oT3EkK8ifHfqV6UU9Je+cPR3hpxVcc83KXggw1lJViQ
2GAUE2cBveQNhU3bC/3mq6RUkW5LEoofftA/SLuJ5QdT78OLFMYi/advIghxCOsW
pBBK5ygKDcj2lUC/yN/sYLrwB2JG/UkBQ3wsHa27rkP0F/J11mMYHFG6KBkJkC7B
vGjNaQNo7m573smzY7R4J8juJOr+MeS85qmyCkp4VGYo2xVUPDAB9r1RLxl4/ppe
Rcuw39Aa1Qxiqc9wE/aJHSHlSL2udGTAmTG/EKy+OrtEdwv/6ItNh75uhCyKYqVA
lGl6nafg2eBc5+dMjehhiEKM4vCeuCt3PJOhN9hbKEe+zjUrjMK/6LR0ZRszGOr+
mua1NjmTXfE7WI/SQNz2movRPvDmvyOb/RRoep21P9Dtp9qVAp/R9pIWk+DMKbtn
izww/VslESB/TQ5Pydwz5WrjMlPIuaP20T/HLfg9myqW3uIQpMjdoZfmwsID0KmH
voVi5Ns5GJjna5KJpJuEiirkHkRabZC4qwsJ1PWm+Ay49Xu6k8qXpCR3/wqxKbUm
WSXil1XTuxyuqStoh/Sr3xFbZl7pPc8zfLmEneu8vZ0I0XHorMXi1+w4u6VFEqhB
MBJEK4UstMIEb9ChV1/B6cXkxKs0Nt8/1agh169ZWI+VEqq/hXiY8X72XmPUWSeu
J1Memu/HSc8vuHi2wxJXNcPIY/sm4imLAzx8fOTNcgLQlidd8y7a697zwjPe4siu
pFUnr57rqcZxADE7pFJRWWGt+V3MwuHX/HUEelawAwHNbGmovm5KA8OceZmyEvCQ
4ZpwF7aGIeWV2IZJ/e/WtrfZ+FMOetmNoMfFAcW1Q/lh+jDG+NOnWH8TcO1MdLEg
iyhG7wTTp/BH7tH7dCXclniYxguBUWn4zG7a7lGJK41kk2lwdkrjg2+coC0v2SaP
/dydZAm94RzPurxXEfFZyhTzxXAIgvRpaeXwFhwrT3aWoxtdWE51hkLVwz7ttKJB
vfzP2e716Ll7nm5edPq6gJSZgzsyAfYTZAVpNj6gHsSMgE3AFpI7O6v2JY2Z5Vdh
xyr4kFcNGj/KmoIwHNoD+LcRVr/aiscXIaLQBI3xuZE91MhIREAHROWSwSam+erG
67r/zpAlTBcFIlRpVfHYtM2U668g7Onw751+GKQ+drHWHLUdPPXG8nnx9SvsVWIn
TevIp+Nc7+7azQbw+EHIn2q7lFuBqfm94e/182YHrDS9LzeoTIV1F7HCO331Z2gY
NEf1dtXbph/SpNrWf81IGR/6+Q8RVm4rFqpO/hfE6rKB7BNthRlskxbxRYEtpJ6M
KLBMZuDyKeoKAgLVYALRx8Lr4U9gT8wc7vMh1q1syIpshQKVB3AbtV3Z3SbVtxhn
w/NWxd7DBdmaBGecLAyHgq+rTnY3B1bp0kbmPSvGXOQ5E/WamTMP8Srdrv46o5lw
bf0ZKj+yM1MH74P9Nnu5Ppyq/jLvxPeLZ8gjL4XhpTbL8aouDudFmYsANn7Rawmo
xfkgZ+oXbYNWcSwJtO0CQ0rdAk23pS97pNfuMKIAVizkpN+txMlv6A+RkkxxdfJK
Xac/XGjbkp9vCMvyfHK08WsffGedM+m51SrfoLvJ8FNDOIOlw0wBt04UlXOoGC7M
5il33bzV7F5PW4cjSQtJepwJP48FiZbq4Mhmr5Hy9sGJjVzIVWra7mY6IW5m9q4m
uZRy8KSF8Altnn72VQa4DbHKQhOSNjWRbsxAO7E4YYNwfhPIu5FF6kKM75UH/kG3
qpsRAA4ZaikuzHzhdkOb09YssoxT986ea3liIXpTqWaes8yJviy1F1/9V1a47oKk
DLHd92kShmH3Yd0vNDCT3i4BFN2hZ+HCBDlDE04IRW6LrRM1v9W1RwSjHGv5PGqo
ZnxtbO5kCb0oPQXSWhhalBvQ1jaMRL3vWbMgD8ISvBA34y+AC35VKvjfjv/bLqCk
G+6fpg49fuY5EpDEp4VytE0N84vG7Dmt2h0Tk8Bb/JWwqhkbA8IxEeXsTd1okfjy
upqddXo8uOcb5xtHiNn5SIocCqg8e/78xDPbedJRbtaLFpaKCQgSKTeN/pZhWvIf
VAUoXHQYVJXPHxn9tQVildTrac8DUTmaworlMbh19i3skdz1KiftVkILlx1kpyqt
D8pmGF7CtPk5Udiole2F5GK9D/ZifPCkr6C/nuWUp36PyVOtvE2U52ELg36Qs97J
auXcGkxog+1iCcIFgFi/Tv1HHWOiakJj0G2Hq54GhhczvZwnxY4wT3bu9OaxDZXL
SSmhEkZ3H7lnm226prVEHqZezReTf1f2QR9RQZDJT1dCYRCMT5+U1B+/hcZhv6Fe
SJgqs0nfAfSJs3JVkn9bPEni0PvdQZ2SBAs1+V0ScXpb5QL8/vGhjkmcasMNK5yp
VIPg0Mq0R9TXBYy5qlXUc00i9cK9HFzyrEjlk5lOUCMC/Q5KsuLSS7JCixL1Ni/t
yevzsm2rvtBl/10j0lZ5MBicmHWp8uLe8BqZll/kNC1b4RvuUAoS5NteW/aTDXQz
1XyboptZs4bU9r5sIDXgbFHw4wdVqhNBHcEHtxDwBDvrTEqi3kg9Aa6zoFeGEREr
/KBGpkzhjOFDRj121o3u+xL2BhfteHFZZnP7hcWTjngFYNM9d7/kwt9xEuP0hWxB
gw08nljr0wkVTq75eYZziN/D2arqjSjJg+ieU+mwkkbmO9PlcHsUCepV3wzg/Frc
WMmj4JwQjIKJ6cy0iqEqfBhfgbsnXaRH6mv8u3LczM2uD8gWelkpDGKIuYxQRYkA
M9sRCIIHds75J/Hyb+lqTAYA01UIw+NqdwGCaMBS0Lscn0lnt42fLybQe4kuo8bZ
VBPJI/jQTGS5FzPE0F55Cjcw6D4qWz4F2X3BhyxjwzQVHNzl5Jgir0BTGGG5zSEk
DKiX5LLQ7VhE5CdkA8mXEqWOWutvynCZEJrhTsNjHMecbAHMHCIyyyLq1NCt8dl+
Bf9ZGFTjNrsLYhlCkouLA0eYzmAqaFw0Fd/vhlC6lZ14GRWh91/07FKT5Wx29zWG
31zMExIHmitjQBtZqaMHotj77XUwfIuMkPst9yQiR4Dt3Y4d9n/kwc6Fp5WU02cp
HqHIeSlivJQTGi1UO9dhW1mgOr85wck4VTReTb7rEiU0nwspVKeTrOWdgnjegNUd
9A1I4hl0IfQkv6wkrQM1FOKDPBOExGVGK1IQsk4nJ4vLZnG72hseT3FGrmrdBQv0
An2x7D02atgzLgRzekBd5hTd/VHnY/Zwh3dXDRN1j9/FQY7rOkup98yBKCl7OwvB
Ahyvb1f1kqbPKmr+XXJmjoPlQj03bl6Z5K99/bAYiniU+cZzXQ1caITee4A6QpG+
ciefSgQjr8oXOj8svDqUcveNwyWFW9yXU4mLIQGP1I3oZjfU2jST5HC/v2dIWy/x
WNtBzTZt3zL1kn7bCJB++TnfVoA3wkgKKbZLEbSHzutVb+Kx2kbIK3T+fjT+1WLR
XGzGbbhNuDiP9nnUonAqVdoj8r1kpTxLadORcNizEJabtazBdG9oKBE+qwgBFagb
sbthZNEjjF/F1zVNrgVvK8ZxJW2ZTljxhHtNn1Zu5dkV0XpqFEeuEAFBmaDBx5YB
/9G87XM/dwR4BHIIqc+FJitVGqjwF4ULT5DSDxkv0oy7QMW+2opi8RpDdXbOitiI
s2J5FnhltkVKKderD+MBS5ZqFbK+llH6bzRnYjTqD222BnoI9OQ7BqbrZRI2xSMp
cr9aic68Re7KouO0fnhJAA0kFiwn7u4mKg7D9/PjyZvFXb58LXqBlhPKdiurLR5w
ZCF6ysnQ1WhswiPI9vRyrpPQWk/a50OD0eXkotowfps6n2Fr8z9U6NxIjcXxyRNY
qMDir13Bh7OOhoPOynhAbBay0My+bLizqOh6YnQgw8I78vSYoHBTnWFLH4WeIJHA
MwACf3tIGFkFmCJnfd9kGX9B4gmBd4wRfB8fDqX2kpG/CuOmrnOYxhsGqx6xsX0h
VCJEvcBfSaqMpMS4LWmT/oHxL6XiR4JAvSjGrJfyAL3HBSjI6fL8E/HI6iIV3P2l
ewVmPr3YTySkNBIjhvtJrcBoDAVe2v27e6H9VCDPqgIJ7k1JVVzcDVlwfyAtM1mP
dhkfcHA+UtIb0aKVgj7rQjbzA4lPzsz/DdD8WlM/QEnOlb/2q0Ef/A9ta0X/9nVU
VLxF2fu3qiKh8UM0IL6shVAo6g5uZ1a4SquTkZY2bTOPdqh7PsW5m4l2TYRhNtcS
qbE3TSplno5X7ZFOxLrkkOPE4ZXCpZxgezkvdZVhAb/zLqFjVCk6Srz8iXpgQpoC
8Hi3nBDM+i5Os5SWIN58rxR7rOSplgejnV76RtTymntMsdwmJ/ng6rESKIbNuB0x
ZZA6ULBUlgBn4xc9TjI5HZ5sC77yRp6E8F5LwbKCeH00rSGSTDdMrce0acXVCuUT
jGCKR2qJraNnpu5/7EIACapX7TP6jUvXf0PjTmWIfk51SK0ooRcF0SOEPrVwLytt
nbk2j8roQjCFQoOykgqCw0eet0ivNGOeKbHqDbSIc2S9Yt30zlJFsFVwoe6FnRjR
Esa+WxgESNaCE2qUnD7V6vDSKZn0DV8kheFTB4RORqMUhDr0RRyD2Ft7U8WjBKbF
MPKhOXJPqxIMBDSvGJ8iCyrPlDAx4Uh8UXR+JafeO/tJ8Io2+JGHSWsrrEzsTX4I
BN6knF0TtwIhIKDnW8x8u10H4wdz3//KEi47Gtk5a0YjNgNwCkIBPm9UmKNHO5Qr
fUL6ypnpSOYLutPc/Xu7kk457/q5d+U7BVmAgRIMfOD+4ZvPosb82tNhDWd8zBdQ
lO08bDco6+Ytbds6mmQ103Lxdo747XfO7IIvETMuePzdzutP3nDRYgCGTACieNB5
HiQDoZUUw4qWvMyJGNSeDSSaPNaPvB7eRdNIOYTr9hvj59WzoUbNUmLdv11s0iNr
KvGVIgVTZMXTSq/0YA6fx57do2MHNDlvsmI3DypwuXo/xKK7Kf1gJvW/Vy1cPq4b
b1Q+Ekxxg09D1DauncgvYrFrbMRsaxvtrX1Oibh8TFl/ZNxYtVRjPta+xqOFHzFo
SB37iAf2q6gS3Ak4OgngUdULvbutYc/0Ti3UdMUWVHUsArPNOQ4ZoUKNu4VvaHTB
7wNJjctMenVVyo450Jwxp7nlvF5WYDqc04UFoJdv6TJYJkJrcYOoNG/8lAkAau6V
UqzfTXOcHYBzIuYMIcNERkMS+ZMlos4R6PUrjpD4zeY0HXhGRQ6R8x9hLUzvUHzf
6JlCjVS1gKFQC/pB6b1FbJO61Kcm7sl6Nlb1fewTfHy+qdHHX6wFL9BvQUz7kSUw
gbMAlKyT+czC8YfLZTal52fffnJC4jtQtkrDSAt12Fo0GJtSxc2NT8Sj8x29yr6E
8N/bfTyiNrHS+kXdu5tQlMYNTgMKUSWZMJ8hCUIFBhJPKQisnxe0bX3LLXboEuHf
GhDR6Zqq0q78TpPzKYRpZ2Ad4kfhz3YMCr3WMt+3/r38CChLWDBw2V6Bd/YB8ZJE
cooJenjLookjKh9YmnW0oBo069MJYbyzqfCN6d7Yjp7/U9O5szTUXlv+VPmcSw8G
YUsIRdc0ZmvCjFswcs8fV4wKvNgbaLeOuKr11KDj5C0IdURadJAurPIPsviXOfB9
5xEd+Ihhc0qesTy2Xu+6FJmd6b0hU/F0+tEJUaCLHs1GLhMJ+rj0nAUL5VS61ItT
mGoy8kJroXXtJwORYD5vVE+wyDn2WZxKJndmvqRoEt3mlSRFN7DJyPTVJasxClac
uliyPivNDtmzOe8lmoDrIMTieeVBtR8MfV/6kQQrY1aFvcbjFK6/oSlfe4ZRQsiT
1sUp2RpEKiFW2NhK1zXeuFHAipTXMTpqdcEBzyqlA2iYlF/vukpwHZsOzo3i5m+r
sfTfpRFeu4aNsNEdoAjM2M59pLVm4SfAH59TpdPYvxOykQYnwkmMHSsLxtxKz+Ef
rncHhGlmTxkat4woEcTqOH6wOlMqjDZEKC7BgMDD30c7uIlLlhOuy2ThJjFjPDbd
0DYfIMgdGaSxeS/cu+Ju/8GA1J9PBOKkpZGl0AQtb4bRu433vF8SmonAAFgKqPYB
4d2TMXxMEPmY4wsuZxs+62wbuC2PffowGdfKVe4A0TyX6DvJG9zplk0S5XRFcSw1
nIdncchCOfh0ve0Z21nse5O+WCoYpsLe0tNuDe1VreHzD/MvkFGYbgTrr3IS43f1
3uP0qS4MxI+JAnvJz/6yHIkYm5zW4XLrILc1mPH2PfZuidElekEKd3KW6JJnr7pS
rtoo9ODz55wGuS0RvA1zOv5KsGckr2grfhjZQnnS4jELy4ML/E1V4NJKeO/73e8D
03bzjsZYtY9e1Yga5r4wd0PISTU/mDfuQJs+OEkTGY9DXJV1R5jI9QNa7vHlfiVs
5qv/ztGx/ny+efFrqJWc3cEjSdkuwQZf6Jd9UEnbgS14mKxUdR/n1FfwZjUYc81H
1bW8EXECXU5ayAJdUtt3EmH+fJhiDjt/NOTGqwKsSicDL9zRaGCs9/Z7kLasj9W5
9raOdfcJpzEHNo8E2gwuhjif7bh0Ado2F3hndii8KgrpGOFE49DaCUV9y1L+XjHA
hzLIhmaePd8naWGvf+E6rSxuIghMjwoC4axmOLOCFZO2lwjlAnj4CERxGvGOIWLe
TRvnsD55oBpHE8ej4pib7d7tEgqckMCB6QWIpr/cwouhKPGxcUfu0vVK6Jb2FTkE
zWsTV3md7R+CcmxSHyjlXFKLQaVYXCGmlGaSj9Qudvm21wgRJL0089c3YLCbM0mu
cFO3CQIZ4G/Q4r6VcOJig7Zw+YqwTvEBh2pCPVg2GbnctSa8XU2SA/YwbBHJE06e
lBGVZak6TBJOHF3Mv4rJG5p14Pyypr310zkeXVIDraCmT5Y9gpLvm/Dwoj284zWA
t4pxZXHNFafKT0COAHlGCDN6mmajdEMzYdfrcKK6qDiY7DMk/+CdxHX25pbMKUbD
qZWkhFgeNlMwKa3MVl7h4xkb0+z0drlvNNcJKaJBBHhMyqSAsEC3Fy+/P3H+EU1L
hNUh4xj5KvrF4WJyGxl2TjACekw6tT1r3Rtp6U3VrIE9Kocv2pWYOw5nR5uFaeNP
FRBlDcFf/tjOhHQqrJAng4ZPBBwLwLAvK+83fWeOOaOUV2fEFkOtyVTyFImG3fTU
Q2YESHGVWsyrJf5RH6cot0lKTD7wha2B1hhPT78D/N7+3oLU21C/CUife9SlIRsr
UogynA0lylanfvhXyqQbZTi0vANNAcuNJDedf5ktGwN+bfhBRk7Dx9BmdOHc5bMb
PynPhD2YJjVJcB5dAbIcv+c8OJ+T2hUPVMGf8NPJzIG5czjPbmv3NZM+ayzuYxOp
EG2iFXz/5UygwNEa8Hb5KoNk5QYH4obqjHG1nS6SySgHjUiwicwpn0Cm0J21fco8
n2qOOhbdbBR/beN6DvzGDCe0JPlGDzUILf5VLOwIxmryatjw/sXm/uvA7G7h+hFl
yomnXhMsOWIfA450F6jcVtK1Fxq7UB5mpE4kPB4sg9hLrpAtze4bS8EMCUNyGqwj
PkK20w/NubfwjwOAYmVlorPgnpxjrZzJTWk8SqsR2AbnM+tmwb7IdMrPJAoqjRQJ
FLGdRR/I6vyhahssmWV/xZsgYkd2rD1wClfZmcyhyAA3E1Bwtke6NDc0gRn7vnR6
179I2gXC9ve1FRXblPktxHBe8wBbF/nzLo/XFtGYibWpTp4aOwuY/LhDOZEZYAUJ
4Ff5bnGIUPhRsHDJK7W7l7RyVcHU2zwWsgPOhhuZtgMfoEf1gMhMpIdbnq2k8OFN
3dL4TRcOzioLq46X4MrbyvN6s7tvbCmv8M3akugzFJEkXGCQDjxowYQHl4zhjJEL
89uC/jAzC/QtZ/avqRri2xbF0mwJUdwpB7dp1GbciDUY3hlZ/W9r/Ul0gzvDBIOS
HKG9Q72MwPh2mIAyfAvYUXbWo6ig7xpdSCDJbF8Fnz6AsXjwFcsghtUch18BZ2Xx
dSDYDcfYyruz+JWnVsgQWJabfDl1bONMLwhNZzjaIc4bW9APT7wGm93GbVwHWeXF
kGFWBmtOzRhs3fwvSI7gsclzNs274EDFpmQ2UZOQ4kmByllx8XVdgBa4PISId26K
H0cYlLOkvRSWpPP07jc/PvONyrDm0OzaUfz+Z1HXH5PnpyGYeqI252fUygfCg8ha
48nilmRC3u1SB6WkAPXpAGtANvUjzeZeT8i/rEKNJGnODY6DBXUyuhqA/wdfpuzL
Z0akIt0jPVOP8IVPH3I3U9D3AwXA4LZMxYI9E1CROEv4RiMWcIE4h2tBcAvV6Hxm
JegdVqgbXIvxVkYdbwHAz0f8ZVNgKJzdSKBHPQLmEcM46roKF2X5Ewgu8YDNzPi0
CutKvnQGjJMGW1z2APQgsiMLv0yKnd1CHg+3E67iiI7DEYmQPVSYgPyFWA7btdGg
BlrNVFf8+Iw+3At57vjHQLnlXhbLKSo0lOiyQi/SUTIxXjwF7DD23JdwKIQFLAnV
0UxxjtWzkcICpEIia24Ul7i4+ObOGdUod5ITeBjfV2A5P16Ml4LGsqmlBJlC47JZ
lx9jITqSUMBcAZoTC+O/IGEPTcd3ZKo2tSciHmi9rCtWM35f0oWTOxHqDFR9/u1W
G+E7SlcfQ3+aipOg9a9iNe1bK2wtn8UxA9DpWKwujQwiG6RVbkU9Y9CqWD8Ajlgz
yu6R+/GlKyYVrgYzRYoK0BUwx9rBFPieO/2fP8NnOWT2uG7DoZdTcRET/cJDEznQ
VNk6+u/L8ybWJxPF9ejkfZC9lPh+CJq3uB1A2yE91KH3sgfDc+8lCGX9exl2QRwQ
wH4fl81Elv4jFWUDj2kKDfTnM3U7/soEM3P/jX8jGdtUE1YiQmPUyr/jIdQf81Wo
NggeyXKZlfxNn2wKkSICag0osVOShkQT+BkUfQU9/GAmlPzn+gtckSWiOKK23gjt
QjbY5x8Q/LhFZgLOO/fDLqyN9emeUu+A5mliqqrtia2xM5DIqQJCaS4wf3TjVb/e
gKILvavzV6oEV/eYGucBCtfxr4IGlO+EHmzkZy5pfg8ki4CWxvi8BYjR4mxYGOAK
WGRx1KEAH3lgir4wN/ngt0XcOe8a1q1ET14AmqKPxPJAo8IDgNk3wsZkBVXsq9Sx
nvWswNcbRljtguJg+gjbva++cNqs5U11stoIHkLDpjAnODt/oObGcHFgvxfwcAhj
g+6x2+g6oFqAVLBvFlV29puyXeJBDraGLlHmAlKKcXzLbo56mkRMHtMWMD7mhhmp
F7B7ah1/4q3Fepl0MWe1jtWxARCMp7VJ9gVl7cJzdqLCeB2lo4TQEsKaI1t4RAI0
HwnpM3CiCGl5PRoc47BZQhE/L+i3idd/N+bYZQCiRX6rTYD5L7AkFpcmOasfL7Tg
ND+fOq48ELtOrsJosj7yhB2d/QXWvyVTeKWDq4g6q8obMRhiR+fms6tGBYueGyu6
n+D98X2zJOgYwjwEFNiL9FqIlo+T1LBW44vgA0MTtsijKEbMmwWXskA5bhN1N6m8
L97QsCVNSHW/dhb2PEvaD9bi/ftt3qKdTmJFRgf5Vz1eb6Mdhdr8FoCsVrnpaEDY
u2HcJkGmRgR8lU7ZsmykePV7gvM6Lh+B63l6E66jyjCRlpIJnQKRg0256nXhVgCk
azyR0h5PF7ClG0/D8odCRwAlQJJEMGrQrdfYFYgQ65z8/Kphu4WOADGPNRr6R8ko
+d8Cmr6PbzFrQ9EwzgH9JRG0gBByCjy9EoF5eal0Tzug+UF+A2mj51me4U2sp7aX
m9GPZ5BERUYqnvpcUT4vHA239OdBAkRMXpo5qaqDGKNAi0oXPZSd2fqsOk5od7ek
5eU6m8kcMXog6Lm8gNCW0Mrpe2mdyQpG2SGzlDVHVKuah/n0tCevelHyuK/odYMf
BWcZRjuiGuKtODl9gnDS4fXzOw9Oj3LT3EZMQLnf7WeytA/8jXa+7adywmGiYJWe
OTYXPj5rdahl3I4RDtOJerz+VjItt35Eec0qv+QFVUlw33c1sYyOyloNZFKLSstH
+Ox7JumM1G/jhjj/fwdurnS0ix7DM5u4b2dcjVSiLV2w5ReEcZAP7AgUfl4F7BSi
eeVGUTuBi8Z8W4kuRNCvHSy23pCkCC1PPgCm8eClBrJrN0u9bkttH2pg0mYOgMGA
8ermcErERQl+OcGUR4x//OwEGRRICIiMxEzMuOy675psYdCdMewwGTa5UUTY2CgY
Sx16QvLPUG3hTtDqasgrrvp6G2Ojjq6ok9M8Khuhg2Ds+5MJQsv0pp/0V37a1Kxe
g9K5GraCvaWYqm1BgTi4W+nwixOg3i2Q9hydRfHvCNR+A6qon1OoJnQ6brFmOK1h
Kxx+lkEnrdElpFcW9sZ+ZmCIzohToSDNjeROkJetvVaD4dHNCdymUuLsxCQIUU2D
odL9RY7GTbgin+LgBVppAUSSlZPNBxjsZf3N0/iPHWExSfRJzxrIEpCIAPpF9R2X
ZuSg7LSvgYAHvk1/ccXMFrTQsBLHimMyH5+6bTVVsvCIuogEULsUbY3KmrusGfEB
tcFdbFRu4NCW2A+hDiTyx3GEixNeUXcwrj+qpmAvnry2bS2PcfXhf8oMSI56LuNv
kcV4Y6WH/NtQRInSFoZHkpP43VJ7GJFTPnEhCVIJQK6hiSpHT2DegQVQfrxugB2y
mfKgp+Z6CgSDs0a2IIFpwypF/c30/In07vUf762oH3sEXEVHNN3uUPrOono0sN+8
H9D24G93HgUDVXnFAU0DCQOgR2TxpaZZbNg7BoZxBI331jwn5gOz2A2+A52IUh1u
M26Zl5g6Rv1BXuXzptcjFvz+i/XdpFDYWrmUSSDsrhdmTe8vAaYnyfA73R30QqKk
qIeuuRCpC98IbuBk7beBhayxfa4G/vMOLpTs7Cl4rIyFK85bSseGZTgbXxNxxbwf
EuY0jYtaFGlAaytHkb8O89/Hwe0Ecc5P3sU1M6eTr0dTJaubkzbGMbHndToe149x
t+7RcZ0Tb0atMcNuQesxeHdDCeimO1NVv8npEbg5ivF1wlDa7UCf9EwXA8QSf0R+
5b4x/D0p8qMVLv8uyE16KAszXhAIbNB+i1agYv0bxZjViINMty2XZhWf/R8fygTg
yB2npsCQH8/ohLjpbG/ME6Gd3ogfoU9Au8hG5IQxEf++6tyTdm5QnmvE07eI+1yF
bSC4KSeaB7uytuJ9CPZUvNC0vMZu3Nxgf1QZN6eDqZ+KRQgldV+RTRAILHGdOpXE
1Dq5AIK9dl+9+Ywy3ZjGkWOqCG4Md6pPB2zUHPVDoNBPd7DFN0ksifWQZIiPvN/b
UWO+MfrH9o2rBfl5p8Mzle0pSbZZg9hZvmREu17MAa4tkQXduXQMiDRJgbl9vxXU
JWs1eqjFmO05L8gJOQhd73FfhCi82kTYL9soNkT/IFivD2zd2c7Lt/AHTbCke9+t
iQFxq669fg7gd4wlU8o1HTgpyS0Xx3bUdZMlRwEPLUkt4dk8C33yob42Oe9nF302
kdztJfgysQmTIzs6GWKMOnfnlSAVLS08K5cTWWgb2aHmyA6cclyTwNV1aK6vlcDo
HW2v5Qlp1T/oTI5ber3MHbzmnri3Kqc4oDSE/WireFCnegB5i3MD2LfbdM7Gkwx9
GygFV/z8e5UNezq+2cOXy9CfTyNwDMIRwIs/LCFbIqDvowLp8ZieA514zMBzaRkA
rPvOONdEPtZu0xHOfCcrTRnB7kE+Gxe4/QLqlvqAacDpZ22Z8qQUmO4vdyT72jSk
p87OvK9XWdkgJCpKDw8cloRDXv6qnRlqAOWTdqmLla/SiMsqI44zxMgs5Mju1GZL
cpU80WwkFnJ7e4Zs5tMbJgRhtp9+piS7sgHG2dbMQ0gcHrE+qJtl/MCyzPFg/nGq
D8U+Z7IItNYhnP8l9Q2PRJQcTPi2C2lZ/eLW3419BHhq9iKgNe2ZRNZdNMR3iI2o
T+lJsKXoSLKv7mnXTW/okXUGaNiedfZJCIr7xr2CCGWd/16XaX5LV4EPi7Jl4cXo
kj89FxKr65DHU6whEV3Fje46Q2vYg7CS+9DD7cun1ElO89Bc6EvaEEewgEBndAYA
UKAr3gXWK/H/5oISkaHfeQp9AL3fkmBT2F2fVkeDphO2CAYXueaQ497Wgthh8o89
8X2fslnyq9RnRQ1yGrzfzulvWDUG6WmeEQhW6ijLwRYr6n8zdYbGBhiIaAFxI0aB
B5MxGkNBMnjxaJJ8UsjCmiTu4IL02xKndjcJhjynyvvj+hV6+yetPVxoQwz2gzh7
CjowuLNwcB55MRHZkJ3S3nB4ksYhndk0nnrzhTWKMcbwpsHNPFpl4coi1raDInPT
HwNHXHwGM9vj8XendtW5GImSWFhvIeaqHBp6CtzY5UvHoJXTJQUFdnWJ/l+U6a5I
ztLpafh4eAk1qWun/eZRdg+AGFLC6ltP7bLeLJLTIcGZGHTz9qL1m/PPuCDoEDLu
XToDJG4+sHF8iqW9zHbuLGSVDtJW5JdDdXkDfJqobnks6LpQRwtcnmiFi8maPh/d
JUvio7S0XPSV70T1xNFtWWe3vL8/OatdSQr6QaIFhCzogDioBG8WAdoSBFeE0SHG
zRoXMkxIJk5IVBGe4vt2B43r2gmEG8iuEidlyv8GqeYa+w5G/o5b5jEeQWYeLKRF
SVJuzhdQx/TedBZtAKQOGCBQ4q/Eo0BCm8EnDNNdIOMgy2iODu3JOo/vrxHL4pHS
yH2AZz8cPB7MjPq4WOJX4KvjV6t2pakWrmEk+PJq/c0jo4ruWEbyOF9auyU6KzRr
z7RTfR+kfbhY98g7JVZMjj4avLzD8R2Ngd4etuotHlEgPGCkeOsQhuDbFR4TMxo/
TA4npK3+N5b2CSpcJyfnX5WQAmHDhixhKDN69WvxiueCC4V6+EHYtguf2M58wsL/
+FxvKkNe21YnJRM8EHTdS2sW+D4aG3sAL8NZ6725u1puZ/p5bzbEF1lQHl6Fp1ic
MtxdNgszsNANMF3p+xj7sJ/svCus3Awq6Egdnk+rjkPS49bkkPi/76KujXfxnCv3
AN2o1PJBZIN9aNlknHHA0zjI8aDjrB7Q6LgeKKnY4MFpgdOgELLd+MWY9JUtsMoJ
fwwNJ7LkTKYdN2NgKcMLL3YH9tBftj9APoVp7wqkpu0i5DyML19E+QXGuyy+Icxp
k8cvDprJK/8UO92LHJ1dzz5fFQIgoMAuNBQzr5JKTbrbAw0bckBwL1rpJ8ZKuxdn
B/lmbqu3n5z6uRM5dFW6VOFUAy9AKyByqBdesPeP6BzAGj9K1Y5YezQ1pnnWV8wJ
rLdxHGqf8DWH6I8GClykdwK0KP7u8ihOw3ouD4Hr7PS9/Ly7odiSW1Jv/gZSFUP0
RrZvfW/vFLJhL2Bjd7lWYrL8ijrO6Y1MWg9letvbWiSpmbRaeHnh1aK4b53OO9ch
Q5bc1gRCqReao+F/N8em5aAvzKKEEOPxuIXvl+sPWzaTg6eemxgTl/F0gCCZ39Mg
pYIKk3x70HPiQLLKM7cJ3GCK2q2U42osfT6Wezs7pkv6bUo7KJAE8DaYAvfmVc4n
P2A6wynk/6i3f5rv3wsswxoiQiLLwnlKgtb993tQeKYcDRsHHVkmV1PRqw9H2uf/
mI+gd8oodwglq7De1oyCUg8RWxPpGjtfxpZ5FnG1E0XXsNshzYDIIpTG5nL6feja
/vBIdrKNWAEN+wpEB5A554Hgyx0MjSVD9Eek8hPkbwVwABcoWJzBTTcawCRTHJ3z
uwD9vfAzsauwW2YAfWxuo9EakUkZ09sQd9rZBF/gPqBylr45l6MbPH5CzQ1VKF1y
Ncg7zZ+3kxZnMkVj4NpJQcOv1rCSCLaqTQEiAnYSifvmywI2XngrkPGHWwSJBKFo
sZDkQn1blcAIfV3b39nrp2Niw7VqfQZtZOozMyHLvBbu7e153PJw5KfK9s3KNS1/
CKSh0zoq9VL3AFSIlcK2rmVkCexhan0+FlDqf+jIPzCaZUMikf6XvyVzPDdZfaiy
sVsDWH6bNaNdleAeSp0QXnxCSbyF5eBi9geDkmfUjhoXlFhQvBpiCZHygQHj2Nu2
DTCI7UNEqiuqcyFya9zClUzjVk7i7i8wZdYCLqvj9532KgIerW5VpgLTvy9YhtFy
+jr5b9yoPweVb/aR1XX+pdOGUmz6zoKEDs4HUnQm7uIsRIHaBpeG2cv8KICxkYbX
FpFs9sbAX42/85FpD0nrPyNMwJV74SYNAi6U11iMlqmGPHmLzf4xAedJRFj+uUI7
R8sYT13zqzpkrlRD1PUOeY7DWbhdqj3q24vgRqNEP9rBiTJd4whZmWzbZ18l8fcA
wuhS28PV1XsxJDbmdtkPYqlwB1xajbfWy/GIMa1qHzFs5JO5+KYkEJdotGYzMeW3
flnx1WbpesGTZsql4a5DRWodRqBw1eTDXZFAgkoPjfeO7J+cnXv9tEDQ7lItrJ/v
ESmfpb0EZ0iDFxTqGk+dn3gbs9lZ7aEU724PgzOIJTdq+Ir9fVHoFQBcYVzZCBCY
Sxvl6cUwfB35+qs+dYT3/ZximbOrDH7gs/2BN9NyR1x0geUHm8uV+be6HbK1EO6F
B45Tl7NNkpCnr2LwMQMpQqCZV7WChnpD4eFVQnvGmNnUB7APqII4NKHrwaaErTHc
6NhU/HIUVhp0pcUfAAJmwhhzVS8ng/gsNW4Dy2DZZK/6OEHktxryT45A8Ahep7Hd
hA0ebWRHVRN7cry+ivmrvq61AYdDTDQ0xiLpaLQ4mRtMANU+a7DcZY693XYAgtAe
YutzUE8SJ1+PqKi1FYOzvSEQKl2lEfpJuV+Hzhh0ENK5YmtxYISsQOaxWCGuB1l1
exgDbrqdBc3aHFjAb/Us726Fvtw5Dti/EWMIvqKWnkLRa6wK4N8vXreYBgAOMv5i
FEEI0wsyNLSxlhGxgMvMbbZCxCZ0Um3QtwzELfA0z+6mpa1aH8J5QDJj1EI2pK4G
d4SJjC8TqV1rUNHCQ+AdXs9v8pn885nE9rAZKwEs3q8sYvy5nfKY6R+xCxykTTVT
Gj1WS2h81tRUBYkpJLnXhe0e6TFjDynxHwqlBfVBzL7zLXFAdYXxvXhpTmP2f1e+
bsI0Rmb8Ga33sR/gLEkN0Y/t4+zPiETxOqSeFOKB+YfxB1fGXVFJrTSMUZx80HPq
cPDFX1sAkwW0ouff4dUlun0Y0xVBC2Uj9J+TbOihaoSK6i6psXqOmKCJ7WLK8h5f
bJl40NWe4doQACjZ7/CwD5RtWJYWR9TgBt9LyEyUaItE7bGv+DhIK4q8jHqSyqz7
oLjWmbCnBswP4oV+MFBj5AD+dZ3mYfwtBc0/EPuGb/NapZ7/yJ3rWWVciwHhDAMt
SiDzMqcOab13x1tPewk6Q/fJ5YEYp/0HCOFUItBKW+vdqW4hQtyIkkE7pYKek9Fu
jEFhVBPvtQP/mofr0hl/6G3rJrnROf4z8rCDB8VzLdFUYHhA+kNdnY1r/zKHkWuv
PiygRyoACaUz6hfqSXsX5wu+NXkncecO7seSUyDp+nkO7Ye36Uwxih5fL+xF3qEb
3Y+N8H0cgJYRjSlC8WzUhhGjtQpe5MQAtiumD4ulBKlGsXf6OYbk3Mqv3BYnYbK1
AzUdVIfYf7XiDAgtSINAJpmDrb/PmBjj8EAqB9hFU3ZOXvuRB/oVP8EzcAMeVaqN
X4Ux0j6gBXocqCYvN8lPmVUydjKKmYXGX0LPXkAF7MizFW40wUX5c9fi8zTdoXxm
PzlW/e/aDAH4B6nhl7f3X9Ky7dKc4U/jBn8TIqgxCTFSyyFECeaJMHWLo4sDTiaC
CA34sYpyfDOhypdkocdxV+d3Gtwar9s8mkSTuUPPYrOY5klj7kEZOviS7491gOiG
Ltv+BhX8rCJxcmXSi/Cg9HphrE5Y0g4uiGS82O1cvumanK0TFGBJ3dDUbrPtqFwD
yfvLS8Mv2HDSRA29FoeB+xf0ydw15a57PBcP+uKyFqP+xtV+jsIdFCYN2HNsORiY
yaCxOoTzRt+oA4EVeOJS90WpA8XbyNH67OVMdX006CagDEUpiwyyyqZsbhIUKtw2
Ef7BW2g6y1Bc3tnPbHcSfm3cdYxtaKOBGMUIgbq4RPNB2UIZUp/eMQkvamqeqazE
MO4n1TEGhNiyNM+xBgQGElcn8FIMbJSRlSZ6J3dx1PdUaY39AHXMK6aTjpQcRB81
C6Lb0ozwkupQHMYWxs3oZMCzCpLZJKIz9brrFS8hd8ZQD7tg20+PApA7rLy9+QVj
M0KZvGez/mJQzYN2ROG4rhL8+O2GM9ZOSEBf+oatPyceUjKU0LjfaUDhpssISos4
cCJhdAsdnqh64eMkbc83AllBGh3yOfR4w/XCIZyYPcfwpOF4jhPjH+nN3C8Lidvs
j15IzhT09zDuLAmTmo8JsVFBsLuLYAAwA9MixLgMSLfskxcNzFFT99xSiyOkamHh
YpkufhAj3qu9SJ8TRKqwCvTNZu5bu4eZ2lVGOclBeou7B3TsOLGWkpKTG+sVj4Qh
51i5EE0FDb9iJh7Pd6IQAwa0VdXI/vD/+VfFoQdLkZzPzJWiUzuxE/0O/JMvuikI
f4JEWWt5PdlBSU4N5UY7rWyoCVd7d89ECLuWU19z93kSEeg9XMZFrRDLV46W4t7l
ioswR03L6t4oAR19f0333HkDRk52Q29Uea5W1Qmk/9j1YVAl0MfuRlZ04LYw4ve4
s/cfdqd2DD7uVTAYQpTD4JbClhYzKRiLiO7hfcBffrZJroKGiwJRvgKlUShX9wIl
SVYMxYCFFiCaQy0DpxfRrN/nRM0Td3+hFsiFfxhP19w0cY72WpOvpv0J/c9rrcNY
phkb+EmUKUxjvgbIYXre07GToL3Bf6pKuoKT0Lh1TzwHVPbCgosXGwXTnqhH/XZ6
ma15WA7kRxGtyL9a6R1H30Bd8MoOF1AffYUixeQ5+6/YtZ9Xd11QkcY3apSMxNYU
YooTdPpdlhjgtvx27CQ4q3dNn1G+WwbfNvIyjUcnXy2GBrEfI0+eAc3cRRp5D3ap
dipmccOliWlMXxlpEKfEprG6v8Kag1RkADwFTSCFieFRBlzYciAGCm6Q4r3foLVe
D2zcg+Ga55QIoQRkwBH66vGCgtzIO5jytnlyTESK+KoNA6SIBz2xs04J1B1P7zzM
G28nF7iEwiQFDhIM9XrhCwMrL+wcJr9YS+RpEMQLlSU13dDNG+P3Hrz0M7Zz996c
1Xl7gA966JetRTS5x7tgLOXerFESP7TorV7RxuwFAk4Xep/znyi/J6Q5gYeiL3Sf
OobnGaHFCFwGLj/FtJr59iM+bMI1g1ND+9x8usHXkF7i3oUi3GyOKUr2D43HOAXd
CfpHnMxmgh6GTgq2VuMIRr/s5JqNXzCaAmRCBUdE8uo7eAgn5dPwaChI01IMfP/s
I7tfukwo16PePJUNa8wgSY6jbP+BED4GZjRWy0mc4AZKWAvHruLU9FJQJEte3iV9
5XfhsgkHGPi56+VOaTW9fmFNeiao9ujCoZ19dIebxgE9PhxShJGAjp9BtwcHdeu6
bl5V4OU6ii0JCZGve55onjSQM/l+BsUZyVsUI3Wn7bze0gr5pdD4gEPIUaPvLF1p
N5xURQ4js5V34HgZZHUXSLjiuyUHSNVGVtQDfyjlBATWQvr3CEFobXwIZhqH5kUf
WFkrILwXmpW5DPh8aM2toUcXsIe//hOE/LCrGGUmCrlhp0DpihlqV8L4chv4zdmI
PYqVUdQepzShGO3kYWx0Z4XM1EaUfvAFeiaae+tCLnGnxenu8FZWgP3WQGk+UeqU
wvTI/FRMbPJXHniG0zXH5JgzyCElKCQ+AAVO8PVdqp4o8M+ExfIcHulYImW0eWaw
7tlz4gxwJcQvS12+vSvwB2DQnWn11PyrDWjufwqalfz2KDG/X/yRjp1XPYILSzeW
qrE1R+R6VTyKTHI6Yei7w5INxC7vvn35TJn/ZL8U82NORhZ0PLRIKZ9u01EeUVxS
QTsPsNWXfCfgVdIaO0+MndQSZhLhHaP3CPsZEfkUXP4htGx2C4fGIyqJL2oD44N9
RGj/8EnyDNGIKZQbz8fDrTTwGvkXysHHDms5S/0E+zzQW9HSwSfcvF9UWgYjLD+J
KsAW/4dg2kPRtyhn/vVAfhgF5KPoifGKZ/+qwkJBbE8TSRclW6J5r8jYUnmNX8iQ
rY46tXpQXAi9kZCTv2j56UJ+mZtAXcEavMigA6lKPkx/d1g+Asf7qdvdQJAKbZL1
fAxp+qtFA2hP9elHfs6EoNtafthtA4fX3vJb84DZXGcw7KZjuWvi1oXY5OTtFqd7
dJW8yFqDRUV6sNy24IwMvdzn0Gw5iH1nIvglkLHbu5Fp2I5XVKKsdnofMHz9cXuK
y0wPtQCHoyYMgKm+tIjECoG0L3orAcFVbvnmknorE0L0SZS58QbIwe87r979Tfjj
91Cqa7tJJhV+p7+EDJTJuvfX8O2eLAZopxHfr0tmOZE0AXEwKnl4ib50vdqC7KXF
VLof+iBlHOQqgrcAZL69FefZYEnkMAQKYn3y+02d2PYOAjgPPKCiOPAi838m9VsT
Y+snHkMaQimw2SAUgV+toDCLGENMAX2a4VFVh7GTrrsUMyfKt9lpNGnvOxvLwNN1
VnIAMGQ/IPMbT41lxlE8tfRxgRD2FI5x3ndnU36wl9Te7gaLbeq8WVmBTktAoFdL
Hu4mjRubT9vVz7UB/iwGUgAN7Og+rTE8Om0n7AXc4zwXGzc2a9uNRTTinEQYC4P5
2Nc9PfKyUKfYMPYPQ99b2fUmSp/zSkCM8mfE6Qu99uMG9gG1GHgCmRVrF2UjyLvR
Ele+mGg53Hebrv0WCqHgVZSolhz7E7CtKIlx87b/I+hmRaVTUdlNqKIiGSUyoYot
8K28JoJpXHlx/O/cyzjlJzfM2c0d+b4dBy55vFrfDeX1hd6IusY4NbM/BdGSRkdv
/vui8AE3Q5MR/Z2/+CDt+MM6Oa2xjwGwqX42P1mkaAqBP7o8CFLhKyuc74znfD0i
PVGDrQ3X/1JJV0/MH7u8b6JPHqjmGoHzhN1mPcPkJQud/q+aNCUlxlxzua9BESNX
DhO0Cg9L4jjM6OCmpAPBG3D1y0UkcfsZP+gw/6frspL06rgZi8C2JUhdZPP32aq4
cR6mDlbUZ82FHExJSQW1H+3OM8ckoQRNdsbaViGsCGoxATwDNWBavQfBpuLnLZDE
1aTT7GjzW5nU7DkjM9gg/f5wcuVGvOJXL4hSdYYC4hQA9qqZYFquMS2B5hRghoMN
A2E8v0Q+MzyHvpP2TeYxpLSrK3BNtgi4sL3kM/U1KUCB03qd7mnzv5n3hRkQSp0F
8pSoyTcZCNwkplVV9vi/bRrxYoJT4Gqe8F/Gyxlafycrb5e8RVnZXfBz8wBrk8R1
c/r6EJR4gTLNQwjFHaxpLFieoQOBo3rSh+WxuDVg+9wHnqbwUuBMD+n1uoywicl5
qFw7Z7D/sB7xbuwdTXdYKkWcr+FOnqy6taHBj7q+sAoItXG+HdPTkMwKDf6iMzo3
h7QdH+irPlVm4bBYVJwsiTydn6BCnqv2WbkI85byFvk4fTgDh5lt2iKjL2FZLHI2
NTNXEjFtLcptUpUsEyA/XM7dkRbqfaYQS9qIIU+1QUcMgdhJ6kpMDBFpZITTuKz5
kVs+twMHlVbGGfdUzZLnn45XLtnLT39O9brZ1k1uWsalBFlUkUT517n9NNVeL1jQ
EqWio23B/GSGLZKxbGT7nl+4+F/J1Dw4RMMp02Y8T4zQ1prk8TQVk+az7BKa+BXE
G7Ao+9uDShJULJr+nT7bO0z3lTV9Kwsxd5IZW2w2g2bOmzB7yc2zG7RVQ7SMJvbD
BLjSZa0H0X+4TuM4vKPIWHZfOgovZKzIfnvnvLrO2gm7WhzOTaewvuowAfuYbbQ8
C70AzzIBEpBsjGcDPt+ZOgR1oIOjGFcjz+XITH7rdqgCe8T7y/rZtiQM2Doi0jOl
SkCllzqmsBY/9Y7IdMYDq5enRXUrHgpVValpuxoTalG2ZzmzCkW/Q7MFWFnEBo7d
NhYEE5cMw4FRfommg04W7QBMhFmhooWBlpCiGTGAHg6hM2ANqyMLzuYJQd0UpRlY
5/d+fNeWkYKLohAXbkVzhqwOZpmKog1e9V0LjX1IVJ3x30krYzEEQeeC8iaXiYFk
uwjHn/Y267KHfv2o05e2jVpyf3TF3H5H90eHc2n71rKFolQ72lXaIJsentO1T5SQ
uZTY6cqA6Zd3QKV+Hl9CMiDq4EsfGA8plyRlzTRe1DeeDt7c3BRz7pM7mftNJJ0i
6ldmdPn/JOLTKuvi94uHjw2TXCa1XnAsFGmopwI4ZAdlbhC10O4o5Un/ltp7Xoct
H6WATEUm29mPj/ZrIkyvol7WCrA88827Iaq4aghmxTEZSxnmU4uoxBHgq5hbHFNZ
wLFq0OyBQQ/NhPl9Wz9bjzeHDjwdVKOn4SEL5I6Gn/n09XjhaYDRfXdzNPmnjIwq
Zhl/v2GvYC8uFx2T3/SasQbThplnwkfbPLfCpqQikXxyfxjCJ8pzAVSJWItpZaVK
Hn7mKl9ob89Zy3ZCKAnrZC308DRlyznl7UU+eoIxF3wfs7AlfBBteiIgSbEdBfAI
EytzZGO7kphcIqrjCClhwU3oeN4PDCuB2UElq42zhaTEgNbnPa+aMPxZCM/3cy77
58USjHwxkmUys+z7/dEcyrRLhl8FtE7xTI2HkvnO9+kk7VhlqmO3klzKVUdTWQmw
qxACljOWPaWRmjNEVPIEYRdQp6YC+Ci9+QNtTxC2i/rIucixXKqUJQPfGV4TOmDK
pLE7A9XgKh3jOk4Ede961NfW2BTX7L+FLmFux+KGJJ4zx6ko3j21KqDdWG4GzxmR
oKGQom8bhrWXF8obE0EYwU8G8LL+N7L8+dfS9RkGPr01F5g7PKKgCa1yTpxgQWpb
ZHstTo0g8GLkPr+uL5qGbzoNsKwGHUM8CWoTaYHco8TUrs1VY66Bg8316YCeLVLn
fRo2Cgg1Z9soIHAC7QKS88tohLzSCgnDzCR4XKp1o7zMSi3pDmEwjx2PGZQhH7dw
XXBi+0SW5nfVw+KwxNCj4Glw/cryxwaq/sonKkOd1r3TEjyWv/5b5tJbqzcfOkG5
vYPJ89TXGRw9JGTC7OefByz+gyRR7XR4DHJl8A5Z72icfpXG1sZ/u7yeUA1Adptd
g78VoiqtczKipcr4nuw4gUBGErSKlu6yhBSR09afbxu71b7Aa+KiiqoeJzIXz5QV
5a7SWP1/pZPnuAYEZcZFuSnUegKmfbw12WcsK0elbZO8uuuFPonL/eqS9sxUoSLU
qhuHoQEMq4m/1/Y5O5d9tNdM+umV3ql8kwFdgFMWJpuSJnKJXDbzmylENBiPdcjF
kcLAt3yQh8x1SjijCST7KMm14j8lAolBHNs2n54ot3K9vRAiSvPvDwH7db7plcMz
TTWfL6VUQzNffjaKh8qwzBvSeJzErQnMTb3/aKVQSKetyIvdNDP8nEmTaZSw2f62
hdTcuSbnD3R1Cy+gTyITiJ9Y5Z5m5L46oFH7awpbSroO8+Eni+4OQgfn0PynGJw8
IngASO1CYqrdVA6EJ6orvEtxaQsNMOY4soG+6uXIuORdI730iXp5ZTp57UsFsm+X
XrLdCHQEAamTXXwzdRPwvlgs5Arr1fro/khq4s3F9HS+jWodL9LmjWQTV92KTgpo
YGL8sWHDCyL5FiIzom7eo+acwslVKOIawaqXWPQeHQwRgOaGzWlsTS92Rro+dh/S
s0MkiFkMvw8JTuitvId0S3rf3DbLxpU1VNbWX5FDRSYE1Wi3E/mOAgrlC9D3pbNR
4kQsE6yAonrtlNM82hnjVzCoCvuK6N7sh99kz6bYsWH6fP6Htb65r+0PoEVpMAjd
E8bA6SgsX9Bv0LAociwXGPnHhMD21NHoJ2NkpYJyhXho9VRHtDa0fwTGzeUJu4sh
h9f5joJVSy+APWzZFX/AvGqnjZzNWSNEcdKC0uuf3czNCwc1q44dJSGzeilSlyTj
ardc/Q9pjMA2NzQuOPjyTw3L9rIl+iK2haaOACNpuNxLcL2ejxd1mOgrPyvhXVsr
BUuypc1lud5VJohNZrczzJDkecdH3Im7ZbSTA9mHtjwU8tk9p/twB10K92EEtMNF
/RlzK+fPsw5XXwz4uVuplmUzIbF3E6W1Y4PzV/sj6d5uPn6BbYt2XSmiWSWoEaa0
+miPv5MpAyAwKZnzwMnMRb27IpvT2/or/Es1FJ+haSYihrfLUHZjL4w5TW2DP0yU
KBOZHdLroqg3hLNJcjThsOfoOV/dYyVPkNaM1MUPIFqLgk+OwjPWKsuM3ReU7ORK
n9Bvs/rBbULe6bvKNep5CWS+3Sh1ZlIRqjJFsIFbGQQiv5p7OpFEreOO3x8Y+vA2
S/8zwCk2bOgp1U+yxApSv4P1fwnhx6XcdIesBUw0c6++twkiCednwqdPNnTl96bT
zGymsK6IvP8QQ+CS59YvMS0EQkfVR1xyt1wpL2xCQBtKvCgozQFIwhNXfrcRqHfW
xoqeJWho6OD62eWQsupM5e2UIFJAZypL2FDfS60QwXcCg4u45SCpWckDcUuPMbbq
t5GOXLHxDN5qIW1QRMQy03miulm7hnOQo/qFo2NC+I8k38104/YJ2UnrocPSSE4z
F2Cj47tA+CbECNfH8bTFb6lYRKeQTzGE6/5McUg1BrdQGHkf5hQM0DNpP1tto4NL
Mf7YwJiRugdn4mQxpmPSiFGScZDbwR2ZmkrvPl3pmphW5W7Www1Qb0LjOHDeAEa2
7VPquy8wocCcl8QNxXTvsSKrzHbXrDSP2O5ztACZhj8GBnm9cbe3sXN46/XTukyo
wDgpmUgMkkGwMVCdtdS5l1O9+594mH9s2Syz8qNSr+N+tcsBmjaxJn2MZo91yEO9
vXxAffzWyx0/i9qibTcCenNB6t0rD+L/XX956/1+RnYrmGi48en0C6Tvjx4+B15b
hqsHVuQRTLzUvuhTQQWmfP4EvH0Q2t77a9yjr1kiD8wUh6yxzNSX3HPBI3H9PO4k
sfvt3OmoGl17Nu+aeO9kq6kz1ftrFSLCchpgT2WHL4z49r7JQRJBlvZaG3zgZctS
60k5FD6lfp1UiBeN3oSZ+JkEP/kASiOavQt2H86a03cNhGSij7rw03Alj6BkHGbI
Y7Sqv8o5vz9+kXJJ9YHLNZCfnehTm87pNyQUsOQXtXyhe+mN1BjJXKeq4+HVBePk
lNII+7DPP/6P3nPBXmCx20orUhZx/84/HAb5RmK6RVh29Nn3VA+eh+WESEaNDA87
ceSwjogdXPjKxpWioLDot2RUIUwQTjs5dZ8F/xkmamwNpKrbq7bDGWaq8DaxnvuB
1MJk9patxiC/CmY2EYowgKIiYV7k3H9oT2UaG+UIcCcbdLQ+4c/ruRZpqQzgHHaJ
GdvjIOEcDAO9eSp8f//GNIbEZtdVojI0U9BrZeddVr8rEfAopN6++UDQ2nHQzVjQ
9IceWcihg1/OtkyzXGYZ9drmN96quSxokcdc98OEwaWQqf+RgCjAfGMmROxcF2V2
/JcwYioXXF1fDC+P0HQWahrvFvVeyZRxTrDFCTaicfrDjqMcrvPcDz3FkI35LoHT
KRZO4FnB+W1JdecfuXl+texaAPaAxX+5jtfEvX0an3P6kjCNVSG1X2N0cydUMVlm
//g7J/pyvfa7gGjQLSzizLdVvOa16wCYJ2q72qiOrLPVbYN47FQIGmzV3eKCf+bv
Y7x90tapTVm5QODtmZGBNjc698cRWhAObvWiNJmDmhzYJHGnuCebRUM01TVaaqcS
XiMP26LpBGc+GrnNPGWgoD7mo9itjuF44oFMB8M6VItmorRrmc9bvVhuSPvDXI/W
6ejJSniXdU+knsPrEYLr1b5dWffSb9V3kNVCuCl78OfT8ZhGpOKBjBrqeAPCCA2r
ZP2pVgISesG9Hu7QPOd/4eOJI/IzaI/1bar9BMpCgdxffB50gj/YEc7yZ4YItLgc
a2B8aBHIBWpxqKAGXXXQaq7ogSIu/NxqN5Rsx71UZxR2zaaHQ3zosZaAAgp/pH/B
SSdd/yA+7kQAKTZa0uKDgk5KyGtd04qoMZ6xBg56/D02UYwuECXOMMsyEoMpiPHY
7QuZImZNCebmBuFsKJMX+cofXHQxcGcdAhdPkWEWfGSn3f6Yg+4xCGymBCMNvWqc
5ZzF1te6X3DxzZCN63XsxBJbJOYfxM3DgV3LPiyxrizCFyTOJ4SiakpNNqvvd1a+
XhZ5IZaY32lCUtQAYmKZ6VTeIMM5/v1WlvNK4ivUnP4AMk1/wCl1bpYZEtGT/Qdf
dl62V1dAmA/VGh8Er3EGX03miUaob2STFV0Cv5p2eOaUdsleA9xBH2E14uFHQtTn
4Jl/3lpKBa1SVedp6B4P77fjrzaOd3Lqa2pXLttkhU24g17vjmCuKu8WpC99n8Pf
rUE0a1J8nCtGQ16iNxHQYOwr654d0Bdfn4jzthRKQnjRTCPfvwStK/o+DNF7o39D
eZiimpILW+ripiXtwfLEMvoUakfn7+L/9Id4MoGLIFP0gohAoH3JieQotwSEJDe1
3UU+8CVpnyrFrlIMYFcngpUE9Vkho9CvFMYB4fcaK0zan/U0mseGYzVKG21MILBw
22gQn7gI4G3faPkHSqPpVAjTMu3fKpn0fwiDZFAnU/5dJSCIRhkLmeXlu5LKWq4S
Ko1dgI1Y6Eb0GYCphT93Mj3xnKFNLzgN9WM2h3m0I25DEYR2MO37uIZy6VYFScCs
aVB5zc3y0IOGcZIiWCUVEcvrwX01WLP8E/0eI4o3JfHC6fFh7M5+gb+bKka2FrN0
ghazIzeJXIPnbxK4SGRIilyU+W+oLMHnAFEJNb1XtXtL7N1tCihGjRssJGkhN2r2
fpMv5k1xu9lTGKNTIbSNFHrdjmqIQ37p8XvbTvCR4xhFPfNX3WyafNPBaVedYh4+
5SYs5zeWQcSfxK4eCZljDC0pRyo4wDfx/Cgza9rOKVqrRfe7rifZqmHH5a0EtNgJ
S0hiEB0ac36ShrWkBdhPJ1JAQHXLtFe0arD0l+r3CYXD/BqP8kVAKh4QyiBPIrmG
QWpEZCvNzBvE3w4CQ8Bkw7/alllU/58OLvA6kT9e2oqrnjTgVGDIvYK2Yh1TKCWV
fIxmlprbUvKSS7gfFRAlXeo060fy3G9Da5yZD+hbmmnC/70r+GqBnA2+TOxknm0O
65+XdTYm2MrUWi5/P8Gh3CK6nFUPqhe8BnL76du8ndr3ibLgi1nnUPKur0Sxiswg
befaCind2OWHIgFyCcngZB83ax3qr5D98d6XiLkWOs7Rq/uzYrq2H8/RC5qVqU2/
acJFKbTugTrKrUWOYhUIwoUY1cz8yY19PAi8/eGehQisD5FpVXyeWUpNuwP7HQaY
OZFm8G6cmq+Rqfcs+tvnRYwONSWBHesa5JDoKuA5lhPIEwCnFg0oiUrYHrcqopz+
fA2oMaxRBG1vHEkskBO3mGrdEyYBECz9q2C719Dln/i8kJm3j1fFIMAigfxKHrcN
v3tfqIEk+BBRpq8eiaA5uQSx2PuyfbywzqHJOuRLFoSV1weQN0Kd+qXLjRNT5/KI
3qeaaZWVG1gEs5l6qylTsc+TR373yoQGWSMSupFIHnRFoBpmhIRdbf4k8M8iWj7n
yaqpq4m/FHyM2mixlYEchHKokTJm163aaUkPJOROxL7gbfDEv3STcycT32eGydPX
3rc4TCTt5FAHLmzCQODouEQHt3fGDdXHOk8Vl80xgjoNTWmMHvGUzWPb2gvos95I
k6ancRMzNYR1z0PvAuiLF3o8BS6DW2h6vl1bgB5Y70SD8amjsC3mopHvoyf+E1vh
TCcrGI6DpF3ZL59Xy40be0c+KzvUcEGWvL2ytAZzb0Y3ryb92ttsdLzxc0x6JNz9
Cs9DV/ICcxTkV1taxj5jpA+2j/GSAJxZ3ZUFQiGRkHL3daelYzxS82HU5/yhfFQB
2si9BQp80VFrVD61/DJtKxBJtedOEO46dUUnBdR0/8dxRxqSClQo5F0hxUuXe0Pd
I3cMFMoNt8e/kqdS6SLvOKokzTbpki9tO+JBLuxMEde9Bq0ZfCfqJuF/2coOH0dv
A7PdooFgVr8LtVLwFDbniizOqvtdHvO8qMcJtMsGhQv03jS2jtJdcZW2amn6L5XA
Q4bxPWWuc8NO0x1zUjdv64XXnqbfFAFay+zZuPQvui7STq4XR4LPBEYOwNY9e83b
RB9rtx8hB/Zz6H72cFt8FhPFoU/dclngVBzW3YfOSET9LVogiA+Gq0Dm9nE+Kx07
N8DeCG7Sg/sT/f0AXNb1O9zv9OaJpxMRWU01ftI5mZUEXgt3dXJcuFzJF/IWPNIb
L+9CGRZE/TOBWsNStYAheEeaktzPcvBr9oNsoe+bI3LVl5V0vD9ihIMxmO+RAUHT
iscCsEPgiSYLwdr9EHjqxDfyVavKKlcLXmo+jL92vjadXaG5EyFFl+aDgsTvv4od
9G+6HdQAtA+symJLhY+vkIoTMCtArzfC4fyhtw/SH6ER/NSrvOBXHBM6yNSdq0RM
ybx9Xc8E2nGBRcLQs9VwWFkHNAYma/JJBhYILjtrnX1y3aFv5+XxoYXvujZJPXMK
sat31axRpnpismZZkgCboNKKfyhLHbaugCPkKbsJOq+nwLYJcEtpE/z/5PWobiK1
GJ+RfAicN6lJQWk2hoP3GladSOD/qYFt8M7H8tTzpNMI/s/T2boEBE3A7wplRlet
oOVDBq9Hmno7cH/B1p+hkT9dCvn7Gt4wC6ynt2u20BhKMteRnU7Vk0+GIjOxipd4
0TUPehC+Ctno4RPuQnLY4v48PtyJUrT05P/G8VNnC2WkOhMzf4lf6oISjpMKfO4c
Sn1/5fznIJaIUWmrCDrasfbIiTtuSd5dLvnObn7r/W8W2tqKSdMEkAJL8AdRPUB9
pj5XeLrfamnBap+hAAIDUNg28MyO9hpkYv+hVb9GdaEEiPUiHnnqV7cbEZRh0U+H
x0Fn3YJFtyM4Dc+5dY6LiwK3b1tCW22a3uawZfwupd1RLqm1ZTIBLwlmxmga1e5T
PBvnH1TI1XLGa4Aa2EnwUdkyM3BWbWrKs9xG5RDE9aCtPFax5N1mH24chtLk2pPl
+9ts7f3hiclUFfXNSZUC2rBBjQxUKmLC0RJAHAGYl90dMnZJe3PgbCsFr2Ds3ost
Jso7Vo63NueoKLu9GJECsD1LXbAozzQauPKcFtNqtgEWAVhVtKj6DEu7IT1W+/1y
oFrfPSqAjFJQIBeRnprnKHyufJUEtxWzHTCU0xBLZO9OFx/bjuD+nHER2vA1nKY1
2itnAavQHsi9Y5SvoPgnm36JkEJikROILWhmaLpsTa9mRrt3OezlmtGyFVCG0+8A
Zo+7xZSdsbQ5zmsfXWEVOaXR6tD6O3ExleQsxv3ec+MWXnSXHR8z+6p6B1aVV4Aw
7tVsyd9jylooed8ddjsBIkqt/FwBnmlSU6w8ve3ajsvTOlkIMYIs5XnqB+1rCNKQ
5UZVscYH21rDHSHh8YppsrtVlRNzts5w6LDO/6gSLfEURZX5VqVMmKaNavtsBhpD
4TIA/UOnKrjqEL4wyv2zJ/NWK8QL7duT36CbrzTpwOEIJmO9YJJyCZ41rMMixi1k
ICQtypp15IlUC0h1n+0Os62Orr2RNECovNKsxyzrpDdIVdrpXl/pKTaT0m5X6h/Y
R4WmdlfObme8W0oxn7fTqqfW+RWwUhwJHPotQSNseBRmYkgcuGO+fd8GMsaREZ7x
iXX3RxnYwzq0bGudzYpFVqpOw+2PLEOYWCookvwx/XPwZnrpRhbgIG/zbeRcKLud
M/vDMpK2N8S5QS/gARva4McEk87MmZ58filENJnC33t+mh0Nd3LVMopXJknQxo8I
I4tWt8AtWlHEtwzMwvGu7uD2lIA+Qrndh+K746asTQS1FaP87paE+hF8+Qvq4ViC
jkvAwPNWaDlmDshuEK/ruDSjzDbYOT5wL5Y6xVHodgwVjQrDJ/Nq9BU7hEx+FipR
8mvUcZE7OcaufSX8LblZ970NaCZkmf/x7937KJAGzN17jIFgPrhRcs136WntCIma
OlTf6bQB0M4ItuH4rCLusQJK/Uurh+UliIzbm/MduzeeqGYx7sIBDHfHTZ6mbWm8
aXCT95rVY8maoK5vPLSkz3RgHDam21JwRdO/MOO34hgoohYJQGf3C374c5Rg30yg
MG7NYRJXEpWdd/QtI2ABLRFAME6MqValwtZeJ3TBsbuM5mpmXhnGSnEtBgSe7pdo
DbXCyOXBe9wPmfjI46ZuKAtNuHQoFVMvgCb02roUiZU62kc/COQjDQn9ZLb5mXT3
SAV/D6yYNlhlgtsz8HGjLhLhKfbkd2570xvW4gNq/aOOmvIxNZQkUd9GMxignSQ7
oFDFyNXbq7xOOHxI1YRRrqh+Tn6N10dNXKm/SUjgeaNLrOXRB/FirwforRJeOJ0L
R7L71uZKp36PdjH0t8LyqfxNgQAx0JMTlxMr/HLxvFUCZw9uvegx05I2ve9KBsAI
ZIpwgvZ98a+N76Ky216yj+6jVjx3ymoEjmEcTGW+43mfLOidxfC7TIavYSORkSij
8eLKxnyqYumgevqrPqw6xsP2tXK2hy/mVwhcMnpsPtpOOkhFedPAYWa+kZY5UfCG
oWm+qUFsyV536h49pjKFqPv547kuyXs96cb+rHySNc8Efw2U8EKW5tYJGRFL4RFb
gxro7hIzL6rhH3ZtkMcnxSkRuKIN0eeI4exoNQ4LaCb2osSFBsDMsVeJ61H9DHsy
E5oJB0BjbUIvBpAYBG6ZR6z0VaokgBqoAZdTtd8je6GVni6SIfU4F4ha7CYsDoCV
eD+IUBmSwtEMfYc0L4FCvBdLohHCa8dNRVFKKtGOMHRgAg6KnAM2vOdH9+9eY1v0
3vdkF+jZV3VRS4APufQNE1kMLRvCFIy8Gt0KNCHBIFEOokYgMxosIDvRG9c7KAis
pyWPcSjdx/FqCjWsrV86mRknuYC0VRmJ3wlsDP8TjiysHPU6LxxHZjfM40onFvXP
dAAuRDWx3nrSuMXaTGiAKNy55xNyMiYQNOTJ3SRss1cue6hsZtqQhPlAj5mODKmK
2+D3sxqQ/SWhYpHsjzEdAO8RR6tiDZ95GJ666UsT71JuJN/6+dYk4m2+RmKK8hTk
OvfAFh3gfamTJwQdolCKVwZsSz/KhpzsqPwE+giVoUnv9MsUXmn1gdnTzbsYRLli
QhmPokX/nbzDmLN6ZC0QnnZ1bXxR6Rw8l49UAU7f5cVVKUBungqNfUGSnAjrpHj0
P5amC++UN4r2poSTEeCuy5OGgofKTecI0RwywCdnMq4j5ZMZ77xIF3+Ep4LYIEc3
nnxfz0ZWkDp+d7CFsukrlsHx6ouNqPfv/LvfdACoyiG9+Qx7BrLEVk1bjCk5GSVB
DgonjK2TA8a2Luzw97BHTYcJF5qHUhfz4RtrrT8HB8zUdEmys3Id7DeSd4xQsbMv
C/0F3R7F99Th1n9ngcEu4N0091nFLWdUwbhmfg2lZhXzZExuHxHBsHMWzYL+GLUZ
daPFQtSWGcqNhICUTpXRVAhTte+L65BVcPZ90DzGmSbvdMmw+tsYUENURyOjqPUZ
702atMfq/gfFQm8bOlTjOB83RRyum/pOIfS6If4i0QDzbW1jDbrEnPk3dhvVwERZ
MILCalnQquFC2u4XByn8pyFZoJOP9ryolvMJwGIRf1RlKrx+GOVfi1x45CXUzzR1
CSykd2QAjUoyG9bWkwmAB+hXSp1eJbuQzg9H3gF7SUblDk7Qyf+3rX34jrX+nN4Y
RLcqXlibyNhijZ6vb6BxM4lAEpNqQGFulYtHcAjc8JFFncMvCPpu7ZZAl78I7Kf/
WZnk2mlxAv/PlC3Oyurq9lIJ6+qYtcscaxItm71+9addMOBXyz9HOhS+fW67hvk4
XBAV9+YslTt8x9M8NBv3MkZsXx0kMpu+riM9RUTjbKO2VKLJNPf0baezPPLxo+QY
QydZBXgNf8phSiuFZtPp7Dy1V8tDXIfIvS8BzOWGrA/1Tc9QBQvD0CV9COqsyj5y
W4a5CNpPUmufFNz36H1u3kRDc9XhznHvKhEtZIreQvCM3du/ud99E5Try5wlEmst
WCOGUXfKLxj3qF3467lquDMNXKmBTHaVtfcYn3ACLb4VSTWrj1wO5S4dLSlQjHA4
Y9HOvUYsXf/cHzguIB/DVzz8LAMeXU60SCLxW+ZuiKXic7YlCWPu9xF2LPkTVwQ7
VAQQBM1n/VXKOA5LqpjDOXFETjMB+G/D3NOfItz3EFZJALKazkjkYafCVxwmJVcl
B9ycKk9wZJEHfdQggzq690tM+1Q9VsXf40D2Qvb8Yqtrm86LW4nvtDpf6aIv0d5M
03ylsTadwNSKsuEg0JTU2VkKsgYgESw305Sbh330WvtwGE46A0wGzCkznwH+UyJc
s86JP7i3+Zo7viUGa0pbFcJ9prUrEbjuVgfsVCqoOdtSGppo1c57ogdpHjIb+DAp
lTiMT/l7ECASqXd9iuai1+602NgExnP1vm0QCdj2oR72yVcJ+/aauDT4GVvNMclA
4v9zIFxdUPs6Df4yjUe6RecmuFJ/3apRNHvb+U+You/gALI49IHw/mAgMB2b0X8k
jmF/XGcX9q/XUdDQW0/t0v0jvj+Kcjf6O9swW6IBtTcE4/uVXaXna1NgcomNIeTD
spapiGcIiTlmsfqqX6KWsbS9usG8xLJHpUxqF+YMicxfcYj08F0k4WN1HjKUDCJw
CEiSLdVcFkNcm7qRppH/SJtdSRfY3HDxS+nMvMy5PM+Xvvc5XKnIKTXapS8rKeRe
rl7dot2G/BkO6srxxQNOjMYRyERnReEw8zR0aU4x0thqklDQwl91C1HbJF91S85z
cuUoDIgfj5HRGozfprdVF6FECrP7+b9xuZCTGsPPfUxz2hAWisYAOPt8qMFI71Zb
T09wAc5QKFRznDGhnR+9xRaXd8JtHqYq/Z0mtxCehH+EKEygXxuaj97X9akodz5S
yecU8KsDdhL1JyjXz5Fyvbl/Dv2EtxjyqQDCeLE8PpLp+7FXHjySJoXBW04w8wPX
R/+bkzOxGrpi6TGN7rliiuSJBHaWXjLdHH7ntJ/uK4OrDTzCTaOEkP0BjIJNu9Zk
kIV0a/04vGhz+d1IDQCeGrhJ6JeV/UV1e33kT14z7L1QEeamAVQbdtFqskM+DUl+
fVY/HM6TgSmPoaMoT2EYuYQtDubZt6PEQ/jr0WIkn8Hgz6Xr3EYqOzRN0mwXNjZb
5fkbNtNtxYkWZXEeAoP/pJPzlo53L9ruUcvHtLUOv9oBCEd7gaAuCWhr+iikh0ia
T+laZ2xkwJTPsn7xIf6NFF1SxXeOLu0tDyMchqELELg2Sy1jgK8vRCTgTMoip+oF
yqMo2OhK5Rv4Oj/UZ4FaL8YlzcYjoXzZ4QDVLnJD4ryLw8AaGVclAl0BVQiD5feL
KhUlwygUfsJsl3jyWsdHPDt5Ayk6zMrqDWjozC8pyTblP32d1gdBIrP4YQIoZv/z
EpNsFR3f5G4ljbbE6nb/Dtd65c2xDtZ+993xbX8/qPPrQn3+qMmI2sXURHIKHxDc
xC5FUhi8DNx89HXiIUsTV+U1OVYZ/4owh3dzjIfRSrvrmou/WrIevJVPuii3GXUw
mDdgtYvyK8wYIKpl1uirZLmlvCe4CfKhH4xtZr8lGgEDe5loGlofvO4i/aL2DNgf
wamXEPuV6N16UcHnk+Nwf8WlY7Htjesr9qTS/LLpzV9K4+DKhZuVq5cf0JVv+/66
5QYBjj2NAg9qxoTcbee/fPq9BG4imypCGtbKp2PwqSgBShucppJrOHZ3lpDWJWOQ
EYb+AmI00DQXJsgC8xzBtjCU0SGqlXDZV4kqdI6odi3TuJFSmQX45fSAuZnhxwB9
4nuuws3BJi5p9lOF0nkTZ6qH0TYyIVhHR1s68ZarzX+STjXy+P88/t5eq1b8Fqg9
QHjMSgKkAtHNNtue7+5oZKUverk0CYzCVYcOKvssEzP05YfW3v5aH/R5Be8Uc5D+
SleJscogdNG/xZSiOSUydq7S5giGUGIKOHECORccrM+gDePP11tEUTNRZYJxz8Er
3FySPCydAVzExZWTA0yw/RcOUs2oxLzKslMOFHSBxsa5Nbj/GST+EQPHp9FEdcCf
qQGaQ85Q3oODJEpG52cSBUjpkb5NYXO1mGm2zuh8kEQjLdn96VlpewH++YDlI+k3
FyVTR+cu0seWgQheQkfmWCz/uMalCQqYtQpDsYC0pT3e/ZgnLjeKEjLWFE4g022y
t6XmSR2My4L8DZklHMcnXhE9dFkmpBNL3LPhP17aEJObRAw9Q1aFHEfVaBZ5v1wb
DArucSByO9vpJpZ+FMbkgDvtbegbDOr9VKfcEf4MiW1StnAQWlRWTYgw89ocvULM
0/rIfxGvA5JI2mbitGF1vJN2AOqmV2zUX1SphY78uSwKZbFxXIKtiMtCg1tz8cMw
pABM3zXC+Ifv8hSK/AXIW1L63qQZLehEGLjxEhzr+BtYmIjQ/SpU2VYSO8jVJ8e2
JWO0pRBM78OarsGXhNGRqtsXqTHg/pl+hDsQF24mZTj54ZzWtTdK7KYPJk7iUgd5
2eZ+GFB+UCcWDUQJj+wm+vaF0WYkOQDTZLHIufME2EOYD8JW6hrse68nzPlgATsK
FvDUgrppj5vq7chvhJNdK2hBJz5f75siDPGWooZtVl2dsQS6UWZtOj+b54MJqm01
0nYU9vSpE6zOjChEyb7RaR07yRXc0WKc96MntNLFgTFwwOT7wAV7kK+id6Bz8/XJ
xJfpGlouE1DZA09ljrzgY4F6Vv2wjPKTHmFllohlka6oQEc51EWcptGLr8QjgqMy
ufd+ZCgcCpbDGIb6G9Pr1OgSgIsagEocCgRHjA58t9YdwNjHLl/+YX798mDQVZgh
qRX62JzQs3MjB1b32SRpncK5AB4LKDtXuAy8LeLhNjtGvQMT2RL8i/6WJeBfQASd
7JzEC+OdUrab2COm69fB3z60gJ5AglHwuNnNDBMOYuic+C6AiiAbc8FsTVcXimlb
CdeavRpB76xHVyDFt0jRr8THuYZGdueMDZvSRjwTkqbsZiUgyT1uD5PaQ64P0s0z
Ez6Sp26rYHrT5NX/NLSDZDJgMYbPCuSDbixJbXZlzb6eScc70mI6WJFjFbbTH8mK
WOUt0KaFm72RHcbX5mq7ytOSVhpWYAT4yUcXYozth6cXzQ6dfN+YpGmhXdzgVnEU
q5OglXjGT86PQgGuG38hEJwt6mR3BLTzZ0zSg+ORvN7dI+CSWB/kTPFRyW2lcGEp
7tslGUSQwsVTpX2aPAOdVMUue18gY3w9siYo0C7vipIBo5EAXvAq3J+YX0yWrcMC
An/yw98iUu+VaMg8HX25CN+yTdLdtZVJopa9h8o/TOXJscMYtsrYgIm8bZE/QpCW
dkrZLSyFIJqYG+r5bBD6gzEO0tda4BQ+5wJelDR7g/fj0NQc1HXfir2w1j4gpNJt
S906h8/3mPBV99xg/oWTj5RL2/8p0dpCkHqBzrrDnqwP8nikPfeNm6xZiocvN3V8
NjN676aNNcQrHvT2WmbvJt2s7umtAE+uvDdjRwmWm7rxUIh1t+5MW7NaK0oFgo2S
k9yMouLMTqu9FBGp2Q3U5S9uTQaB/d1dEdcqRdwjcjYT88hKUD1BsvVMGEUfNPxw
M7SyCW9qQDhj3bFDTCZJJ/I0q4iotcATeJp3O+0X6vJMMqWUkl5Qt9pW0kbSZvqo
p7ttn1Xs57wnEtUb0wpWLJw30Z0My13bo4stFsEuiACgYWuobIcLoxT42JJLF5T1
xw56JOW3oZnB8Ags2iiYB8CwsM0LwbgOqpP7Q0ekgeP1XOsZKvWuqIDBsxUTSjxk
Hq+QltilBIfVB7XSjKU03ICfiieDe1QSGC2buaaY6BOGQctKnxTf+zq4d665vduw
lnyNmXm6wEGDauGifb9LaAwqhqhav0UyyF3JluVyhgSIzBP+Z60cFXm50twpZcpm
xblF6e2QG26ZsHvEJ6EPakYma6VGAlcYZ9/Dkj/AienFGY9w+5a486nrDwLfLv5u
nFTyBqfHmffS+eYvETgeWga2JhVU0yQw/D4zK4DFtcm5PJx/1RgZUayYzkwa6tO7
U2sxTlqhcOyEDJy2KhJEy+QWaKrmAI88SL6U+knea1FTzRqAsnFu+98TEP+IOAd/
7BZT58MsTrToalfrtAxtAsInKKNnngCvhgAa4EbiYTUtg9FiD0vlrYHrlQZKbELy
AUp7wjBS1WHSNEcJUDO+/TMhz9LBqLw5sPcYGfT0NxJTzNdog7GO62KtxR3OwId4
ivnXtspuCy9Drwx8paglmRiLe3aEJdJWt74J2jdJCKsLq8DUMGQSgj6NzUEcDfIW
kIOm96QuxahdX2Q6B055zENBut9heBpr21d23T/V8nB00q1OdmhBuXB9Crcy3wB4
/aprS3xUR1xNNZeHcKmad23OdQmJ4VckUmnbWoBnY5gWXh79pBeTQkBx8zTr8SM+
w0SOIFiAJxzTDPL/FsXYqm+BUwSEkDJ7/cnHVwuxmb+k3hnZr1YTzsQ5dqdCWp8A
6g/4K8XAbf3uF2JxzpzqKlxbagDTMyp7WLWyaMqAL1tiy6lXq97TauxBmVawbeI/
RA5c/rwCBymVBeEq66ezvDJ2VmSI1QCy84FmKpY+nMbAK3ATs2t/UkLDZO/wjRpa
rCY5qe2PPoYs4A4OHoFvKQnJ9uBK0D0yxYJptagXXjjwnk2ZMPognIlbbgWcfq9f
WD9RRt43wl/+tU2PQZQXXcZ8XH0p3mWLPlQWYWXaKTqbDgyz8SmM2fhYPwiiamlk
TzFrSrDT12LhhOUzqQvpEzqccudIjFXoeR1APSAUK71zNnGHgL2Q7Hko3lGFz0KJ
flMBGc4Um4lb7y5Nvx3Ix2L1nigxQoq9gTxXeHjqQMGovwtocdf86pGJmP9am3iv
AoiVj/YSVEgrX+ld3LmKVjH6DbLsG5YGWxmlN28+3UbZek5xCFFA9RYl7ygtAC7h
MoMZc2y1szeNYbGOlg7YOhdf5h60xu0jiAQKvcJtXNsZPfPWUZSLxjGJuLA1rTOE
uSV8OrwaYmjp1pRczMlgUcL9pYbXhSfTd7vEGUnec1XQPNbGFOWy9GV0iro0qU1j
m/edSTxOOP7pOJbAMSGrE9ZIcMN5+gBXOln+34qw4YFQDqh2AJBPIz7atgir6Puz
cNnsyF0OhkB0f3+eKznjbssPvWVttudRJHJczEJP8ZiQ6Xzm6aFuP/GIzV3QbJ9P
Gl3edeappl6YVHrWdEsWt3FFOfGQ26HwN+xh5QpTW63F5okgpCPL9K2MR45tsgbC
BtJMZ4qsgU1EZzZp2HUYE6JJJliuUtSwCqyiOyfZtbTvBrfT9fLLW24aSsEFIpBv
WH0hvOIqOOde7zq0wMS6HvIhQpG5bEfC3nsPSaKXuxLmhfRD09lA/jZ9v9/oYbmn
Ie9MTHhc5fvtyEIy1HYuNeuDvX5mMXtJrkzjTQrPki0ZglYA6jJig/B1yT6Tdwv1
vGjQ3K7+eciS73LKDFf4GIMLwcCK2cSCTd1bb9/+6UB+/xt4bgIARW7sE0H6PmLc
k5ViaYDVfePCPQAWPRabjJ4h52yYPNqe2QZXGqwWwwNDvamgGnZjk3PCzUchLvKs
KpnKpaao1JAt/GRg7d0Z6i0FHkT3xcWw/J0sOA9DoPs+JAi2isyBWDoTkwx1Renl
p7hTGvCMWoPPD/de6ahPNmPi65HKYRZcFSSEfkfMfl2rKLx5IBXv7Wp/GuYtWBI/
+uPlJSs9wLI2O7dtYwcXjLPK02QoZGknSpai2HIHZoAiEkwEa5R/AW7oyWNBxaoQ
3AnsfBQaqnQBYOOIaj16wOwVZjqC+MtCmiU07eqgYl6alc11tMOahXjoiRQFP+bN
8vqGt4vGig9B/iOWiWtp0DEBakeGV/OAlS0eDYRy7UiWMmA5bqJq1CCXpPTdZPWc
l8Mrvn4M7pKdcI8V8irwRQU0hq/ZBipxK0hcjrYBRqrxBO03lZck9oxBuFAasBCM
aTUJ8ClYD3yNN+ZIgNmMLI5fqGSfs5oKCVTiDw/2mDHSJOeXwg8uOIKyQWaV2JDP
+zYep/SqN6j71N7N437ifab+JJA4kRmh1362e+nqCHTqB3zAEOaNLAOwXpJMGxhZ
33dn5B3ay0Jgj4Et2eh73Xt9BP0uPoV6EYj8VOza7S69gEO+y35U2IFxhCEPlaaZ
E2aUJQTgTWITtdLL6mmohQckxI5YqdtmSXnuOGm2CCBAGuU9fq38P+VZ0uRNlK+M
VuwwCED8tvfxasMFTvvqRHwQgjbbb2lIOD+q/iw3Vcs3dH90nEG8/y84ToQOFkOi
tMPIkgeIPTTLyS/AK31Z6Q47Vtd8y2P98MQTER3PwWKVUEup1CPtwfJZBxhPMRYb
SVIV1qJ7UKKvGO8t3480YPCLzRgyLaMhMeFGU1TqUtkDvYAngf3Rd32CFFUQkYg9
9tX1fFcAruJio4T/yYZXlhuqVUnkIgX+tR4P9FOMI/YBd5ekUpn/OY50V3tNgcgb
ZyJuE/JffMEiaLKmFKbwEzGxbCXvvwDxnVafKLktFYNmSOVHzrHYRnV2cyNP5paF
rvDLr2VpQpzGQFHJEjipVvOB/bFF3e28Rc5n63SFUBMcsdnrHLzkTQtJRJUIPekq
S6VGmrMUS8emoAqb5GBkeGzRZ2KWn1JDaUWsAI1/zOY1QLAvlJLsCUFajyQAK0ta
4caKXp521B8pTDn17gbEzRACZ6LY4p7mQ25zVbs315hyNWaMesuMUyLbyvVtSMiw
OagQgmsAoDqDkJIaeZ/heLl2N9MJA/AO4Fo/5iMb8zMR2M3PYHhy81DtFiEi/F1i
WEsze65IC9sdNPyH80UeHtpVm4qRP9gWghzqnG28EUcj9+2pkYejAw+9JJ5kEjQp
nDWy2+YRzQwvwZcEIXgdxf9uK1tCT38Y3fe9ZF2JQzzgQSHl+QFazaEFIkYwr7/z
cFKEEN6UtxIJbcxWKQ0CfCDmNdhhegbHWItmErMYzsK47ognBMzRES+WFsMZKBT4
nkRnFNqntjyJtjYS8QgGi9WaIQGK3+GEJBMuUrC4OwuMkXA3hcs+iPCeF3a7rmb/
AY3xzm5krMabBFvB/gTw4X8eIvAxLwQwTMT4rAb/kIOFRM39PthmHhoYYOgEK9Xy
k4xevYiqxKKIKLt/VSdMSZZRakGRV+t68BI3cdioqvUFMriOjnLQWnVcp1bm+Rhd
Y2rcNYayTF1M/4F7L+UrGP/0OiOo5/NaLO3rCzR8R5oQFEH6UbKJw8lihiFiNcBG
BG+u5nY9bJeYkP21k03OZnUEhfeid8UvIWgkB6RcNuG353Zv20aqtz80IhrZwLAK
9S9f9xv9mKF7TwMteoHb7we6UmAXt98DwSk4tQXlqFB63RGBduVrF3CsR1+t7xmF
oghbv49r/RreBVynvQYxKNnrjNG8nS7nTv9CtJFQOSK9siovfkVnfhdtBhfmw+m3
o5/UNHYKUD5goFzi+IA1qkSVOPr68pJ8M4XDLu9b2bSmi16jYi/FPW4u+PZsdKBM
r3NvVunod56kuQucns+m8GYkUFuxG9LyNHAEszlh/glmOwNAknct3AjK9xaCHWMs
3xWiNC+GGYHqRGcpe8HEFrDRV1DByl9U/QhVH1iVYRVVSLMn33xjarL3wvmxPTJE
7yZaBjoeDY+CCR201bWJkBGiORgUlptnD6fY5sL/7iCjDPb47UYiNz7zuMgD5SBU
V2bCeb0VvxPgeUX9UEPO9qMS9u0guWFD8WgkB2PY+6P/nNSJ/13+J4Vgt3fOrSz4
kDiytUiGBro6pY/kq7jN0ZuV+kF20NU6unZgFgK9JQrGq0xjsiCjnHXh93T0lsRX
jwqwjySsjZyLJKb+EpAQju/iJfiQvA5ZK43LcGUvgoWge5qynRhruFmkujkO/1An
+ZCuvD/BasFB4IyPCEcEeuCBH5a/hWY2608192BVsQoUlYc8koShFvDkz+prgsKm
7mAkqY/XbCjmNFt1zCF0mIrbTS7jlowZXNerAvkyEwL/lQOP09MXxtUlD6M4j3uj
nkWFiqmlr4ACWSKIBSh1BsD771d9ctj0unN0tXedrMRTwG4T8zSbWSRzZUEBJ8BL
JOGcZxM/yIRTF/YWCIu2jJbqziT5skudT7NkkabKXJ+EsIKq/nBL6oRpwSE4qiU1
5wtOnbbwfoKRelWrIiCYN6EB/caJD/jI9Y2AdWrH8uUmbxy+vSVL1k1UBuoMS+gz
Jwd3ZqgBNpx2kq1E3SVwZOVGpBGs893UmBAliPE+LwqsqatRXMwF0Ckth0cZBVO0
Hd0ZZ5OHO6mcaFz8YORDOQUULgAHcR2KJ+j+QZ/6jcrg6ic2a33zSGnGe7kpZF49
WWwvx5w5KTRiPKshcyemg4+Vohhu2P0vrRjI+NSM4YiPzJkfb0MiLY+cLWCAENYr
tfcpwI80WV7/ceaMhQd1yzHTKReKBJhwWevQ38O8Z7EocRaTWMpiOLwgEbUlYHwS
wTJOPCPqJLv31TjvruRRJ8V/aXXG7/jDCdR9OGWJsNyzB4vye9KSiC09e30AX0dW
g8I4/FIpQ11JFwnlfqN62b38BdAo/IFOqGfN01xd7K+HOpnFK9C7Lo9ceddT8k2L
Eg1B9Z1QkWlkWwOPYuyKXTaMB17WsbTLMybQjrdKjA57CuHCqi5ZdaPFjp6lcdtG
HBI7ZD67MdBgWP4ofiEit8VzBToERV+zeQbk9YbbOf2i3mgRjocPzU7U0WCTBriY
8lbTZYL1Zd2KT84yuO+J7pBk/6kz2Za/jrIwo6g7X/ulwKV5bTpdvbiNIwagVujv
w48usFmOpjC4WAjwQ+L6plBQy1zYsbAEwgViwJ+itGOavdrw4qcweiEynM5HQy67
gzNLZed1knWgBsEgpfrNCtqUxQHrMI07602o5TcyQL0HTpM2J35zKjbnzHzJqSwq
jJrjQjtSCIIWoTbiLjj9/pfUNPYoc+SniKHv9ZSMcMaFs1+ura0NZMTGdLVV28NT
taxHSQPXff3xCaNyNpAxiwiibb5QJN+k/XrHs8FQklMyPW7Zp76Fi/YZ/HhJBVYv
x9gzjQcqssrFcalwESQHcUsQ798AyVXpQVlyO+upuxzUrjXLT+FVFXjB62xXDKKm
ECXfgA6qVEgsJkRXBTbbxa5oPq+i1fec44F5+ywzIqyPbu02+5CECaPREOgn7eO4
zSbkpukjSFX5Cfeho6WKeCfUns2jzPMnwm1KIKZDzpgxzqksy37rsVc4wM+FTiqy
idgV6Ye1TyWyCXm/jLx+hJIyAQKEhLbcjKkNTsOnxSMdAXE5AcbOGaLCn9zUftII
eUWYTUbI5EHWnOxcdvXJZ3BimByU98N9jP5r3X0kw0J1w54zn2P1KmncJVmLA3um
MexCNhGclypuolJqcYF0hD5qCXNV+liXECq3gPTJ3HQSY+uZQml036A4GlyUP6Ws
d11DnrARvGWoRRgPRdqaOaFQ1CEVGKszdCjVf87+BcV840ipCah9z8N/pzPqYO13
AKoHPB3NbLu6tW3ls3pG6GwPVp9Oqjsp7THScT1SAv1K5euQS1XzXnaspnTDW4iI
h3030vpqVko9z0m625J1/Tf2562lZX+C8AHQCnaxPKAGIHLRf/VAKSqEXEG+YBGQ
Oq3KtiTJ1jO7BnMnKbDdqflRYmLX2rjR08DocQPjNYiUOQQQvGbqf5gMLZB+6XEB
ychUeqJs494p+10f+x4uKwOm8G8ZbEyKlQLBlZXsKA65nwuHbSdREWL3CvOS91oi
pGQOjVrari12XJZhuM6X/6BBl7PaB3tMvaU0Q7NxoTcvNzS6M8ieDpaq+a6uZfk6
uxICiaozk79qgFaP2KQfajKmuM46KZzJnPqcWNAnAGuxKxfl2aT2r9C6ugKJUVpl
0myLhdtchJoE4sZkalzSgt1IsDREg1gS74kP8IHX0YHP/IJt7tnARrTaaqhRwAqN
cx4r2ef/xC44eY59NcXr/zKV3YFYfUka8ZL6mME/KFKw0Tb4UJQPiO6NUEdI18J2
tO2gxdKabIrq/Z9V75T4K7A8M4O43S2ExkXQOsdwHRRnEi5v9ZE/LA4bfOIjzLRb
Wgwut8ydtrobUCzRpeCn4Jq+znLXZHCG2fOaLjqxSU3TVtzCMssGfGjJw2r/13oo
88ztZELMMG431vH5cucU7haFnGbQTmZjmYk06A1tRazmDIEIfVVxRgd6IYcvWNX3
CfPxk32mZoHKcMnbs9JE2jfSgOaysU+NeKueVVDiZONqt+kYu/ihh5F3JQwUWFPg
9njiJLSdibAlNvZdTC0v6/M3OsywvGRBJfvVj9P4/8E3J5y14gRp4dzFAsu4ghFF
hV99Hfx6ZT4I85rWO9rIEHP8Dlm8j4gvIefts1JBaQxl7PqwSklcKqv2QEmPcdMc
khLan5W5grahCFNZQh8WhF5s3xpKbRQ6yMiYhGcqiqlqQxsL6/o+0o+5i93PTXCG
BP+YzXNXob5ij7L98okbz0aSw7fwN0yYqUUQCcm/hfgsEBC6D+hz55MGkynNeN5+
muFpx/MWiv6wtrkAnyS416HnFVZ4tu6YklHAWyXFAJ+BzAbUMT9hjsyf9jB2f13D
Q58pZ2NhcgFsRxYLB/UlWtom0x0chp29kAMwGVnFOm4FtorZPLJe3KOcUGzOhCbi
/XEx3pPYfhRgQ4VWhSxxjG0wekkQkMrybpc9bto+2Kie2BNzXCRYL1bLa6ZtOPLl
6yt5KYZ/i3sA+2E8OhmH/q2BeDuK/j1sAKbGQA8Ed5AVhs5vFuGTsnQhz5jIc7PM
Y05m6UbSp6mFXyXu36g6jnx2yRb2PmZK1NKU1AMoOBUt5Kk8EIfCSN8P5F7kGWKc
gr8fj7gTlJJGQ6JlHPyldjRoheEHN0PrTIW+t3xs0nPVy84MrrYIjZbPXhCwSMJA
r3SE6tw0q0Hhuj+58z/eB9mYRUPLkiZZGnj+VBH+O6mngvI0D4cHrOutpiY8e0Zu
DXU017a9Yw9xCllyRIQXsldH7weYANqpGxuDmTx6zTUQfiXplYGYgov9zf1xtg9Z
avUN4PT3SVI8gm+IVwE2ZACJ4yNYfTzp6UN3LvjqorFnY+1+1kOUejkjeHe5R0/J
c3i3De+UaJnnFdS3aCqNbvH99WWkDSyYh9u6qU67sYHCOKYgY/z+/dNJx4dTnbZw
w1+m/K3GYUlDJ7rVSHkMKe6Q9hSOaLLy9NAeSa4VG9Ispeyza+lqK5EUAvNT+a8N
e2H6/1L08eHsS+B0FzQNeQvBKgGXvmfUvlrQavqpk5LmNajCzYnKfB5aK75gRIrr
twJYC6kgH4FkXa3aX+QBlUohNyEMQlrDl9DOZZE8HGNK6E7NZHmq3E6XlI01XcZy
P7nnH5o4Tfo0wc3VyP3J6Bp5TodyvfT2JvBWlqI2mUbjKLD8bEe7xpQpBhJWH83p
DeugWKvKPh3kl3orvz4+WDNBZ7BnMJaJA+Tn45Coi/dresm4mDXWSwO436Wkwxyn
ghIv2gcIGkE7f5zjNW5OnEXK8JO70qpkJJM2CBLvMNkCRYtHKNJffDh2jCMwOBHE
xipduNzvFTkvO7Ze20mA754NuecL5qfDra+S47pNRtxP/ytV+rPSydTKtOA5y+CB
C+aZG36Ue4KOCkhOGdgMbm6VQj/GmPM9AqTWa2MubUhl9o3Ty9AJBRbTxkQue3oj
NqJvJEKppG5FtzbsG3sfsd5SaNfNghJXtWwP2TWqduIJasGXKwoaKBvAapMYOScu
NSsJIijVUnWwxDBHQfaCY9SZJzmPSuogRGpp50qD3p1jGQ/BAwi5Az1J6a+Yf+f0
+jEB5fcmdEZWvGySkdly2vP4dzahnFmHWwYT8HJhEbfaGKNb0+fT0PQyCRCO29Pr
r5Pz7IO7dxEQRrYB1ZzeO8TlldjZCaRj8OJb9uYK/GNXpSsd1nqbAQXb91c5TT6i
AN6HW1i41PyCd7XvMvBqnaZNfICelNY2T1mDKJosCaXw0JPJ2XR+N977aKP2gAce
+7nhjiEAViK/W+qILrgQHkrFxHB6RFZJwe8zwtacB7wMVIaMEnh0fKbn86++ZMR5
jwMfbXDOhl8mMG9vkelW1I0vvayH2ldHSmkHs4n3p0EvZKMdCBeJKLmF3JZr8+kG
7u8B8HwXkHxPvBcqWKxnSflYDL9DPiFvCm1UVT2AG9sv2mkOcT8Ux8aYL6i3iAD1
nATlg0ek/EvOnTPTKhEmnE28XgOhtUdXfSxwfMq+kZwudv25DqYi8kTV/e331JWA
AOhYt+3lhM8wfZINjKxs7x+QXoMjtELT1YzDA+HFJCy0aiWxnaPld2hI8OjVd72s
xI9QFYxZm7iuaE5lCqwZX0wojlrMKkKCuK2yuPc8HJvOtTePH7ONdpANLN0z991d
rQew91iIlQ7Eqjab5x/qDTCOff4EoT/x3/j1WTn5lLAV034cdHcaS0ymmizAF5dJ
aOfIioOPenvg+AP6TLi7znrVq6jTB9pVuIMThhUHdWFSYZBIQMApaOOcxlQ/aFsq
NidOKJhM6cCXqpcivXoV1qzzLfP4yCFxYZCp9rXISUAQYdVDtmmoBswWgqTcLXav
TbXTUZl0KEJHgcD43ywQx/gysvcMgW3+Hlyy9evPmJ3lYrp8rzFERwGaOwsLEtid
OMx3TRPsbZmAnOwMVVoVNakwEoxCe5ymQpJdk+GVjjqhWOZJq3ukEqdIyQwyr9u1
dyTQJwB5bU5U86xc9/H4TPvKyB2GNEaqS4I/PBJwRBxKcARfV/js7Gf50ilo/oDm
YHxHoSUUrF7rAvOLRMd2FUxqcS72BDnBSN//GX5txZfMyTV2ABikmkvyNb3/H1zz
uRmzR3xaTvE+QJ6Ql68a3vlJyy8jr65YF907cIOqEUM8nKTcbHonM2L4dpbkqyFY
r6tFM44JhZhlmjC/OaMQyowEv+FCIz6tgm+t7KupyPjU5gDXalfSZPOhkyFiaNMX
7vTFciTXvrqdYlr4DoRSKF76LYvs9A0rI8M/1S3U71bTCSWqboG7j+o2tcr6cs2E
zDqshsSpWn4UwhBrUfOttP44GWhBeH/vITVcfzIsgI6AHl8L8DBw9KnvnKLisxT3
q5gjYwJ36VbDn5dmSAVk65vK4soWUcL58t2CDpe737d6Z7YMVOTSt0IwU5qV0Hz8
h4039zZCUWVsvLZ57JXDoS58ufTZKg9UgPsIe1y7QG2qHcm8KnfjsolBDCW76VtG
0IVgJsuQvlyu4NvNUEefdGIaJfDfApS/GDGXKeg6EPRvUfaAiQb5SsjkgBohRWG/
PrWUEIsaSNsCOMJIVeQnErjGbMxAPHYx0KNAA2rNPOgcGEQRqcrAUtDVBWaYR/xW
QYdXDcjYeeTvoCV8V2sb+J78PheaDSMybvFA1pJTNMzWzcf8z7dTUCIfc5giTRfQ
hKIlWfGjuT2NU2ZpXsbWZFcvFdnDLdjdnnKDM7SuLXTqGRyIucGbUGbyxGm0L7M+
IYpTQ4+E5uecQHTLDAsTykKGNLXV/uXN/NPU9y7f13U7MX5ZHlzmRdcAQAybLXDt
3dYUd8ITvZUZ1F34WBCU7xZIZ6DKUxMX+LhbxYoxN6GGs/lwE7RaFuko3neIiEQ5
9YgHABQxYcXnmXQEeLBiiXLIRfkhShjXdAaugwclvgGRaadSbOImAfU2PoMBa3OA
KwE+ol0CVmJwFJiITCJqfA2lM+qcxkL5DybqDfzJUqFrKa1+pbPGZ36frODTd8tF
r6FqEJj+p5smUd9jdjO633HhmZ4JczOukv+xFCvMdesPU48WIM+LhNb6DkfZl5U8
R5e765Muzee2JnFICFFteMC6chEx9oPT0K03UUNYeYBsFrN03VJUNWoK/UxPE0Jl
TPRel86FyQEc4YDvtgwrLqZrXx67ONXGBTzm6FMsw71KpQIPlwve/SCe1cfNAxGx
peAAk9DNtTaEb+DCOQdX59NuGBfIXBI644TJYkS5suCP6KYDGdTHMX+wjBTHNe7l
qwi2ArU1HbtbTjnifuIis+gXvdSo7I5mLM5PZgtI+Epvhs06TCMiX1W3MIhvY4d4
fFvecZuSsiBNwh6X+HaXP+wknUGL3Hvp73SBmOuUjwLIC1JJHVEy4FLMopqR5A73
ie0lAJUTxJbOlMi/weuDr+th5gYwfwM0vw+WtwX7+6jOlDhFm/tSGKSKReHYsAV6
hvtwABXx7rMfhgP5NaYzZOOw6b8px4h8nlJ5BlJBqHb8sBA8UMImviMChxcJvBaN
NKc6PJF8ghkYS0DR6kDmW6C85UBEX1LRkjTf8ehLZ+lpduAqF3KdoURGJmDHOLIG
Tv3R6RyAfpPpan0qAavVyXTCwy4kWBQh0aUGPcrLr8yU/KuohLNYcoF2HGSMCbG4
bC5sRTtXBA46vJiIFT7TfczaiIJJOfMKTsVSfyQiKx4NCCz1KjSiqMzv5i7xZcNZ
CBSom5RSjSrHTSJ1nWpsR/O2wGiMyitau2W0rIGvJc2JBtzVWgfpmrpSiuySdy7Y
dKVrV2K5HG2MVShlDBf6BrBcZyn3tRlomWxZ/nCkoxtF8i2SkCySEPzSwXeIugbr
TVSk+OJyAefQ2fl+Z9efAyGToFOzFPt9heuKhxCxVszQQ51wzj/6ZnYwGN+F39ag
Jn/Oeh1OLKgPigiMnaUYT7wGF/e3dDAoI6h8YO4Myv9+h302NUVV3Mn9saQgZg85
uPavWaQ4rtCx7eJVKb4ci+vH7GpKkcoUp2TMKXPdr4HQHmt3iPKxiNVNAPIWDKIs
LFQMnw6xl5lb22fJyGCAW3g1gNzGgpcYjdzYyMhMMoYvVEhlky/sk04RPhVS35sy
YzVXiKqSJu8LEfygj760LOW1egeB0RuHDCsmyfhN5RYFRDw63ry+tZ/mjLBeIMeJ
idoDVyiHyaOshFIKXRQlJKA+5NUm+6lOMl5Zsma89wKuVoFvoW76nYMMuV9A/My5
ke4wFDKzcZe8QajF11YPoBVIFjyliupDDco0uDWslltFB0PtHRUZNCNvlzI7oPlB
5kM0s+pLEnLWAmAarBvWF6hbDruzw3Yey7lTgQuBejc9Rem7CZbEbTzpWnSpbfwA
5vd5zOuCYYfNW7ywX/+eXdk39/ZALAbrLJTsFVZI3judwfTpPC1HXHVlfi+GnG7I
AeIXPYLeBPz6Lptet9wQfJCOOrZ+gKvqqzC7k3WauyHeJ5C1Bg9KhN0fAV78kdDt
Gm4ymCkFBwv+R8viIIshXE5uzUUS8PEbYApCKyBYA9gdOhZ+vekXyedDZ7E88Tsk
KOJ+cZP/ZzEfDkcEVXnTEhGRFtshoLphcoDoBETWhfHr6XxmCu2VUcYAnPazJpsO
BuUOOFe0HCKOnGiLWLZGApZUa7doD0r3KDRDwTqfbyGZBVJj3L4p3UmMwke6grx/
77kopoDlZOG5eav9GW+ieGDn+m9CjzNIMnC+gJW4GtC2Co4riZ4kEPawIW70EDbx
2zmIMWktCp3AtBjL8SijLUjSTbWOc00d+ra5DXppRsjgMMQhWJWfUSowglY7EmmH
yZ6oysZ7pWwsYekcyZllPax7dl6mOW7fveczLkasaHUSyexkRqOi5G/mf69v9Yln
XFCAg/ap0Qc5KJyaoW1grIgAHecn33gJRnIdn346RGl+ZLKKJxzEKoJqmZ13y0ex
h9y85CKh6amC+nicKoc5QZSGVL9RJ43J0o5zFL7ftlKl7EH5WHVL0zjZtVgynMNB
ci+lq3Hoy4bbPaLtq9Jbmt9NjyjeC+dTnf5KizKpnQDoBOx8CeyNar8YUsvMzhJq
8SrWfmQImv8oxJ5rzYwNCe1WGb+7+uhV0ctnJEVMiIXeCQLqHIcD8Rf2mSidMz2a
1vd4wn3X0Lf1SBK8e159NXQP1Mxx9EUSW17G59wrXtb2Q8NxhnPl/6zgudHac0iA
8B9hwr4CmtlWtBm7iBdBCND/tJVEiCZsbgx4elJYpl/ELahT6Mo2rFNNcWoJ8i/f
v2eux4engotfjZL2x61FKZ0LKRdnOc1tcFIVpcghkY7Kxp/Yuogu8RhWMcxy1L/w
mXabjAG1B/G3Wbl4mHoPtpg74SH6i+7CxtHqfytlMVxsvw+SEoYQNrVDbTmpEjYA
0Wi4ZPfqMYIPxnp+FmBkiI3aKrPF2Kp8azkKaXfib+oddWN1yIkg0Pi7rtBoB9cj
G5rx2rFQlGMlQy9ejAc+CHuXMYmPTcouCZDlnXaBMJGS9B43LiV4yBZb7N8mfZKt
39Y1IWBgqj/jAwrGTodTyFbft14WwICfsdUMaRiQF+OGcBL+LTphBTrgyk/IQXqG
cppXa/Cd2t4s4czaAMiXouyJkX7auDabC6nqTnMTTfk+fPqL4bTCVWDAOiSDQG4E
iuPwaNk+Qq+NaSvEullOgd0QZKGzwFL5mE39K1lXEX8myEqg3M6kVHkDBN5jt4/p
/sYeRrbXpxDYE7vmU64ntD8P9GtKvp7LHPS5QRpUl7EsBg/sN2qrscqf98AYMs64
OAMAxDnnEqVJzD5gZStMqhEkbvMeTRglz+KDTdsQynKJMQye5DGkPrs4n0rGEhWM
mdvTgUq3HOPMb+LxjVgFbjmDsDuFPs1r3jvGokdKEvjANBh8DKkfwR9GnNpSj6at
maEKkwhEDOTyQY09QJyPBUAcFSYAgz1kxV3qxUgmoftqGo4+RqKJSyISTYNat1UH
hSxtNoGaS+ZQHfYsh++pai3yeRQeTH1GCXPHA8Y45AcTxg0uWRRwVV8ZdvncHLoh
niBZt0/VZnoBAUAd8sjpetPwfGFYpDF6aLHmT/TQ9k2guhtV3wT1NL3l09TIxb0A
2mPPOMp3HyZspQbAS8WIB8Ei9Da0eDJxn65zVNRAvuQwk+y4uY2YDEa/RJa9RuB0
WMg4So34r2znPg2EZzUzEoPrLmFumKTG8SOJi5NbE1YEA4+6JEC8yhhU/cRbXeIU
M/sivvYiLSknc1w+QtGnQAjmAnYRk7yBtGBu2vfRQ4qnYnOT/weKLk7JVN5VGQrJ
xb/kl9bB4YRaLj0nQxXv3lpQ4K77HAtzbk0zwxaj2P1ORUK9BbD4FBbmPy2LMCM0
CYvSjsA/jB6WUXrfAUYdIzgdUAFLqhU7UPoFRVo11M6eMbPD1f6prVbZvyP7DyDv
R+ryOiCE5KAiQ9aoSIjmkyUyBxxRU4rnSD22PcVrzAzLCDG/urEieByWYLGkaJ0e
faNacOWCaMCtahsPBarznjKIBY1UUUOrR2wz6/RZ52+Kpf7SfPHAQJbWdKYgOkIi
IcFHcuXTFaqIiC4kmLVVFOGU4kp62Dw8Z0f07/PKT2GmC37GExC39FzjT+Qd6190
Lg6Wcl52hErUPWRWc9l1wk9m6AEYdETID5b2BStl5ppxyd+7Dh3FyeBmZ5a6BnIj
iQ+Rxb62AXrg4oPLQoew3/jyvNts/stV5/Cht0ANU4HAuen//LZQNZSgYTUIsnKT
6EKiKW7Vv2BlLIJTnalaBidxG9p83fIAQAY+Rld+6k/jj5p3K/0v/9o4RK5pPbjK
/cSZsx1Bn0xoEqD0do2iDnCZP8utQ6ojn5HGicLX212P6I16aLZZGlDYn9vEg1NF
yO+Y+zOTv5UcjbAcouqJiEgPhn4DmAsRZMDpBcfbSbZjWX6fqeyfIePSLLxaDlvp
Q5tznqaQql3KOBHV9kFy5S15q1pKldLmdlEZa/JDhYUU4E3gJ4NHfJWgFoVpPSg8
OkSDzSNtkLGH04yQtPMZzdOmcQJrRDJUEmV15LE+ouUiyBtbqEGcNn4L/bvZ9EHP
cw84WdaKEdOzd30g5Yca+yhnlpzLW0qYYjWYbsG/x5a5Szh8q52iXFseV8fflHlz
Rl57/wCdWstH4NWmIQIcGALRyaIfOM/WOV5ZkZbQQh/aNZQh6urOyZsSN4Iklh/7
mTVY2vr7Mh9mvPqfHFkzRnQJ5qW0bRM2ezX2iX94MmsyTuaU7d6A08QjFvmNXpgF
Ix4VHxH22w7DDahEBznERuuC97crNnmoSK5aQLFMhulay9h8XI5JSWpRFvgTJZrt
nzhiOpC51dYjUnr81p/UjN/g5m1RklqrCG5ye6zLpW3lXFFEFV4k4RO8W2dKlEZz
PPEZkhfSWZ4kQDv4Vpq54xEonwak4eCIeFZLtVGMciwGSEGyOcRFl1UeTeGM1HLb
Kti0YdjXQIdB+2wC3St5AoW1ZyIGfIXS83LeRpap00KCPWVQH0teabsePvwdNkX2
K9j5wJ6lnlUjKt6uuzOcwkkhafpHjKMUbh3Lj8XM1+7LtB0zLF5I2kbKfBlQ0VKk
ZV3unst+MmSjWnSBDH+dIIyy27AktO9ki/aTeReOpAUBOalP8o2K+mC61Lye8Af7
4mmB9lLm6kOyxLng5+8Lr7fRgKFa3BrZf8TmN27LTldA17dMNpHxusKfbpx1apn3
BWa/h/y8B0/8d39ytnv4SsQxGVObVRLbF2uTeWu5seQwMEjMfS7R+rMkSVPjQkEL
GalQ8TmWkFHyf+4dKpEJGeyMwTO67C83heRBdZxVUVxGrIpHX6lCBFNIlRmQaAdM
UfIUqWabRxsaVay+aRh03JZlD69BdKsWw7aEeOvY2ftuTA67ylx9fdP8PAYbokVE
ddcpM/4TDnEZpuK6pxtcfUXMvZMOY13NEbnHAfx99px/HJsO3mslVrMSSAeNgvfA
H6A0zDStLtg9BQBw+zsXzK8mFfmrFHnuk9Teox9OWu6eIKU2ZLnH44siidZ+cUvK
Txg+mrvWT9pnbTw28mwtD9rLHOUvEIHNGboW67bpeeCzIwOu/ZgQ3wm0FTb3kBbl
ZhvbS+DcFznhT+vbNKKB8XsEjSqy9Qq9KEOaMPpwge6IMuc3TuXTixJLOIelSqXU
vpyaAugY16qgGpo4PkMuN9LJRla6N1V5ZLzg2s3fCpW89nas4UG2jR21zJKi6odP
g/S/P8VVeR6HDZlENXYMH+2+Lqgs9ZjOYv+N1WWfRP6kMeLDmL01N0jo/S1mAkei
nf7wXKtGyTyRZHeSosvOWmpkWO5SdNIb78TTY/HVkbZk12UQV0q4I3lEsXeYpA/b
q2QpJ/PMzBXMCcxRWFsQ+7QETbyUtzL67lxigAIPaF6Q/tK3+qExzWXGgKGfzRHd
EkUP8dwwL4zyih4a0dcZc8MLcnzlg9rWD2tuXXV+f2jSfAv4N1LxPqXCUflKaFrI
uPtjppgAr0bGLhyZNYkh4ypKN8509cg8krOfOvgvvlYkg4n0O11MosTrOXWr4MWM
gFRBZk2ZoytDuiI0is8oK1VTqa1jrpHhIWFTn37qA9HEs4WK55ehYBZVoVgeyZMa
kdiQ30l0lZTcyR6NzZeLNaYqPLnIsF6AaSN6YaAyerjlbU+49QMDBpb1Ulxc8nS5
2tkHjEPmXI9pLYA1l7vB6eCwdb1/ivdlHFn0wA0r33n1YMYCHt/v0PJfEZ5rML3J
pABHBRTiSc4cqEY0+SR5nMcYcmf19urd0CCYgCEEfX+Za2x1Uh3egHF/y1zIR6Tg
rH+bKQqjvCQ3ppM1YPq96iAi6p9fZ4bWj1euAEFU618YxJEb8E5vyGEfSS52iseM
trphf+kRNk4wO0eP94DdT7gWS/UgPKKlvFooNnsFSD05mA6olvtoaKrsToXvP19Q
qZsyi0wt9N5WiJGzMkCdG2bY6MCsI2Xx1jgrjPE9zwrPT6V7mg5xNbCshXiaEw7T
d8NG31hz6QTSW/Twb5XLdUoCDY54sd9G73Ig3d/zi2Ac8KrDowKVmuyAnIiq8HqI
rZ3T1vqBwkj0+KJuMboU7HbV3MasJoECDPGkhuHwXkJ7wuQMfNQ22TcQWlM1rl1b
DG+PRQ0yB3vPxIvWeDyAr/8JPjzDDCkSZu37Imsr+Vg63tZFAlqUEaO/sgIh6ny+
I+w1PKDVA0vHlexpBrgU3THzXrq+Xvzxn+09B2p1NN9loFkNGhdn7VulRpAUOjQs
VdjeuIswZkgfB2o9a/iZf5335eGjNZ808cbFRGaTl9NZxcZ0EcE86C6OmwFwaHg/
ffxfnxtqMAu9bio7lpz2uSLHKhDPMF3eOfbnTj8ftSvHbtNNNxH6uk58wiZ9zTdS
CEWZqwrg+TWnL7ofTjIA93E315ZM5G0/CMfHNXuwTHejdDW4Y59MaU06AQ0c0/me
ICv6rFItC17S9dGVQHFHG7PZNLXMOIuCHIb85k62UQevvjW7GPV7jj+9jnrPSIDp
9HgNBe668FCSLiCdNfbKN5WPYmyEvbY7Cs5E99Ph8fRH0lB5dmwYKKZyWf+Lp+wm
/j3WdC2V9CSfYgpCz2iMHbUf1ehYGdbsxGsBp88G2Yc6QO9A94qzW/FKHf0K5UFq
+KwcD4319CU0OyCXwc7a0/HYAEwlOoC1YjVttBluPem7A/zKjaIMIM7KFCzquyi+
J8ZIoR/AmbLUnprfmb/Segny+hZlxzvL33v8ZbKokAytaTqpT6fwjv+02dIL+Iox
brB8QyViLlZoRY36qjNSO0nOdV5bXlTVZp1blDNZqW7IjiZi8GmWgYiZDj9sSgOt
Db1nDgkUmBpLck5sUkgqfo4jyjcuGeuLJdG8TqNrt4MaMfK3Bxt8RrYo8dgAu2Jm
kCbzbkVXOMvMesTwsNjFUMgAcOAfw8rta6S3Jdz26/PNdn7YEt9n3a5RPh3AaV3t
cBy0PR12yFu+B1j8NgVopJF5H8WcSe/bPq9DwSgmitGWeImmDgPswRrCKZcM/Xkm
S6LkKfKP+rA3dBOufZoqHeO4Hg13ZjUtPqYAB8g59BbLr8BXg4NL0kNMrag1vjvT
TxZf2bYhBIPmC0EGt3dRj0paiQp23UzwOf07XR/C7YO9P7oII2GlvsgWmPA1ZbRy
sgtQQrADxknrUrCw1oyDVHggwjuzQFRuu3+JfuNhSHMzGb8zWjR6osPv3/dYpnf0
5Vv3iZGYRoBBotm5gFEh5y8B0P+2J5uWrIx5QD3wp5jv/SbpiB72vunVEnbO/uP1
GLJMKzkjX2fmvVR48wArigwc4qW/koXUsus6Z4uZDBqTHGjvcRz79UF8feNjgi0K
/G9/7T7HhNdiNR0wsS2Mh6J2ci4lMg4ODtUikTE+hQcD/7lRODih8iBBIqTxU3ak
dV64IkoLWTglFG8R1sw/MyhhiMYvZ8p8FTb8wyRTCSbJQkz/Nr94uVgH+NRV30AH
vtbf3tlzUpo4B6NTcueeJIN2WYWptRw1aQeOiGF+OktYFpgjRwCg60Ey34t7qgMN
XfR0oz+udtSodWqYlCzfMKE/suGBV4aNcbhfmI19CA7GDtiAGXV1tdn9AAAACSlU
SHnXD3wwk+oakjm5Oa2KExSvoed5pWRSc/0Om+uPcrnIxDtaD9ywmhaC5Nf6CSN2
AAQ/+2fX3nfqu9jYd7Wqh3UeIBBsvpd9BAfFbkD9X8fsv/c3Gqk7+DSfm5E7jM1x
gl/Ar/ShMsYzIwMI1gs3t4t3Iyqy3HsNS7kNZoRFvLa2z79tKxbP82SP/63oV/6p
Z71Ltq4xMbh+XMR0wTK+5NzbyWs0Kw9CEJVgt2LvuldZxrikNhrxCGzvU7iBVYaU
DsM8xDmsuTF6qbVdTYRPld9hwWHB2iobE59vOiknSU7zQiRCxaCEcawJTEsjnelo
EodsBSLKVpYv7hd1nPUETASIVYAHpXlz9WuvSvXhuN8SzdYATmmGTtg02PoihqF3
Zbqnpe+xQyST2reYEf2rdt9zC92Ky9NNBtIOlQkAtr08QQAG7Dkttmu9INa5cMQm
rqNebJuJHtksBJr17CLT63S2AmuBbXZGRWEUY2BHYWNXkxW+qyBEi20erfu77q7t
oFDoOwoHAVVrHMclf6sPqzGbLMXjZrM1Q5ct884mJptC1cHv2c3cShU7kENhUyiy
QO2uMXJfcgOS71KWEckP6Mlm7GwzXp9g9TzSqd5/gJmb8U7Rsf76hOYJc8iRJSxC
nuvdB+dzctczRAaBuAIDef1aFTF5yntOlv/oJE4JpkmqJVYJh8hA63Cz+iLH/jdm
jNwANf8sK5N59iNMM3qq7imc4eTUSS6a/uud1mdguEdUDnAe/Tv/9GyUyG9lMDbq
srscuBb0TLzvb8Ks+hKcT+9gE+GqT14i4bc1YgRY6qYumOeePkR4eAqBPol2KpkF
trNL8ZS8AJKMWMswQ2bU1zDBgb9wFb0b/eN/N41PUQfuWkucIPp86Nzq2D6WxCzU
tfsdw0G+uAwHV3bplfvoRZR+4yuC8ASxssP5Ftfk1cAiskD7YVEYEtF0oeKufBNn
2SH2vaa6pTjoAPwUvb0fPNTSr26RUxDm8STg2kbaL+6hgP937VsqUQ4vkwXGMRSc
JRsmRUPBAu3iZg0fyscPvQzvyHABNTyqAmvHw/qZBRptR4N3upgfqBWZcgUVuF7/
/WOuzduSMTZ/YAc5flVREFsljXJdsdtK7NRE18EKOn9FLBn5bBw79pjrEK1uhSar
/HebVO2P4lPFdUVjEySaKL8Qyf4/0Zwmw+Pg7VqhfV9eQSiDyq4x9FiB4dytoOak
HdmuTCC+XP+nCa/qDmwEdSXiV/ZAxPf/QnENBsgTZVwROI9DtT3CgPeM0F4HhQh9
fL9qGAZ8i9owxGFbulgqkJ4ykgsBqPUBxZGMiFzVwCt3HyqWgCplW7zdihVBbJvA
rXpOGgNfcUR0KdOzSFVziKkartKXopV+URF4tvFXIS8SVfIgrwoKiJH/SnGU5RmD
lBP2/JF2syx/RcHURQXrC/z6cyf15ubFzpstAjN1zOZtNTo6KH4K534MMkfmKAdL
+J6Yy58xzDaBTFDOsQszcICZVlyHMegFsuUdwZKJUdKhdFoYAkUUfTF2uw6AAAd+
8bWsWNszhv9KsfQlwG6wF9rbRU+qF3khlCV4CAb6w69goZzyEaXCxOU8OWJvmP9a
fba3cTnOHJrYny2j6eJSN0MgmyQYpv2iq9ARE1jOb4NuEyOL5IdxaEUcLTtbKEVC
+EjhiM7sDmteFuaPsk23S4D3kavrcj0wH3VLHt3YlpYFp1bdMpGiLhv6F/d83Wtp
rEjF+NwBz578b/AlHUN6IbHIT4/7PSxGXUv7Pkcq3K3pEqBHpRENmbmm8bqk8EK2
WV577DcYeazRxCxi9JfYoBsxl7N/sFzUjWOOphxBkICtDayPOChRhAECoVt3gRll
9gNr9+bTAewVfOP3YuWLpl/xafoPiBTEqs7LMfMLHJmI+WWY68mDKcJ6cKr9GB5w
Lf5qxBIEYgmTY7PT95uNfKLsIOT21bPrVqHk4Scbp+C+FfjepjLQX2EQGmguJaBv
stc8xW7w5u5nRH73PXosU8QjCxzZhTFVIInP23ptm8k0P4AtWWnitLK2keEaFu0i
9nUH/DpL2gOgabqh1edngMFY9hl6gEJ6xAJfN+7knFzNuRNQGmfUNoawOg9cPxmy
MFdsfaKXnsGnhwmkx+8ybJvAMru+BZUtt/lPd1e2O6Qc/dIph4DaHlCCnCAOMChW
XBngZkSrC+OxYsgYoJ0UsoVz4jBy2AsGYPJMKJ7T9gw/eXqGdwkP+putbK33vOPR
ISzq0lFLWoNz/eVtxDNlNh7No/bQi40IMyplqqWxGMMw8PFn80g5dD6Ob9JaUJQf
xPa1FCEIRLRVzClfkkcze4naaiPgh3FhlKV2zg5RAK10NUNUsu3TZNy73mCBb3g+
vqPsxQ0+1Pg+j5z1n9+HuChnw2lUWywwPQQT/tP38jDD2uu5n+tZeFYFwSZvyK7z
7/GiZNPmMYs0SQmJEsZJxZiJSmsewHxiGiDAQZSeRL0bXXuM/BaIQtZg++LTFBtr
mZVq9xEqtFPVtIqLteEAPNn+4VVP59XTXtdjFJ6a7xvO1dEJiF/i4yXg9bSrJjCo
KxTActClFTmpgIPTmrumrRZfwkVcLV7Equbnfm1IIndNgoStEdnQkTO4jXCbUPO6
4P2Nx//brxGjYtxyjOoojlx6FQ8/ZM/1hoMah5AeaieInPLPFyCx0uuzfF0KU3V9
IhVtfrdU3nLO1mO6nJB/3UNAyIQ1OV5pa1gs04LzRgkF6ga0CBhEQrWUTexodQFB
K4MjPdhFdem9jXOT2qVWp3u4wMRxkfjJoeyT9LSI3m/Owgsn2u8palHSqi1WCBA/
yZ/03qK6mex+8qSDcCHk19PlJcCm1+hNbcqsBbY5ejc4iI6g/C/z+O2xNPNoP2z4
hoogjWro162+Gd3MCAHOGIWr1HeUlPb7aDeOBTHmFiWNiMb+eqeV91Q22hOuW9Jn
xAS9b2N2gNR2tBTU/uDmH18n94ecNKMELpFLBD9Idfz33K3T/gJUqmwHOe2pFgvt
wRrA8nQBUaFSTru1ayu+VfYAxOvfmgZy2LPLCcCYN129lQwDpY1rcAeCqMieAdkB
jf8g+dt9jLRrys/+tYG+Sy7QK7BgIcVwsNuLfIbC8ujeqhXa4c53RmIP3M+fSeTy
NqLpNdtWFY3QoasO12tou0daLfDK7xms13wxtub8YPx3UtKDTvt/fhnEoqXA5cY5
auhcLkgoUrx6vfoI4d31pMLoNXycpy5HcGClD2bsTj0P1D5WjXMRJiN23ZWscrPk
cW26tSFg8qhGBMBxu1LONafhOefKkEj+XP5DhAHWDbg84ke14n/1bJSVtvuHZaVb
K0ukSc99otIWM/TojfikmkD7axwZfczqGlR6Ao7uom3c9fXrxlZ0BEc+Nmk4glEJ
l5/jGmoaYGgsc754a29qQim4Jn9mkYqYaCae8FsYV9yxGuLt/Zo7y4olyl0zUt0N
S47aJa46cNOShV8hJBFgTX6SucEvCTHq8WGfdF/sePQwRQfiyHfIc673z7ExiqX7
y7eCk6+rtH30L3FTmBY/lktsj+00DZAQwG15h3dReBmQOwEann2bmTfR5Wx5IKBP
CCiZjIwMHcH0QdCuXGW8SOvdppDhTZvPuo4EbXUKmpKmBK8efYyOIAgdHrvaXB1m
uylbIh6Ttke1XXFZues9ibajBiPyWOlaNu245bui0pvss7JtLBasrCgFraV4Jxlo
U6jLclLOMLSLvOvay3TBt4pVTY1f028kOFJKVk3lLQpEY6gZR9fZ0QeatdmIVq2R
MEneLz8xkjuneYsVlxG1/EBwJGItJOAH1TCv3KAnmFkj6kr2Fe/H6TfVXOel6o90
mTyb1LoN27P8IxIowV9D45xC5aOnZ0uw43/35wOHbl5YgpDiqgV7zuhTxx7qF0zA
oHlN625Db8H5DrncTdzSFlvTe1qfuikV60LLzr+Yveur/cK+hFSYl8mNjYXhaMQl
XWAN4ppU4uePnharhbJ5aRxn1FO3wLFbfedNIteo8R9i38JQLr8eMAT69GxrqC6y
2sULmqZL0nZbaVmVlAjpEM2w3h4mCvKsRhVjK0d3CbYkoKLYg8+dS9kEs0V/NAXh
Tyeoka/GfbxCDt1klantnvn8sw8J2JJzWU3nyWCfe5u+vrYRbx4P7i2Tpjitg4VY
7FYh4Gfubn+eBFUZl8+3QONxc8GGFhjjNHhxr2z83q4n7n+Evklb/PGdYE/68aom
Vew934IyrWeXT0AN6C7cyx3V4W8Lq1+uAmm+0l7Us6vyFWWmLpf/27McrtSIch2Z
oPKeJp1LJ/nbPPIxux/aY5K/LHc1zUMYfoFRn6foxIV4osmwKnDE9TURprBuHRin
H37WswKunWCN2HJp2zdzcS2Q9GgfnYEfTSOOXqGGzTUTF6Kt55U2DYk3rFOe7Nwb
Mvrs6eIsT4EPAnQ21QDoz1OIYE1Tmcdmzkr9coObdkXzDJJg/e5+/dU9T+rtvUc6
zo6VF2Xq7P9v3xjLCgLCrdc6RFr4W3wQmeQ4D8nSzwIKAwhftoIXCk20uvb451aO
+Yan5E//2xqQtU730xur3OzpfCtwGWKy1duuMUMBBetccoYiKR/ftCOMI3cneLka
XmJsruJSKyp81sv2m0iz8fu877Odn/WRZwP9qrkH4i2eg/mWQ00PizldBl+RaXy2
84o1NScxgoRKTx/UMrAvjTqLqA0uJy8CoMaXpsJ8kCL0aVHLy2hMUV6aH/Dihh8V
T1yVqDiL8neSC9OKUKkTrQxrrcgUS8Xy90hxZOnUfwpPCAq0BlWFL5lcWEpIL3kP
E0JKdJJ2ci71F3fs33YqJ4beuW7mQSFrydGLsZ3dLN3SauSMwq0G2q1VamfAB25B
VwKCmwO8y3dV0Pc98H5w9YRcIJ9W6guyif+2+ezLhFtbweAJ411fkqk3jHNpt8nD
N77jQ7Ei7qQrjQoIiINEF4Yoi/H5KAK/N6YtytQHUucCZ+hbLrSCZxKBOctMZpLQ
K2IKmkFx3OxI1ypnakl+XXSTb/1PuAb5uwselgpL6TyXekNYZbjngwLMRyHCLzHu
V5iJa0lp3A1R+LCnxXWdIet3GHNnwyE4XpBG2g3GTDZL9U1iGsKrzMLh59Ukdgwx
CQJhSPjUe5u6PLd0g8eqyDwsprKAEGCzpeD1y8MftzUnYKS2Kppf9mTrkd8enHof
660LYqMKo+HrvUFFc3JjJGx9hKwuS8/+wmyu1GDawnrlGoPl4d4gng+AF+6BEi3O
t8VZehMa07TScAEl+5/K2tPi10ST7MMvd6gDDVq328qU6F73K8jcMJOpzHhRpMGf
ukYd8KVQM1YDcm7s0VKCHc6/Q5f1o04/SDKPKA37UuSGKY0KYWJt/WuFwud9tjYh
jKtZIzG6pUE6p9u9f3xSETGMj6RN4jXYHJHkQLB9o6JTosdc2f0WNCh3fAk7dLna
f43hX0jQ2H5xKCUTzBa2CIdbzMJdOhO5XUxlKM2cZk519ndmidGHMmq5oWmJdgWc
WNq1aB8LZ7dBlXwv9UyY5c57PyShOu1CsdhPYfsycj35LQDM7ih8tyTEZHiT9TMe
0VsRzpSb4Jx4JGkyt7TWQAQgjnmSZJekzuDsLNVNF9g7tL7QX9mSV9lh9iFr4osY
jgZbQRZu2bJH88ph6txrRjgjSCgcOvCY6VL9tU3E/VBtFrt7MmLFFhY5agUf9e2D
fKjgNSGJbiuJwdh0A7lFUOZjTHiR7ms/ubyX3LcwCU22aBY646ELBX8YKLDTgxyj
nDqkDW20Jyvl/iI2Kn06R4+3Ryo1T0zD0SOzSqRpzvnhSOKlQd2ZX3ZaB01/05Eg
5O0PKzVXdxoHVM6fhjDOKMdwgyRO2nKlDoUYG61YMbxBrPOlYPVT8/kV3ZBSo2oC
8Qx1p3iitkwoALMah+bmOD79QSmwvf0KbzfzPQKN8hgrD/1G7Owj4c0343oYemfI
UfP7qC1+9loZUEAASeCc2XRuXaS0Qua777b9hUQJU3uR2Z7+HaDZr67/shujsV66
0SpzbpuD73bc156TKBp80SQFvQrckUOYwUW2eO0fug5rcgSjxNfI0t+zCs1AJhLf
gf5Z6o4+5Af7Gq/oj2ChLBsASyoEJIbF6k2cbvamthnqpnpvvQSV3hLwLyxREVgC
zvPucAcTanKaJeDYT666n+2DzDjpSGx1p4YzpUrc330RIlo1fV0A9X59rvpAu+0c
4Br3yKJYbnNxUm+rWE5XVe7uQ47odhSFNlOjYRJDjW5q1LgZ2oINQnCp8RBN+D9k
ivaq71ihwZIO/jC8tSC8ootcwcjhKpYpc3otxx6/+5+CwaeV+3VOKP8ZyBsijlg8
4S51lzh/0PE9UFzWipwZKxxN8YJ/HHunZUMUF86pKfPcCuv0VdEVDdnRbqX4mPLH
a23hJWhEV7GfjC8yZVERzWiiUwNypTpZbPFq+HwPdpgz7okdFfqc3fQ/6M+OEeY4
tyjiK/lBEiz8Nd/605cHD/X8qY10HrCvu+7QGkFxNixU9bvDLBnDbLgWaDa4F9BV
M034I9iD9XSZZC36sFV00vGnCpWkbHhlCltOVNo+0pgzFIcbh0JrXLa5CXyw883v
l+7O1u98xpexet4BeDj23E0txWwdLPD0dnraK6yf9p1u4AhK2QQivdk8RYynWhPt
PQFXmb75i0gnNFVsn2Nn5+M94UE4KXx9CGnk6mZqT6ifN2K8jDCc0uHo/oAnKI/q
hhEPjdyxHrAHdIgJPVE7yR1PW8uvdQxqkErqT5V/AY73eBcSdithaCPkwnIhoBCt
53ns74RJwzY6xj9HNxNiDddEuLXxglzrpQqaDY1CmcofR7WseIr5zfPCTWccvlw9
XYeVCPrzyj6DdHUaj9/bphqzwXUfGtE7Mig+8UZUpeoQPxM9z0RqBUaTUfqiEffv
9eFE+800HvjbxsDUVGNokptpAf6OlMMXwen6WW21s7LN3n+PPSVIrvwun5LD1dZm
D4HNR81UReLRSAxDzbkbp5h1x+zqsiWqQs48WslspDrEFirEx6pKDtMinU8SIG/y
V5Vg4OuImFkYxQNZkpFfMGmxK4Wf97Ai7sgAlcAoVOeSYBjEXCGpE/2VjtrvIweu
XX9hUoTsPfdO62PNqzhoHQQrZb/LSntGTXMA47NnMdvas1OKPjJS9SE6GhB54rYr
OTpBzEmoUGkkqIC06Ta2ynAcNKp7F3VNC4SqNc66ah2KflUhgN306cfHJCKSo/GG
Mil0V9xOhnY1V7ZKHKAgokpiQuS+lEB4HiLpcjtDX8GTHkm6s/UbShwFvX1lmGfP
DF50J9p1eekIXr15gVfDYiRQ7pX3fABoKx9X/+Kwe9iQheW7LWiF3HlHHS10trUN
B7gRRtEiqFjshSJ3uLJPliPWv9RAhhCQEVZ/iq6o06CYBbjMVzLg9mTJmnlGkLE3
8Eju8wbRr1cze/VfVZa50eM/WCU0vaO8x8TJOfh5Q4MIb+4KpPKgatWHFMM0AFcu
8C7lmen8QAz90thzLi6ybXvCzCCt0neIN+wc/f42/qIufP9PFKEmAeLL1aiVwDbO
vD0piQQKNFADPHqmyG52hd9w6uJZ565X/uQ6A/A7MenwSnQgzjxG/xKWPKg5fPLG
Ccfi9oUIrd9BFga26K6zZuN/UV7EzgXslsMOf6pQhzc93ka+u9kClvLGNNEyw18o
QABcKj9wOVJMaVEdkVJE6Cz6s7NlVV9ZPsVygBZ/VtkGi8ZfkeWLGjuoyXIHZ7Kc
5fsNTHL0eH5QMA1mzuOml/BGsetRiqtn0vNGx95SOw4ltA31X07248y8C9WddwUw
mx0aA2D1fka6b9nrhitp63Dyn70ELHiKgeO6netPP7IJWg/9jZZsbt4ISPsZRxXo
vtx0CqbviTrJ+Eka2obbY7WmlHVRqm7QKF4n+xfQq5p6QI8nU6wK9keUkdg2cOo6
ynf5dcG1qvV4CGPlTC3kXMeO6RZddH7UDoqSf5Ybr3+fK+UhmV4N/iUe70K/hdMH
8lwMwnKlm3Z8Q0Z/7sq52tvEVJahC3m1UXCMU2rqJuncWLMCcknLlKmL0dYk2yob
/YUl+03LO9iVdY9m72lQ1/oOTdaWzNFinUiMWNnDk1CytJb32MNAyMtblrKdT0sb
znfI5v4HJEiDJ9OQ0seRSrDh0Sv28hn1dNaYlK9SpmnJt1V4ixP0x8ISz36jmdin
O98GFHTRN3+0T46URJSP7RYt8cMGoQShSQWIvjP8KwpXtCM/jZAXoXi1ICMuC1QP
yg70x62e//SGfq5cCBRr1FZzaplhvrc1q6jQgrysBDsS8p2jzNM2F2D4LRJE2Q6y
DKNgh9QZR86MJ+VgRmdemFXq5+L5MHJJR/OZtuaA43EgXBW1A1BMV1s1fuuXr/cS
h0UcwyXpYJvUoCjKhJh0nlv3gYexENRVSaiDok4UzJpUGfHvTPo6cRfYdyUxKarq
w87WqAPWLzq8oNoZuwNAZza1azXBXl27kZMg/N4e+yhbQ8BYrz/KaUcXrmlneFAf
1uIYU8knZuuDfFggrP5RYf+ecECo3YMO/d/J020dC9WOiQ0MwLNW597yCVSljySW
sKOI7qERADNjY9xgmsD+ZL6qDdPBM7aH6lfAkk06ueuzDP1GK264Pk8WatLr2GSL
LQRzldJ+0h3bn5B6ZvHQDbg3YFJgSPVGPtRISIk1G8CLXPWuAxZWBZstFesV55ww
yLZftZNzunBhRpiMKSngdoTrbIqgwWwZgd4ZEP+WxlTSQjpxMvLWKRwB3fDEte6S
2XrRtIyjqNhAwS4t5DoCN4qxxdrlGJmC17tY1HgKAmRFPKhtZz71j11UVd6ba5KS
o/5G/QR1zTW5B7sOz6itrBU9mNpFym8OG8I93+NG9sza/EY9mNsYT/NTpFEgLcHM
6BJIqy0IIDNmlIeFaNV4Vuu7o10bkTHEF65ZyrL1mkLVTZMVDfKQlsHv/ISdseZP
0VfvHw+23kJlBWFwts2qDivQ/QFfRyu2AVkej430pWjOa7S1H1hEXKzltK+SIFbG
haO86hVYPgXeIcS0XBx+UwVeN89Cn/ivUP9Gj3fs53YxqENnKxw/a4rNkq5hRxBi
zgkDbNhPJdBe5HfwUbsHG8ALrtVYxZleUZXr9ObYRFlR5gYAMcVnS3M8GzKukDBZ
YgJhgI9Sx5DuTisWV3y9Lvz/bgm7Mmfoh6DuMuhCQMGMpx/Fz3suRPz/web+08v8
Ls7o9wQ79ilqMVp9PMjAv4YDMcL82Rs2C4bU15fn2cDAq+KnoOKOz2oM8xGbmf+O
i0/nLpNvBzqjKuUNKgo82GV9s1V7Frc/S8OIIq4EF9nOdSPeW+/M67q7xJ3Uzk7t
JP+0K6V/Bk/ageZ6K1ZGAGiiv44fOpCBYOp/BdTKHsie5vNYXM2t4uS8Ov7Y8P8s
CMvijTjQdKzpyJLMxujciK+C9GE95I/F3hK37pycp5aDGfjSzQ1MfDCpa5s3+G7R
X6y+p8k2kGS1R/AH7vR9wgNrJwcJYPUWOkfZk8mroQ8Sy3egj+0pVavj8M3vudIT
s8fCSvrf26dpRiAz0+zkoA2vGPcA67LrGbjFT3/k+DSRWcF35bOcIH+ckboFdBjt
17lA1cH38aO7jMRkwH0QcyvsITg7iq4AZhjmSmpeHYGJyNXFvCJdjpI2SaCmu8CP
izaoAa6b0ViPifVs/+cSqnEDLwQGtYt/72hfR/L0Lgx+pVNKjT3vVMFXjixS9p6c
YZvC4T3Z8VoglKOzPl2WB6pz3O6/bZ4+JL0SnluL57myLBdUUKZ/ghwLmoOKUzF7
82N5shhmK2Gd+gloXfh+LkmYSJUT7Bo8CIRRl6WyG8Yb1qFzYdwsNXNyAgSO+AwY
oXOu5nHSxsjVsmV5hXbj2MH2ICCtSnwpBl4g5KkLxI75FkDYRBVfAW6lYq0uob+R
NM4OOS71lDmuUmIzXpBD6YmgqXHZYcqYGYb0q0+Q4iwhz9DdFqjANfK3NlFOWsuo
mX3kNfMAlbcnzpsFT5TLFgsonusEa5CojfVQxMLmKjdYNP5f/fvH3x0auTxdX1+U
fKA+VJX7m0ZKiruSLRBZnNArbRAamL1AJp9Ti9p7k/Sh2Zi+nKD2g53qJP2U8CjJ
TccbrsYsPN6UorgXdNQ///sIckOy3fMBwxxd+icDkGAMStcv0Q4v+pn2sHLni99p
hT7dfrcsD5ZEDyZRMR8sFNLHFXx9p1xX7XLJb1uzOJygNOJKsg5+i9zyfeSxNNDK
06yYv6+brJWWIjr//de3/SGNYzYnOdsB8iJ9mLMQoeBWlCkaPhM/PgO7kdd9ghPa
YDDGo6Nfm/b9G/7/ayTiNYFF7l0GvzYopaWjwcVTiFg9cFk0ZPBDjUq0OKOp6Zhj
GWnZLZ6MaqNL1QEkG0ruSJHoJ8Ru2RskbwZqSQCIgxKBOyZ5RWdwZvBF8WJ6JwJ2
t52CoIH3fU050L8VuQgELG1+GXVxIPEkPcmiArT/H06kRE0Uz1TZRwIGBQkzJXGs
Uo3SmoylZ82HAFwoDEOS4MJpdn48mcZDcddFJ7dxN/Z6dPHcDVZOkp6LKdPfglyS
s4zwT8UhD3fNcROSZB/r8wi7RqZpmr5HEMvmcfDNBwxq7D3tJuDiE2F9YUCl4g89
n/jJl/IFFkvtfGyFJyEw3PqLU8emzsnJHeIsvsH9mHsb+fbPgQtKl39I7aG1g8VK
CxWHYAMlbPB3vUIO9yh3GiNuOXq8tVpMzVh5g95J+40PGzs+d+ll++McvfD+eqi2
38sbm2wDs504vLT52anCNT6foShZpF492qD/7m+Gi7llmwjfbYoOf2Z5iACXDCrl
SC5HC15WJJjSSLJgvBnT8q3JqBrrZoK/2ZUpaWO7E2+JIaKNxIx+09Xh+a5EqJ6a
r1INnG2ByYDcybQQgXMrY6FeWlS4PdmOOFK+P9wDvfPva62j3Gq5Uz+ZuBfnL9q2
7wjLq/mOHkGaVX4KuOhEoy8ga70YTgwM5sGgMmQkYz973cu0ZBJUdd/cmtPwXVlG
XRbPWKarg+4j6xylmqSI+Mgru8sSDLAt1r8fU8/RaRK+XRr90htz05r1fBxgvB4m
NvfKzj3em2JapisM3Rsc7eyWp3PKus4V3to2BzjafsLctkeYeqwOghihgjVlcolu
eM5xSCp0ge1xZ6bdyn3hjZB+tgB79oweSRiyK6TTljBfD4z/J7uj9fe+2M8/x1sU
o/cEJzqgnYpQFKqJYLfWJMwzm7JHdzZRTRIUIpf+36QtjUR4mRMpW0vZPt91Q+eY
OAqpsTA5riTK+h4G5xrXgPHGAQivll7KcgfQR/2aTm5oNf3dqwyvcJGvTKhPV2QQ
9GiU3rPSaN8jSuK9Z482tAfm9x8oaOzGsZQsluxW2VpHz+xyMKSWltC/5Z1mfDDF
GmuA/ZbBnb9+NqlA7YPxv+IgqI8L2IGLVSzBaCv2Y5wKA5L4bBFEvzYu+u6uYjK5
G+5agO3nx3SpCTqfEjgYoBSJwc4CZZ1xDD/6DDv9S7MviA3s3x88WPKAlJ6YkEss
X3L6MelA8MUdQerG6iYMamCx1WPZGL2m1dcFAk58lBIJaYk9JIzkXsDB75bPo6Ww
9QxqwCDR+TYv+XXGuH1Z0/02YxUpB7qHyujVG0Am6PDJeQT3OKSlAO098X7tA+O9
uOWbppf34G2cfPIHv/PUMPNwHu+dfLrwPhXzIOLcIVBz8bUSRmoN6syDOYDdaCED
8keFha2zaNzG3FNO/oFIJyTlgybEQdG76EPi1uMQG5LJ01tHDSHtl8RVFWFW6rJu
u7a0Zzs+1eqcekjqwi7rGwNIMlr9y4FdD5aLI1MXeTwccFbXruov43d7mDANnAvP
VfsBrOFPo33ABXqdXst8HI7iR1xmd2JPxwoVf8VJnSqqGUUFonkm0de98FLbBrpD
UsU60eWHG4/AMajEEnLIYzfDFMnvLlQC5tRCPjuHnh1qFCFxIm/UTBmZYonDpsqs
SbLBU7lfWvmcJsACIOr1YmO8Qfw2df5c7KimNDHEnK2RmC3O7EduTtVbgepZANXj
57PvZWwXn8WbWW0XvduJXc87zvW/6BFrTlBCUoXN7QSWi9xVuvqmlnyLVjaGf49W
0tmGv1dl9Sax0yh+yT4tZ/XGo1AmOOJK88trPZwwr1/Ymi2gxH5HyHGm3825wmsD
WFuWpB6Y/Lo7Lte5Ij/sDPG4sXIaRk8Xc1c1ru+cwkt+NmMSzEEZY32EIs1jLORp
g9GmHfpSpKp1kx0wGOpJlX0efy+r3UWOdDlq5iKRFQWmiqlTzrdNqn3iLqbrs0jW
L2U893FWzkZYn/RTdT10rX/zH0yV8hGrEnObURhNUnJUCOy2Y4X5AihvsR7wPrF8
N2on9hnzrigOZYspf8ZV2dbvvQ9Cxxt+Z39gC8EorFT+KpWYONEGepzNM4aagJui
fJGawsKz63ouqBnp6vJ9UjrRwveU49Ii1PEs2OyCZLiMAgXbSk6qk/wHtzIWHaeS
3NHveZLDpNVak7Iz+pF/X476s2yhkNExggl6ZtfLSw7+TVBMdFZCOkbokedaokoy
TwGol16lkPTMlQ1pqVpKu0Cbv9OhbEawkP1071R0ighXCWzEwz+OFR54RraCyKYG
JxQO/8zzefWgg1uJxJ4Xgkakud2OHR+blhmAAMCiQ/5P4NSjP2OdhZk8yOtDLQtZ
fsd9HOQRj52ZF8Kxiz8PGvw6nItLT1rA8qVCDaqM7I5cccVBwOxs76ueIc7c4Uqi
9HyJdz977Eg6L3ZeQWqK2/RJnMCCplBYS2YoW8FfNSGjVcxoT7PC1qg4XjABzchE
7w0xgJBRXA6Q0sU47cquJHm85bWtalcdEvXLGRgJgw9lt8U3PD46GkVBAtGQctCj
8THlpxtOAAz6+SoEP27m8LBcKKEiyhOIk3mX1wyMhWHWqpY1fwi3MmPtYMK+a4ge
chStx4Zfq2BFlvRgJ0j8DPrVLu+1IbaKRA8+HXmEA7hyJoiYmLC+zdN7aeboZ2NV
Z8PpXTNUNEpPA3ycEvcvjYCS4gCY8Xm5SO4xP7ij1JU5UElODA2NxDUxq/o49EY1
X00uIA08Pw9bAelfiJ70CRjMgP0KfbDbxfODxeUFQFN7H1INdkJLSzY8Ir6dkxGe
rorsNMyD34ASkIS5YGY9apOuMF7IdI117pVwlCrlFdhidv4FnDuAXZeE1h6LWjjj
VvKgiH/IUde+lGdqBZJSC+AnbcpmDSfbuIzuIzK5tLwjprfxmMGI9mry+ox19/OL
lSo0ox7CV9vt7SMGPitek4jrW9uWqKQMoeLlAmDeW/mz7Oe3x3qf9NBQS7ng0M7w
iRrbYCu47jUm6eQ4HkfMb1LDczibbTuJX4bbLjqZXcyLJryGNAMyVs5HHf6W4/VB
Ngl6VurGcGLemcHCrSyST0EtTrCty9Yh11TLTbLTOvCiDiLTPvk8NpcYEl+Memr3
mHLlPiLKsanxgrxdPzpRZXGvFdXIfqttSOh2PhzlBEhD9ScHAsXD8Yv9o0eEvnDR
GwNRUe98HZi9uGNo8w20dL7UxK5TQzG4x1YGdux+QdyvjfXaHoLQrm1A+wj6M0Iv
s7hQgMkh01r5t5Javjb2i9Of/7Xp6XKpwSvl0iWnftuZbSwo/fbtBogDPPPtVTGG
6tyH6UL6r5Q7rv5DZpaSswh2w4vRA4cHr4P6g/Y9Z9A/1qqzPPHi2r9VA1QSBPXe
NV05BTB6BzZEzYp+2oVfz+HrNSp/XCD5LCRHSr6aM/D/kudSYWaR3/TFojznLlq3
IH8rKMaDVxR2Q0nscVyv2/T/J7Bzzm2Qh5qdYYcFy3p4Jzkcb2sSIj6bj0w6f/RG
GOII4V7jXWeNyPnUR3K6rtylsen4WgMVZZ8W+Dg3moZO6dt4B78BF8PoOjSqTK/s
F5VMewlpOHXu5eCgs2/+rcYXtMf0hSEG5izS2ECrRNUgboVzVEtgqql9LxeifAmh
Lc1smAAbVatyki+cvMJIPkxM8JHvffIxb7yt4TWu8OraF2plLFOOs8Dw0arITyLw
g9KG6Qu1Zu33Ap9cnx4J6r3E0U1ZgYTEf3N3ur6fvbV3cq5HIqyfqFSdHvG0eZQN
F/0Ft1e1HH9kKpTb9sOJUhlpgiVikGz9lpD6CNWGvUJ9Ugjq9shcQhZGxjcq95vb
3vYG/yMzqso9idvtHk2lJC9OjuwE37NmGXjEpt+y6r6L7wRaQS4eBwH8NYTh6vgk
Sz6qAlVDVLAlSFuOA3Ezd2Eb0stGon+Ni6qbozd8swWuNjbZhp8av77x6bUn4a8Z
A5W+vWEFjL+8JOv4kVJQDCJnKiowIj/ye9JfZFuGat5sC3FwyCdemg2mJ8WxCS1P
D9V5AZLcUwNzL9WyBrpNXcKssJnYYUtUV82T1Bs3gtMu5rX4KwU22xh4F+HwpUWC
P7K7JVKrvHjsIUhpTV6h2aeETIRVtQ5ac28J7jr431SnbFsIzwqYRZ1CCgGaxeG5
KODsjBDuH3vQ1LQvUNAH462ENqoysU+GgYD50PYs+mpJlcIG+09ftqikmZmfU7Tk
l7pdA1suuIn5YV9uYqJw1aVEMGudswD+SdWRJ5t2riXDw5du+TCJ8lDlW2A4ogyx
akMs3yWM+zvAj//H9D2ne1iCwAx8jwM1ZxyJxMs8iXfW1p9cBq3jsrSsoEwyIZQl
dK8OLVM3Zx6miKS8FYnlqfkCi0R6R9oHKEV1V/Rd7Q2JyYswyX28RzMlx9jdI88c
Z0wFldRLE63+J+3enVG56EcShsEBnEB1nKjX4ITO3WyG6FfHyquNb2+VipvrCoGJ
SXHYRw4mGpgsk7ZEDqSpbxTTH/CTL6bo+UcQEknjTgTLFu+kHtXzRskNawYpC35G
2S4uGUzW9wMAFVrxO3WOxvrLKzXi0alxDQCEzDjyBDHgYwEfjKvkMF7LsMtjyA3N
51pMW0+mt/mwU4tjOl+y8XX2jUwdJhQbHUHYlZd1FtQt0YvJ8Q/JM83fYMwrKC1o
cV94gV16c8YfT4IuLu8jmNMc9mthILlypEwhsXrhmhfzwYtuirSeqeje5WRB5uey
1LGuxcrAb+S+ojKHG2nr/KeQpFpfyyT5vs/SoGV/GzaxozSD3VzIM54YI7/5YlT1
aHrtHgrD++i26UavAac66gOUw6oiKLxvI/yTfWgDnPm5P5nH1CGAfEXvAsosMulr
mcq+8V8dWQP/IUKRWMBQbahQg6Kbe2NIQwclzePxjQk4OyEvPKbzDWYK2RJBs8UI
yYgwMxZNBX4qqn25MKfOq8j16CQK+ruArcIWYj7vEXfxeSlBvuOWVLroCwrjsvEU
rENAymQuUd+af7dSTpYcvM5Z3tye/Ynb530ddcHIDWr0ft7Bj6aM5jLAAfWvF16W
kJ6DxfJBmacsZAXoBQK7chpIW5KXw44OjsRLAPgh/4pTSBn428C8KnM5toN4eKkz
jgvQlV/+C/XTJISuOTEoKDeO0aL5M7JdQeWBBITJeqPGJ7hzSY8Ib37Spy6S9aSP
iajljUNJjj0orKgn37L3fTsNHigt9og0/YfJbAtTQYU2VKZxA1kjVV4yMwEEUXt+
VVRZv+LGixtpKFIRJ2XTRUusBibGRn4L5Q9S90rQQ8gipLdjPK6P/lDUjDogmcp3
PD/kaSSVzwM3Sn2IYB2TMnu3GdarY+Tub+haFdyG2eMfxCkhOE/zrgEIpQDYQF/y
HbrEUmue9bApb39ussK4lP+m3RqBdljxpDgvgW4Zqaqg5rd1iect6nqsoHEGeC0c
IjbKqjBGKhUvPd074t5JXzEKW0cRHrwyvH3WUG4btX5s+mYuTz9HWllqBXJvn34n
MBTJq7Ln20Ij4Sra1ig3C6n4bnK/Gqqq0S7Ps+S9O4WxaqrQTE127aJ+O5V9qp/C
wVbFY/Cdvu/LFld1tefeYXecFe68o7Cp+Q/JEEwEOssGGf+IVlMeNeh4m+yDnKx8
GWFwd7FCQoRle8HSWy81P/m/mh0pK50ShN6cLlbkOAYXw7w0k1xv1PYiZnYo31uh
ZgbTqE+T9BguvOVAdGwyyE23vn3YTyd8GFQPdSylYwXyVOMxvrKEnfw8J/sTcPpY
H0aavkk4GtGgaqH0nzJb8btgC4XtapnJy/dbVYCfM9BhFoRlSRqkXfdExspIWa3W
pFOYXC6u345rf2yPLO6LBRFFP7Y9oJUO5iJRbvRtLx41bwNCiq6yfg2scFS3w6Le
uks3elcRUcEj3cVx7j+k6kICeEDtNLXcu1pIb9cprGG5vGubQrYpHPV6NMTGDjNi
95wOnXTFKZ3gnbxpSo0dS56GF77aMgJy+oj/LKh9BHvC0Knu9QMUTmRqtRg1KOHi
QeWDcOc6rWVzZLOpCAAxo7bxHRlTJrpe/kI+2uKwt9hGZ/6KNb9mkUlVChJyTtmG
KQuXew4htjBnmlRNqcqsIcIOW+tp6tSYHpYfC+PbtrE65xs8YasJn/d8Il/ggSeW
huVTLJLh1lSUc72f0JbzLckZur8ZWcmtMW4iIhKfMExM3KADXyFJOMR7fkYF5jvp
CEYvV68/kziFwNaM99hSLVKbTMztGnILD/5v7HLumiNWl2/CQOQ4jgSwePrsKSo/
fICHa/ryuYoqwIrWTAsMGCiZ4yqULfqQ0THE05HWoeNWopNT5uswU7BPkPLu//Jf
v9CQyPFrG7toXJrS0HMZV40jfOodCgDZ4GeWy7bNbp/BV7x08pFrCt7GaKWmapf/
dgeCO4q/oGjteLpsgF4uuHtIoOjUX/ofp4Wll5OITXRC+kBDnrZM4fmRu3ZJn2zh
aQG9p2BsDqVafv6k1e+h9srKk9U2S+SwK2QT3xWonB2WMXYhNIbVRi/xYxIjtfqw
jRd7c70ok4Yg8iFPsuiEQHPFQrY7k0RmQMzXs88xUv89l29BH8U5QwS+TeYMwxQs
p4Oh7ZZfYvr6NpC0Jh5A6Aj3if+6ON+Z87/2eiRYDBcINab2uh62Iry3y2TzcdBt
GYZ5MINyrq38wlnU5SagBMC2hehaV7Ely31TFLEoU3XKqyIS1SAkGDjoNVJIi0R/
hGt9T81m5EHbalJO38ES260pgnek1XtPOYoy0LKCHwdEGlDMjI1JNJMIQjhO3aM6
if7Jgtgm7SrC3GMiB43E2ranwC0FYIHO3qCMwqgBZbz6IjxZEzY6oVof8hoLlbQT
vePJLEmDc49+bQrWge1WwctH1sX8yJN2/jHgcSNubKooEp15M3ItEYSnYd50wS9o
+ZWPdZs7YTCCyAQ4ZdTAKLxuh+I4o8mZLVI+PRToo3knkBUcMkJOs8rG0bt1nqiS
LuDtlag7OwOOD3QYdmp96FVeBo8WDZI40a3xZutQzINBeN6eXyatgN7Jk4AZAaFu
emwnMPp415fQug13BtsYeFG2DXYfAU/jqrxykBAcsGDn+lxhyuQFTj30Bf7tXD6t
muGMUL87YRESbLWp8vhnVVY1+vzxyFyJXRnIrVWMSENeSRIwRFIxf6GjvsjEDGlB
Fs8f+REpDuFS+B0kzoSkTPssp47XdG7+Pl085JCjZAJxauCVFqwgHdwIYMXecV2/
+bBhgBaRGaFMxyeuUmMm1pyH+fQp08Zg+86+56QPiaI4oIraGOU2jrGayZd6MM5D
uhWoGc6qyeKgbcJv+57Easw3Z2G1moU1XSuG0T9vldxtfPvmo2oiwkur6cOkmdLR
8MMKh4bU3wEFfXXYgEkwufCCO8bi7KmgKQo4qD2o51ayVCAsKU5vLTVEj0cXmt5/
IEoxeJVdSRJclOqtQXtdJu5wAm/hUpoDCx9SnE+Yu78+rNFMKaq1ZVMOYcKwYvIo
4ItdE95l5JITDaY3L68mDDhhmOwHW/4CI9uv775f3+eDGQsPfg+8VSTtvxUNEkwc
JdQomPlLjpZkgWGoiYVk6re85JFNiDyOs2ac4FnbF3HBzIcuMrQJrBaqRdeqQwJV
vZf35Ab0kB3/MStgv1+gNKEa8O+qQjCcNUluMx/kTVIUou6p5u/OJuNLVxt7LS3Q
YfNd/ZNuOruHU3wdcJlkI0Xz+z0FO6knZFjsvi+/7JtOyS1XW8pbbR0+gf0EQhio
98vpxh9L4XAvIIquULksC1+BqlwYy3Cp5uH51Z3plrFMoXxf2U4T4OTN4v/Wq9RQ
uuNEwH3MckeeC0ZKbZUS8cZeYgRLnhjHvURdOKn/aG26mkxLxnP6eR7gNrOn7yJL
/dNCHhfX5Hnr7boadywnynFdpokwdIhwaCKzIG3poQhs1oZBslyUWKAHC+JA3OVA
uy7y+GY3X1grib+QgMJahVlgzhiZjFGbOBYrU6QhBqqISMfcAkNldSg/E82/Vsgd
Dk1xgDcZV3emoMbAIlYKiDeGZ9mTzNYWRK694/oS5OQ5YkHI/b9N7KaHyFtRNaUv
joZBYWRi54FN3F3o/LuCMZttt/LF+PLIu2j1D7dxnvR8bYADw0h0Fyejz1raDYM0
SdAgxMI3IIdEQMCrAZ9mxlkNN9ZHuGiz5YLbGhW0qDuhe25XtBpMLCyGhHi5ek7K
857aPed4+Rh6ytwbchPaT0xeFCea6PBo0Ulc7aZZGqKEIHFYNgrTR+wIuRJ5CFBc
7nGkT7urSdXdM8z2vyHn/89mG0TZYF4sa+6qq6+w2nKLoi+5kMowSU49m+fdgudT
HASv4TJwoxrmM0P1uYVODGYWuoqQbgRpbnmqN0FROQ9frri46pdUIiGbH5k+zVr3
PJ7v6nKpOJibwdt8Kj+LiQBaZ9FIsa/8DnFCY1Rkwsz5qxA2ISE1ctoSeYIOytpa
L7je1eJr6BQ108SmNgy6MbuiS9N3OBgWq2s1GEtFmIzFOGh4x6EQtnAPRQQWa1e8
0p8bMgukegUw5GsQ4JYzFE3Eldhoyi4wf3+FbKTHWhrUKN9OyA7D8TXfBLMa11I2
K23xuIUQtGXDcptJjWsdZyYp5VkfYU0BrZM92X6FoAtd7YzsfiU97pmbYCs8Wbdk
JD6yc8vSQEG7wMFse+KOzEVBj1IkDPG1e+Yi6NT2mplfPO8C7MZ7+I0xAYYs1MzX
+FGJutnxf2tJ4wbTApOIPyWhMT27XRzViuQN4dI6JYbuliK2l17+7nCfneE5N/+J
jjS431Cr3yEWJeeN90PFkHjUZRz/pomUMhQTYKDEk+OGP2QlcsLYQhzy6B4XuWWK
eOJGJ5xXdzokA099/0P4sOsEQEnaZLf6hqqvteV69wK6vy24cA37wt2P3DNh4Rk9
+J9pFX4D5QJwZTm94+tlVEIKDT7XKvL4Av24UhpWvSMeyVYaaXgvqzGNTyPtQDN/
Fv5DD5c+ZTZLFAH0/nnE1Rw/Z8u1ToS+G+x/FpZnlB/OMpJU0ItdeSt3LSitIT1A
bGuwibzCze+Rz+te9gzSSt5qMOj+mhbu4TYaqor0JbVWWZ2LAejwaDxRSqyj8yxd
mQta/VDT11eFKhOVlF0LowceFkSBJK2Srpng3DCTONvvsGaRUfcrvc0iPOTU6D78
jHeIK5qg79DENs/9KZpZCMFR/9GM4QBCZPtsGnm2ReaSxM5ZE9UwcnWjWg8xKziS
4JiYVOy2d7+0vpGPJHyWmqkjmWemCN4SH+NFRMgJnFF2SpAmvLP7Pu3c8uWAnJrf
zcogR4WGsZ+v2jd7FTKcir6B5YdW3E8bVrhMDiGNFQjnnZcu2wCGd40Q7AbHvOOA
C99DkgNNMKw0xIn6R7LNWQKxM+Vf+rWhWl2wf5lefeeT5iG0WfM+ZUzUv69fqvrv
BsR2zBItWolvLJA2XBxgxMfAiPNSmPNbwZVDDgFQGZztD0XS1I2HQTsLqZYZtOVC
p/rqVMxaWncPrgZ6O/KOksX6VPs7RN+qG79yPRapC2dLeQLRvLBq6hF8j3BfXV5F
Os89UbMp2xxu6RLBVXsILuEOpwfmTk5hdMSvpZf9PxbTtdZg+erqtzCtNFm9xHsL
gbomqMkXvVewBCchOcE6M/erj9WuWMA/BWBqKn/UW42WRxXv/EmPyYf1A/RJLAwq
xXPBGxQrM1NBDS0IbvznaL9+eaAYwHydcxhMHTSyTywreGzA2BQJab0zMF5L7S+o
FH6BP2YSkq7sC1JZKnc3aeytTmSBNI2qNQYDzVIgOIN/jr3b07abZ58tRtWpZ8dx
f43z0ol+VZYZUG6Shjwvdrwo5btIHYrtlP+wrRVcsFdLasViO5TrqYpN4Me5R5rv
KipuWxzV6hKS8TU+B0gJ6rOxb+Iy7oE3vDS95gB2ALJslQzteqMSUUOjTik6w93E
SGgf/wYOO4W2ID3PgL4cIfL9lM6X1eObvvTCy04/b6KxYA9MoTA/XJhcKg6XMAFb
BhUCAwsI/HU2u0027SlMfcI0q1VjXvPufW5B3mFAD729gEnKJmPfr3r/hTW5sF/I
KhcRNaVo4glItYhzZXJ1AsYlBObQk0uPdWLLCLRvj+nb9dFUNnfK9S+bi9GzlRyU
29voDTwgLe3x6yltqp0b7FzI0LfQlaETJplPi463zAeY5EqPGREAv7LtARDuse0y
qkChQ3jN6CDxLhvDqw2CKVxjGOTBSkNqhnZDcBwghnkGboDLzfJ0aY2x4bvACZ8V
GH6a9azHNJJvxJILttDSxwC22n4lSoPDNTipJIVgzpIPb012bmcI8j+ma604PaZ/
M1aVsRGGyQMs1E5iCv66nSmtSMYjEup8pyEwn5qFNlxE+Emafoi/ByBMhGCvRf/H
zgTAJUviyzwNp6TphXZFJ8xh4ugyDDACOFzDSfYLRHT2gD8vLU6IdMA/GCnynM4c
yDXUPcFf2GYi52M0VoHd+UpDvXUPaqwKHh41SqNLm6p3wPxBDLNfGPwd3fHRqMcb
nVPLRasvMS80GsWzjCD0hJxTPj+85JlOW6bCczLgIpRHFebN4w2tSV4RgomSrTUW
RIH/v7sEmKOztb5mpgk0E4tl9X+mJsyjoT7Sok1tDKYMkmau83XsqolpZD8Y38H/
PgcAPBwS/AgYVaEiva7wykZ/+IpOFYXGNtM5luB1XZWZ5PEllsGZiXIrIBfjhLdZ
q9fxZ9KVEyRRZyprURnnHjM6rVz+mNoh+Hu6ctFSeZ9XoD1ijkvppabia1GY4k6E
cvp6M/+wDdelcDhWCxgjci5/neak+E4Ewr7yBS/SqocL44OXo25KPDNDULe9lF0j
bm9Katl2Gewg9qbJal1GhvYe1INhitwUtXTUjNPEaRGOqmh3RUxS6XtXxrYwtuG6
bZInbvaAHQ9eccWyjfOnrz+R45SYqwjYrrFwvw6AOj80OsUJiGAyjMvM9Suy9nBz
q8RAgt5rHAaKIj/deVoOtOfT4tshWPzEzaPiQ3ZBYq/fE1hUWah7dpXO+dlIGYTT
7t1heVSSayVJDQ86iD1eDeyGqFzNPYXoUMlHS1ZieA5saI5Hy1EPdjAQBJ8n+fWx
4FXQlVlUNnheXEGrXSVWWg1a5AxPX2TvxR6ERtCProIEZNSIJA/wSJjcdzsOFeFR
NVeVQxvdRUJZzcK88CbOwZXVB3NJQltQsekevY/a2E3P0+DpYO6+xOlYgugFsTz1
PEOuD/7P5dy13igyndRVcDrviYKpED++E047K6elhYZ92bJ5iuY1dFe/RZz89akT
H/EyNvjvCfiQIg5KHR5ToZDAalaX7ezOa3sRqmD+nspwcsk3AMrKAV/tKJ/uAShY
cvtEJ5CcYMXEdjOf4FQ+rnEvTJR1vpkBSxYdsUArnxI6Koel77XOmd4xK+cydKMu
6gwlOVfVYC8Zt3CvRdgMxnjSkjLqMkEopBw1Ea8jLK0Pu94n0elOk6QMCM1H6OrR
yZ4D7ZRPCSZPPi5DFBRM50ps5srTAUhmEbNhU7zToO4V6L26+nbuDN9EEVXQtnOB
+xZ110SHvGy+m0QgKfoVIguB1TavIF5R2O2yby5V4CfeGRK5o/VFzaGWsFQHrN2u
8HLroRacJfFtCPIsP7+tAfztk7dqH+Bak/86KNi5UB5UYB79PNlMdUeleN5scND5
gZVJdbnolu6TBjx4hBduHm/U0MrsBCvEh0dn/4+SxZ7+BfhjJL+ji+EA5uA16RsK
9PPEGyzEvJl5e/DedJOLuEb054X6dGJjKudEO0n0mIKp/fHigU+4L/s+H2DUJxT8
9feOHY0twIvlG6ZfnAxsXAGMVxefc1U3jhokVittqosGDZO6Fvi7yR6bW52/WC1x
VTUtGmEa5jcNtUBSI7k4Mfu4nx6fGh5MFmctczhwZVcO6eICsZTt3nNHXX09ehSS
Pih/8DpNNL/LeQ2W7q2a3ZjlpXWYDytVHdMGqTDBuwdzVqnuJBnxM9Lu1XM+SfHV
x8n7yC0g0zlT4+1LgwkZSwQdJSp2PZGutEAVDPCCRvalh11vM5USqPfPSN583v+G
wdUk5O7CdRz4Dlb5H09L8CN/Em3NxsOYqo+ea5IrUkQQBXXFNRJ5gU+0vKb+Udrn
kiLg10B1EoYi5fXxOyNizBkMne2amAQkIRJUQoCvpIPqKzG0jwHWnekiEayywzvq
1q+YIBEl6x1E6qmWxmdUA5xWxL5RklA3OokEIFEiw0kFbxVc1jX1NjOYtFF4bjAn
hDqEHZGtU9+ucXLOEAZ4hvZ1TZEbWzi4etF8NLd467ps8xHrsrNHUvCpLR9fTxKr
Yc9/rBxZm98YntwGPQy3gPTx0gf6rk8zAjir68nABPVlJzDb0suZ1+j5i+92axVv
OdwGY1gZgdpAUstD36YFjP80GlgG5SdOV0T+kqJSby3Hg1KaSmAcQvcRjs14NPzK
NqK/KXAgehQHvBsbySa+xKFS7k8d1UwaNGDdEH8gYdm6SWaM/X/VGJm1efsgQdoi
JJ6Wva8zrhEM9/bBIwd82sJ3dwPc1GW7x3lQG2FKGXpi/tZYdCc9IWD9C8bcyHPC
rw4D6ocIMMuNiwggVzCYKF8IQG/go2eLa9SLXAFLP6VR1Yp4ytcmEf0z05+44BMx
PExRHWtUCFOa06NrtS1L2UoExuWZ+gTrbRt7E7Q86YsdTjH7AGiVLUZwyjpNisFA
LZxMDV8t+u6wft8ft0V8ncPihlo8XkLJr4SXtrLm1ueJ7hff2zj/tqayE9TH36Bc
pT6AiKnibFvta7pQp3+AmitQbNfv1yzkdGJDWb1ppOABGT6DAy6tJkYqqrsE9HJf
Fx77/6Hi3mjkwFjAt84geoG/da+uA8mr8eJwZFMz5V3a3InMf4Jxt1C3sv00pUGj
czVQrC1W30X9ktJiUS0qfY6Kz/FklVlrIacUnL261oZFjXqilNWph+ZvTCyoc3yu
wdf8bOillfctBDcsa11wxC5ZpiGX1FW4op8Ny/jeOoq6hKzNJrOfGrK5HE7ZCgRs
135GsjPTq0y81lfI0+B8+BLzLC1cLyT2Dac5ZvJAYF7fUeVDMWEC2UBKuoTLwv3T
RDOqoedG4jOhaeIH/y1G0avgAw3XCXtf2eEsdgObLRhW1nLoglO0u04WPBZ/C2dq
LjvcEfz0AFgUsTD//Gax0ViHJv9VM3hynBxoytx/KpWF4IAngg2j7rm1xNGHmpwc
xdTcki988sIwQpAzwdAg3OvouTNuD89/jGPPdWIUt3fhxE+Ngrb1GwCqPGTDRLzz
+RFGUyekzh5EOgiFNsTG94x4c7mcWAYI9qPmmofRrwSfXRYV/az1rCKqYfw6Kq4i
RVSdAChtS3puTT17V1p8ICiGFLnHgGCMQm2JvtDwo4aND73gZUNZyb2rZTmzfDka
RE3J6Mo44nxG/x3L8fb3otZEFGKgrOAeDDwSfdTruFEOeHK1Dmc3IrOAy5TA6rq5
1J1R4Q4eW8SrbHPZwBae/JBpHBJvIPFl7kUPvSwqfSwAdiJTd2KC0m1deAFcK/6a
FXdTi1A6GpMxhzP576Bw0wlTclqJOXhydk9yTw/ycTZgmzTSIWyN/+MLQOdqXfmf
srid3TiSczDCMtFVaEFMbuNIRY6qf1pvGK1bjF8zFf1Apmed7lhUM8xUIbGSOJ2K
gIfnvgwy2EculcwDYU2sJOBfiMrlI4GWC/WNR2dxgCo7t7PQ2+rpHhtvJExWcfrJ
TZeXHa05J0XHbjtRRIy1qVfolKFe8MqyRnIsdyOkjrbEGnw+pqAEzlmFzbsBRuid
9wl9Z09wpBmFPhCDE8I+7uTBOLSZsE9oAGxpQLx4gM1gMVCLPshjWg+SN4UtAIbx
nzOe56GMBcLvWFfAnOBmW9GN5BHVOz+7VwGOx3yc1zF3U1NDVQJ3FncvaTyEe3ah
SwPzPLIQ6KPrMIMnnBGcS//ZKOq3Zyu7T8lRFA2h8WdQ4WhqBSBHg6vPf/8VCiw/
nZQKlVsD8/3tRmQy+t17qFQh0ejdshwIkcE8HUT3aTb05DJ3z1fjqE1SpRV7sY04
8uAx8VosfjtuSZjnsR8Hw/zE0mRMj6lqiGPYRgA7Z582ELjngHchd+ICc9PIR4PC
uxdMX5jeyxWgaRc8qy9+4hmqfjop1tr23AntLpDp926z+tbqKatcvZmw8oVe/Qto
vU4/MXlVNgo5NGcAAcXWem4qS86iAUAUiLzirjdhoh+yrpGyjXOcVfS0SBmEn0Y4
6EiwowoCO6lsDBhBGHtPmChRe78c/YlywaA3tpzTbY6vofzhW8i0LS84zpYWRl19
oCf+TTJ550Y0yCXhWLITPkcIg7AYpY8p6M9w0jRvehrOCT150DNfBC3aBIkLQaZL
aT7vBmZrTdnGw/3ZqfLUq46kXw4UPBTSEaDk/LpZHTR75Ywghxg1f0GNcLGHB7Fv
0TC1vmqD15aZvNsGmvlVeEtjduaO3OlzY0YrmjZ8bgqQGcKRjZpCy3Ko4tkTC1HJ
raje4cFGmkZZQT4clTiPL7qB59vqmUYB7pwWAbgScEQOFegXBSy9TPzI+jrUvEG2
lpPMd/utgbj4v8zGsyHtCkKJGA4YuUM43m4r+nFzawUV47SVl/M9dXlBrg+eGEfO
oOVAF+EZRnhZBSkT9/zIg9cZssQi33nhZp3FBSWi2Zqs4P6DerVmzo7pemJ48g2+
iB86AUTnh0ZXGF/h99mOWE0C0kucidkPfFKMefGYZtaZJ/az2EhRNmqBMF6tc40I
KxH+tI3Aat5NEBfqGlXcB5gMgnfPkDLSZ8gNDit9MBzAyDrsOlL2okpzYwV6xRgK
qQLOIiSm4kWRynsW+mwk1g+X/MfrXYvIzVV9IG2NT20cJi5a/q5GbT57RUqXhBdt
cbHqqL4Gw/BviM4UN/nPqeL2IYSzyFNUqDFald++M91fb/Hn8WaIDFv8+vxjnxvq
Ps247vNdam2r81zqJslhKjadYV+gd5ilI99De5j1uD8Bxt1X9597uKOXxPmc5H5B
rKKX+EaSAGSe5U0jkuB3RFBx9J1ghc5vGQ9bFABScaOD/23Wubb5S3MTh2o6RsNn
Q5PR07O2uJd9rnjOaxXxEn2aKeoe9v0fd0VtHRDjn7NQIkpKIvWnh7jcnHKzzxPC
wBkU2i2pjr+PPqS97k/ZlQCyAIW9JL6dZX1a61yB9zOEnkdnw6EDpVKLYmevzpHi
/hJEglpGu5EPbNk501KGVHh7T2jBFL+qJgPA9EpWjJVTX8k8i+MVGL43nxR72MN1
6rdyxYZzpi3/f9SFU1QnhS4ElRr1LARv1EZrkqMlzuAItAW5ta+PyQfyu2txZvYJ
FM8i+H0+K8DhfAmAOJSU+4eZV3J2ZkynNn4N/DciK0vkEj8+RNBwpBEa5XxtgpUT
vwRY75Jckfzgma0OPYWj27+iTYy7rUbnN0fVKe0MXYxMwZ5J5mYx7IifOT8r4FN+
XC2yLhWme5uYZdhwHalw9WyBnDoA39YJhdIUMUp7pl/3mth+SUVHiSYDjtBrkXUk
FjNsmjeOiHR/wQBQaGrr/Ei60D91N/WEBMneXFX34PBC8HKezH8ST8m/u6iVC2o2
OqtiVk4WjR0Ng629zqfgB5X5VVRP9BH9iU+JojHOL0oACaU1yXn7VBoNqJAUNdL0
axb8MLDrFfWTxj+cHiccH5xcD1nwzs3S6vR4uNm9dW07UxxTJjQN29o45VgU7cN/
5vynoh7aRCVC5FwIzgjjUep1Hf8N2iOUux21ezhxnuR5SmGUpF730efLb84imzTi
399E0uQt9iFtHSjxttCntfKSVZyP9+IWwqjcVQICDNw8jaI4QgXpqu7bOFffJhCG
xGy0Lhs2vVXgp2G+SGmvCny5S1p6XgujVKxbghj+BcBGk5xYw4RP/VmK/w5pEjkq
DaCiKcdgqGp6Vg5nv/krRl871YrQSiShFbRzs2fG3DI0pA9RTEcOjL21yU9+tbfh
fku4JbNKytKZVZrjPY/PGS7LhueB++qBuEtAekvhQSseNrm84FQ71SwZBn/YxP4E
9Ns+iOFF8qS4UURm+627miR1CGBSkRabJTWqo2VXGLV4kGFD5Y+D42qcMhRp9jHG
AH1dMoPhMjgMJgp8aCLL54jZZYhJWMUvYEBnJCTquQiSh3KOpezVYUxic85BoDob
TVP3i9IPyCakU/fdyiPXDiDSm9ETOppQbcd7JbEigheV18CMFx+wGv5g0vJlyA1j
8+wl/253Y//MBHF5TPpMMf+IReDNupepSlc/XM3is4xoC0//uE2Te/lUy3NUo330
h7e99gHcl0nWyIBZ2Nh6+5qQwKoRGUOA3jkUgoe0BlycjzCYm+nuolk85NTtOHtD
JLZRYDXxqJr2SWBlMrSiTtVKcKl79XYsCvu7H9Uj0PN/FVz5Vg1iJGiJJNdtX5ZW
rbLCwjcIa12+IIodN7O8AmRPdKr5sx80rcMrsRDy9TfWkn7BEHZ9NvbQHccpWB6v
KzxwyB3LIckToBEeI8e/Ghp02xikOfbtaxCzuonluiteiddJ5MUlpPNYMD2LOLju
3jpHTyljpCYs9zk9b8ZOZ6SYR6VBpBcnl+d5IAY4tb3F/PEoGvk2opc856WkzmXn
FRWbD6QGyqt9H9zKlxIiURLR8VlO1oNOOdkXydlgUjs+I/5vtsNf6MJu4YMjUu29
Bx7Zapjyq2gWis51t9uOzJ00ZO6KJ7qluCme0TicIKLntRTN8E/CWQhPptrbAA+Q
7i5ULW3HZg61Z6Ly8OXlR5joUKULtlO5p2p+he97iSUZZV/tAgbjyHc2L615k3M3
7CVnATGhypIXkTg5zwKpfBi2Gf8+09zKYmzQtNBd6dLwqs5ih41HLQpYyurvBzKA
BSBmudz+pza3+MBXyckgSpKeHzpwX8bHUjFKKBgHDrhx065gBnwKKCWa1O8pQn0Y
fyioccGjntxULfcFwrWX+rYA2BZJiusFtRWWpO1d9g/KuFJ6j1W3BpAmerwUMZKV
Ps/AgW3VvL+TiXWfVOgh6SvBz8CAt5SuPdO+PcBxmkU/TsXGLfVW1yRPIwDQtBLv
sFcvmIYJmSw/K9mx33lpaC9M7kdzBqhRgrMW92LGY6657pAeJiCe1hDRqMazKhQr
Bh7dI9lBq1Ex+HcVpB/l6LdlSxpaWPi/vGBgXkH0OoLApG0Ryv0+Y+vRk69MxhJo
85hfIf4YqBXx8vqGVzU4ykRozmQGyqftcWrU3gaJb1D7yf1Z1iPkXn1DuxpN8GGu
tGFkZMqEknmm1kkO2oH4jmpWJlgkSa1MyQdtCH1wj3fBchgI4g/5aRAOHvSsjD2v
iEN30h8ouuJSsrWk/ROIjOhGQhxbukZJGtcKqu2GSg9eXkM7Ecn1tiBt/HbhqGpu
I4G76LVoqTOWQI+u12aPAd+N/bPiE5Gd5MAuae9YLcxYTabIabEp5QK77u5eLIWF
fFdPAvMVJ20bNcpXTUha4a2nXj4/x+h9BFvDdW2rlYwoBP1ud2GXfMS5W+ioJXFD
x0uKMHDgShy7JCabyeE3jLJabzKNH+AtvuqEqdNkXiG2X+lsddj/vQULgkDhhFB6
lJwVjqQcVWA2fONaYxa8q2pR6G/kZRyzQnNNzxUkr4k1qillhy3Qd+f5f7Ac77tv
l//iyMp1SNKIGlsSOJbkAE/DmPF4UOl6iUzlBhSM9UVUPBNEaIBdpadDSklS2LVA
6k+EmKdMcSKYGEpNT6bB050riGvayLMvFRMlx8Y+vIps20oYYenEY49TcOwa0aWD
kNzTCQ9Eou1gXlwWPS1ApRmko2tZTMzYJpLTcTZbvGnVQYPGtXoykTPcodrPIb2s
IYmSwdKsXnRl+VBh5XkufUEGyoAiKx1ujYo3y49jEM9BwbFnc7yCRNp20+jU5U4b
H/TKmyC229RIBVPxQE3hT4QDB6hHeZsoPKLcQSXvk93rg/TwJh0naHuR2XySBv1N
y5pds4LsdA90tKHAt7Z0INW6YkyRLlChZDSUviy/pS/FFqQLFct/9utY5sZYgp9Z
9XUfU1hANJEmVWI0yB+B+6/whByVAPedH8sY4ud7O4S+O8ASlT2MjSImRlFjHmz3
c/Fm3GcTs5P2n/BlPPJUtIysNdlPQdBSZC8R1egfXZQhjOA4+VQDVmgtn2V2NqmK
grr08WLjumUmfws3JOvaP2COxJTeQs5UTDBBaoBUv4XCHtRrrlKV5ojDg/O0ljqW
gtkY/kg9to+ZqL+08oARF+VyY7qdsG0MZDoKxA3zjP72tY6J2+nZInh4rUXGWRE5
q1yE3gl9IJa6wb+05DsIquYKdFkR9Fbpa8LtawEo6kb8RbHZNXtYsEs9avUlLfPO
NPtxFrXn0xJF/WQycShViOfhEyTKnG0Q+rdv23KmSjwz1BRypjoHga7R5CtUBOgi
pP9hZJGI0OLlbQtSptWfYJerZtSptztr0T6mbrjU6VuyYlxYJH6p5hV9MaglgEJq
NJy4lrEBnwi6/cS4GeWVN0UrOQkJUTmuLojIesu9QzAEsQcPg0OMSFF8OM0iiZmI
JgvoljicgqB9XHiF4VC5W19gHaHukQjuPTYe34qDLRLMi4teTyKxfziU9joYGcBT
7W0jsYmEMjiEIc/dikTNtoXuYoqxCUXIRlayqW+KZqG/h7KT9I9y5bil/71OyFU8
mga55RYKpK0Q3PVsE6Wwc5Xl4tpC8iMJZOI+BnshhHzMGLxebxhZuBazKn11nzx/
Y6Gr3sxbstNKJfutYmdauUoXZht+mP0gj6f7CsRDHg70qxUOh+E5vMGaU4i8jf5j
JXtGSoqtT5LkyLIXYAzeVS3UQ9adJS2lvAZFqOpWINBtMCrhVSEwWU1UNLlzDLK+
95jA7zyWsPtFeg8PSj08wBGiwERDIshnmMYYr+UyuKid/cMn/WcU2GjFpb/eWLNT
QhE7V767JLdbdSB3I5jSHDRGMrXdwJvPZVQr6dKrjji3JFUJqVsbw+gtqbHPTRFg
cIN9XkPcYeIjps8ynYsqpYghA5QzSlVW2i4/gpU+yvUsX+R+t+GIq2tyQ2lUd0GB
UWyCulbB6X8iddNwpkfm6e25BNfIChNIhyYDBPp/fjA6Jyhl3WWloVHuKuF4qKD+
gcg/7+4yzYr5l2gyZwfHEfni8RrdF2llYNIChNAgIGarVLlQPKS35SfXYiZleMEH
gC8XyvpckfPDjYrkGyenbWZl1zlTawAhjP3xWMzlxOWkJjeDmeW04XdI8r74FoMe
oKlxX3X3ji3aUoI30Kik/AIb2YdwWuy/a5+jK7azJqoDBW2UDsTnhcliN+0e6/6F
rH5dByzhd8JnNqk4GOeZAMKf4VxiZtLp47QwO1w2zzSV5riy3Khmx2MXA882FU5y
8t1H5BRRO6xLm7wm+QUrlPv/4dAEFNWJ2RuIuq2M0zZwBvxrRJmyHcG2HncquT+2
N/StR3mA/iMWGl7c+Jo2Vx+i9FaBVwx/PhzdUHlfmbHU2Eik73RCY0KPcymbqx8n
hw7AqmsCQUedNJceQ1+wYLY3ia4wHYpPHF6NSGxwt1ypz3WEySTbqF3YjGerkDS5
BPEKmOwKur6FZ/UIZCt3Lvkb0K4ySemh6q3BCGeZvmKJNOnSZFpE1E13t056xYe4
HRAnsYauHChhNMjWdIXgfvnglM0PaHUzeWoWuG7ecCbXCVu0xyZrn48wkof9UeuM
BgDLgu19YVNEZiyOWqQ1G7TQ2Q3DftQOTFpkj70Rrnq5WdHTdSp2q+rfoHe+aDUb
4Fa6B2iAEWe+0D5eImZM/k/CB2cDCU6lQcUQ4pIFrB+Ai74pgZ5QHOdhzlNnBcab
wSXHRPSXfC82FxzuvevNOEC3dxZeV0BlyprYjkaTMJoWw476DxC6EBO+axHlZ5yl
DpT0j2zDl35Hy3igB31bLG1HIadE6yl2mWF9yW6cydGVQQmmW+2Toncl7fc2zKe0
cWQusU7BaQjM4XPgaKJ6AXO6KttI5LhoH6GdEDBrZstJxvV4lXi/mLGCZKFNtcOs
MRFTTXBICjN3aw3vsvpbCe+jRnRxVY4hbUS3Qq+MrVUxm8m3GAQ38GVIb35wYRTs
Gr6yJ4Qq6FmO5GE/xeKalK0942VK00GYb4Bn6lnAPAF3bWGI0fJkDIpBL//nVpnO
moqlOWr6im6kaPcUhPPLPUToaIC+if5js7djXl9u5XQCPacqUH8CBgQpRHX492XF
VPUSEKzvhSKMJzTcyYydj4XbpI6BLFNIpqEHvcd0J8lj3Qo3SKtVwTORwtYpm8gP
ow9s9yCpzzjd1L0szu9s5+SavdHmjvViOSG0cbVdP0zjHzmstnuzroi8dwd5N2Pl
AmGnawVdtg9WzKvbS5QN5lOovzFcyXjGlDZNQait8AK2O0hhLwovLBcx+lF0Bqoi
/YOzyH1COHUNVgBq9R/YCmm2wG8WklZSiO7fthfbj3hRfugJf8OqEWtJCWjXY72u
0+yvQdxxjNRfcAd16u5Fe/xVYDRyRwXYFkyLOfsaFw8n0Y79v3vPQlOaAONihcwX
wXi88jSpYJk+ZfqbyLbfqKRlaulkl/vHWv7r4dRJmnU4hPy2Apl2h1agQVrOAJf+
/7uPXkOF5nfpQcHeuNc4rBMiCt6yN6qix6rS3X1Iw2xHMJ6KcebwpZnCxkxoJwMx
SAp0nIXGBKAGxujm1AJRkBwXm7i7NPYSJi7G3IZeCQ6nslx4EoUCRMeUxcIhxp0p
XMuD4t0IbiK4AFy/dIk5n+nDjeto32nVqMEM9v+IAy9yWKaluwxzq36A947qc/+b
k4YAu8E8/KWOQkdvrMa4qpCDjPTFW3sEwxFda/7EHt7SYGqhf+p0b2jHTph55Vbb
Nezt7LRe8hKlMxuKgtGDbmoU/BKfOFNXf/M+lSmSmmH0RodCmrHzqR/GiRvAd5gL
aPA3tFqytu5Z+qvFpc/FEXp3krwbFlniSNF0o4UEjl8fPEFq0yquLiPZxvweaU6s
PSkSyf8VRJAlMx/ogAPAGNg4Mft/3lLJd57pyeUWz2mPaep+3GIYVoA3hRhwp095
6O36apl47CdVf8hPW8YmKDVayXlAFzplm56BdgvooCCGNBOX+DRSvKuDopShhn6m
1pNv1ObzYOGOe6e+kFVPn1y6CNB1Yd07HCt4nRe4zcsLRWLoZ8AjkSH+HOkzN7MW
NtryiWHLZkLtxJMIwUfEZ3BLBWjiZ6uenOfHEB2Q+6QnzSuPO0NGNnIMWOJVtxem
0qksGcEIqPwiFkS7yYoyCnC9YMnlpnXtbxSnxj5u+4t+Ny8NGeOwCmTp9YcmXHPj
gNmjmt6K79UlUd9K2dCcGSkn1gx9mFxWTscLiW9zJyzLL62g0TJbu4OeBqVPtigD
IDmYCeFRcEZBNlM1aVPPSqnLHnf9zxM2ZkfUk7a0fk3fRb4GYHqZNNJokLVT4VRP
FEOuX9MKBHVcPEc/G/Wv4fTgXHtinlWBiJUXnGwluzPfysNwiZ+kWP3iCZUqIiFw
vdC45/Fyiis0K7QTKltIfHB09c+mfZNNj+/hylJndHG3QBlxAv3/QUwMD+MT/C6t
Ca/ptqzxVwzgn/UXPwmi48ktRvL6lnzFBmgyxWCIbEV+KMqCdcHG53jRaOMK4TNX
S4yXd/fXwOXoMh3nM5TylwNtzzfCVWogb4yqbQ5tqluiLoNJBLTZnT1WuaxJYt6c
7VzT2hfgT90w/GkzfoeaXewrsFWvOnMuQFsW++90KxI6i1+/fR9g8yczV07hooF+
Q7N2NhWRJiybHkDNaaJh9gbfUQFklXZUrM3T/VUwSvPPojCs/VoDeneg+gzxHafe
Z0ekbIUBO7TxnnpcsB2c6o3Df7TiV4oiHqLgsqESO7tnHB1nfskE92sRpys9dQeu
HZynNT8GQ8yBGMh5REMsYVsX0ge2f0cb22DbB+8Irg64DlBluVRhrfqY+xiMBuJl
Pjr4382OyF0CmAbhn3nRtL5Vx8XXwoHRTUF5+W+sOa07bNm8QCQwO2II1GtqhPzf
DS/jQunfavo12vJAEsYWYKTdkIYXrmW7qWqG0drS6X11vYlIMnunFIj16b8zG333
C/C6ZNA0gRMikJeuLkkcFZHvvYQYocsi6qqz1VnuWw+U5ely6W+16qJApZxEMhHY
DXuJelwcEfsM4vmGqmhZZ8Q3R8Badqq9/rqfohTp8g9jIB1JHMucRC1BoHQKMjev
pvcjYIdsIvO1ht7p4m8dv1I4VCfUvcPmbC+RM50edeXgkwGB3HHRE5KrAC9y7iZM
ha87cREpM6GIY3e28oR/FaNfLq1oeaXxXk5jdV/ytz0+NGBvdznfvCbtbKbRa/r2
s8XnQc2OlZHTRuzJGFWGRHKyKbJ+lxejPt+bnu9JqNwIUgkHFcv0zLdlkAePVM6q
62R5ipRIft7o+FYPQ0eyf+mye52/8jviEwt0nSCZgZ4Op8+liKogeyWABAtVhaPF
e/jYWrmRKa17mdXiBkqGuwTW618fhL3CdZiT9gXWJEtvsJt5HK9q/3vRe+NbuSRb
f4M2nLi8NImgdw0diXsnZ82Rfp9VMB7SjrebDdY7hHAu2tWCYbShOqsaWWMrxkPr
gBqpGogcSAAM9Jcgn9qBzvNurT89JmKLSArRCL82HQDeFDmr6dnguZ0DrKXDFJ5h
iZ/bkUQHp7rZsFESRnXPZ8xEytjD8CE7KssFIRoCA7vjQi+muZFoFpRU3P1rq06L
4Usm495wGME47cnAlCEGjHxeOKzIvXEISL73KRLZX9KvKcoAzBzikBPcVFZ8lPLL
R8UijVpI0RttEVFYGqtz7JyxnfT3IRUZ6xkpwnR9OrQSRsY9CLlVr7UUB/KDULP3
XKuDuBJDL+C4o7jyCU7PIrr/3jfgzxDgzxt4+aIJLkdf4EiXSZajVLDD9lq5vwwA
gpvfc2uopXNRS9NKghdA155AP4GkPfoujmIxvoimU4j7H9rFqWhgsR+DOj8M8VZq
3VCR+ujTiwCRPrPd3XmHDrtcq7CnTB6T3sLyXyl8fvyN3KEg4KHHBo8SXoS2Z7N6
NgrV9nPO1fJ0MxZ5WVWhfrtQmWNoPoABuybM0WyTM+XZjUifOO66EKVukql0ijyR
UYaQcyVHMPrKE9nMcYgSwufoI2+0Cmw7gIFcbqVydQaHkeWThjjbeDdUAbs5ySrK
nKv7B9FvCX5pj2K+lIeFcGhIc/C/RS1/G/95q+8ibvkM+c+rW/HYvVA18hk12xpx
tlhVI6s/O7BVFO1Gf/Blkke79GoXo0seV449nq43XR+984Tad8jUuW6ULk9ugIU3
rm+kFdIcjp+gZ5fqB7ENh9hDzKChG6Z0oNnTcwpx4FADTw9l0q2Cn9RwcM/h6oGh
mBKInveXXF+926tsTx4oOtghVXxF/fCrohOrKcuEyiQNQflfCuVhYjQ9U+1qjsHe
sP+4iwG1NR+se93/O9FjviFwedy7a0+fuPj+akuci58lhlB5wDvzPQbaKHvW4vBg
UzF5A+NUfu1sA9whkJEe6Iluc4yoHQncgsJCNzWiyxyKZr3PNaV8ZtDrmbLeFcr8
E7LB+HvHftCnck45S19sqhf7czINl+2KQoMjUmmjII+UnAfMnEytSI0M4BT9zNmi
yjsi5AXFIQ6uckXXhRXrlZM+RWlRZmvjYDzoiwcRboeVEqczh+u2p8I5Phx85+lk
hmlVP1prExGQ4qX9//xupuuhvKfpYfM8Umfv0hKRRjIhXGKrp5g/A2PuSj8Y3ryT
8Al3xLVag4QwL0QjwVcj+pguVkBGcPcUkVtO+I7fD3cRGTHjREnL+o6nDG9Ah+OE
t30OhuwawpQCOu9oaitmbXMibFlqLwC9EAMrwFTRbdGsUgGDFuHNvkCk+jtsyNax
JTgSIngg4Xnm6thY+k+Yz0uDYOjn3MNvgU+w8KE8VH9da/cokiJrlKyL8pfutBiV
5XCMT1obWmrychJ9auzsC4qxVe6o5IYI8wQJ2unUIaPgJq4HS9zkELg038Rx3OTd
rIfrQoYSisGdQvCNLnViOblxcmXgyKg0DE3paXcXWA9j0wKOyCCAyh0UCdAdESnl
esN4Ml+zwYcJrgLe3C15VLvls+VncSlOudvQrGIudJbLy1qznpa9eeNQ9SkhAvRh
OKT/dIrIvfrHjMeDhuzZnqkz+tsLH/cNlweyPXKd1jwY97ScN//XIyddBs6BNden
uZLYyJa4UGnnBqVoN+ewpAayujYeGoQOrcpuClvf+fJIr/CJVcfBkfMqt2Bs74Be
ErH0vm34cv0wYUE4ScnMLWQ9dfEaJxCEPsUK7HJusPBrtrQfJmnvHDX0Lo080szs
0At0C/mps78JADwdtiaueO+p32RYPcQLaEie4/pX014fAaneBq59ijpG1Iqss/qf
oCpeeSVw7nTPQwx216Suca5JsVbVStYUNoNQprslw/KDjeYpgef3PZXWBB4NAcnk
hNY7nQNz84VnJLKB0x7Vgg8s8SpImj7trzI5IxDjcdG89cho1jrynNtq+fiMXzxv
2Xrsd8D0p5IGLzcauwLMvkAVIdA3+lg/fEKUUf7YtjL+Rr9kx7t5L67xv5gaWRTF
gTQi5D3qd9AozVqzEXl4sWtplQQ/xsOT+HMol+hIoDsWrtrQVtQKyRn69kJo3h0j
kHZToNRaDftOQjNZe1sbqmFqpksbC9ag552eEah/PElRMXc/1lAEYLUCel7bCXhI
yId+RGVmFX/2/qsk0i7G4Cvj+OdnoX1WvTFEFjZn0QKmo97cDlfGA5ieo/x5iUfK
QhDnnkBDS9mHK1Cab+4n4X5ds3Z2oEu+1CwOG0fFleoSNB9tNHOR0IuAoDNlfQtM
Czozqoe4W2M2jVVNFc3n1WztlU+9KSXy+uejli0QM2f8D6RiHVHxizscwhPooioW
rji8NIUo9125Uy6R0X1MREOyz+BTlE0KBqLUdZPUX5TtuOjU2aJbN4Sl2hAXQL1J
cc5glVv71JS3iwkJUrUO6MjQzzITkChsXRRX71of9Mh/yfAKE5DsP8MoaSKpPJWl
L6/+xI4J9FUH29KmKUf3zDrlHz6Lps/+6MzCKRkGTICWgHO98gPH94rRSY1bJP/h
XakwbyfXAHG/MTmXcp0XElp3cga0TsTCWsZfjdfCC9orWZg4uDwTb7Lqv7kyZK4F
DGDQw02nRjLD5Jd+1dNTOQmX7yGvETiQEojt22TOg0bgY1QJsG/sRJEEp0nyPjcv
dLEAoZW78S3GSk8pvs7C3FmXMsk3QqOhV2MQ/+tvkCoX/uD40kuZWpy0lKOHhA3a
YVPee9A/4IwYmKmlcBSDCS++HV3nQDD8/Se7sK4n9vFcInDasVotjxUwaCUuM36G
ahpE8SeqQPsLVJAzNcKlnZBaP5DRiGe4wgQJV2HujZXuyTXsPHHi9N8yTjqkrtDs
C2eZojYL7J2VI96xE7M99o0+CGs269MMww4wC0jeIyrNQ6ViuZ45cQc6mCYkvSeN
BraE90mFoRsUQC6gzbD/2lMkA65zaD8VQxjDBpvOWEQFxv1shqxhVm63aNE+BV1r
mc4dRwU4puuV4+mr7YmAL+tkpMeBF8PL8/1DTFclLitqUouDqaXh+7rZrmW/IIba
2TZwwLlExhYU7DxpTW0b1jY41QQRmxhA4GMJuiSSBVG9XcolxoEcda1AXmOSIGle
EgKrQzJXlxwc67KoxIdTCdKIc5YC0O+0TkqF2JPRa4wZZb73wjOWuC/LJhK4lMeX
EhGbbYGh28Lmf3CiK56dwVmXaduzFIcffVOaI2netHSJ17aIhW2yTyNf+EXQxWiR
6olLhInIoZiAdgpPjr2wvyCvXosKSDKqwcdtifw8fRxB4krwt1a5JMoG8IWNhxMA
okSC0aFasPFYJ42Vf/C0C1Idf0yxV+2Yq17Ka/5tBpUE4hKWGCCQLoeRghgBjMgL
f50tIjZA/VwdK4j1atUlfLg9+rAmHAgBxvWPHl5qx1n51cB4GyI3OtiDBQ6BaneR
iifL+5BHEeh8LcXhLBr9IV0clPrx7em0DsBdjINRn2bQqEi5Fz+Rif8w9rjhxVPb
7uctyFOm2nXY/zemipUqpuGSlLpyxwK/OAWGmLUAfrN4I4HTWvfkh10hNHfUQgXG
DeJ6yc/jhYAJLztHvAmEE2Cs56pxuPMLzwylyQ4DlmCbgQwzw0v1XWQV3tW9/Aeo
/OtZJbb4LlHKkZa/g6avKSgbaEq/AcJJuhaK7jrf3GT6V5GGlO4vaOU4I6xmJgj6
7dpn8m4C3fifehTImUDQwh2iQsIb3Hbjs0S6kLM5XW51GnzZyapGuhHOIo5t3O5Z
N2Mu4vCBwkHI6q19FTLuR5CV3FHsimfVhvKAp2bshbP/zyuKnWpgEiVdWDdwemHu
KJ1/37UGGJ/tMdVKi8ujQsB+c+tYUBz/omjwR4bhccCJYtisJfP08HYpzAUAi0xX
m4uW1o9IN5DWDNyl9VAs1Bg5Z68OMOi31zRg+xJ6c3UeH7tU6gk6Q6H6ELobRyRc
IBw4wf7Y1v+tbMQpAiYdjwAvZ2Pz1LXYBcjZaGrm0o2qLYk4dAwRe4SUJT/8ZnHH
VY+KVXKt+eZlizYCrjCez6FlKsSkoIjAzH9aVd2NvJ0VQVujOMQKLproHwJ2GaVG
XDYOviSbIiRmYO09eI8rccye/YNM7QbgVcSUlZFWeuRM6xBsMZOjmzocjXhjEfkA
rHKOY3tycn2bnMwQ977W22eUqQ+zXwl6A5f9dkGUwAkJyvF3fx3kskAxAHR7adhY
BYMgdD0ZPjwpLZghAJzaYEP6XN9iMvNTMBJrIInWq47xYn+Yt7BGHbgMF1NMUQY7
B94AsREuHa87hhrPM4t4gr68RvZZm03iDupXyWEYxfBddRMnUhUmCkoo91GpSG2w
HS4YwY2X2VFYuW7X+fnHM26L5sCLKln1MwSEEliAQ8sr1blDBek/0MWz23fJ+sBl
3JNvUWSFK2QXmDzJLdHVCzihSQ6WyJbrFs7JDCg4z516xj5AOcElup3QtvN5SJkD
e81ABSnhODV3oY/s7Bl45nKQlMHm+fvTTVbpt7Ic82LySakh3Dqrnkaq4Dry1VVW
3+gJCKiJSOiTZQWW0IugfHYgkP+Z5cjGVN/dbPPjhJTKMEx8crX2QAHhvflebFc3
zUUIsyBNtiQC7Rs8GTnkeh7nvZko7bCdcGCo4Lu+C6XmC6htekwW0qQw+PLwX9i5
RxWJwCv9AyRFV5XJ/YI7wM8sCON6ng1XNcd8chfLH7G3al916Q0k3XuMJxAZRccI
Oi7TtW5aSn8PS3sefhEFiorseLXCaebTw8DQ+x1cBsw2Lcja7i8Am6YFoatYGpui
TapCvuyV8b+nNrSLi2Y04Oge+8gLETTTzMVQF9o5uXjkWBbikta/C2CBZ8eyF5ZG
oUp6sK5HfvGrkb+cyMl1t1sgHkPIa9YAO8TjttFp9+QMg20Y9DOdqaBt2vKJwjJR
ZxdIrMvplgDe6mzDlMstakNZ8QanlZyPEoVuSJOntgUyvgMJEOkaW02kes3FzwgR
wDVw1xwJ2H1lSrvI9CwcIiqx5k5TCiRVdGDog3Vk4/UoFYtithJ+7RRcTw+7U0Fm
pLGo6OaIXbpfXdgZyF2tHTAzeNYrv5vACS1qgtjAlvnQTXPeYveum5XRXH2rN60C
BldZEYPwSO7/4Kls78tvGZH2ebewchACwKNYU6HmW4Br9m8TLFZlXL/qerz3+mdz
GXYhb/G8dl27two/X06tajKc6Yc6ttDflWBj0Bx+VeQ+/PPMIbdVZsSsSWYccwXt
1eJ4ZMHMgbpHdCLPbDyuRrJtgJvA13a7gJMolzy9TV3DFOwn6NunNT4HKaV7VL/8
dwL/woIaGb2PqfGsgP/cY+hAJPmSpYEd+w0GfG4yXaulsBCCEQHTUmz+k5YLPW6C
LfLtWclF/unMrHiIG3/L6egOLXebsIt0331vhTe9a/N7QUiQiIayjwS3rJwTBpRS
w7q16EEDO0V8T6iYQ3pHeGr2gvaeJyK+lrPta7mCvFfp9qlsTjhWGUVednGZZjEM
QAbvcBQbjGB8n5pdMjXSbrLdBSnOeWymRjqvY06GsyO2z+gEx4qTGXplWAaxUSXD
CZN62fSdMOGg3ls+RVqkl0Lf/mEXKrQyHzKZl0yAOV730nQvVRIWl7L3P3mmBVYP
9XCwLEfO8Do9j+O8Ov5iXm59mEnYcFoJqI4FIoZVgN1oTYQ+rvXxxoj+KSAtNGdp
fl2BYpAEktnv4V7RB03jezmRHnca3JhxKXKUzG0TmB0uNJzrl5WjUJiPh0/rEKHc
ccudFfKaqiNpiS92eGf8IAkFoAwAckz/rYgRSL0tddbusBlRH+5yNH3VCatVjgYJ
0Q3DFiGc5h9vcsU3Ii9QcoQ0sR55bIBIt7JcCJwL4nQ8Soe+L6xIJA41EYBJkUHv
ryAh/0+xYUzskYuKdeAl3JKv3uLF/vM5x54nEF2Tjtf2QKid96/K0jMIw2/qgxT2
dkJCyZyclpIB8yr4lA+Ct5LOuzKirB5x72kVVAjnP1ahHpHOYZbghOSR/hQdunqC
UUK/jGSJJ9e+N2h0/9rra4v5PGrFGndy0pRahNMsN5E7VuPMKnrteESzWKqODat+
dV03rtb3Li/l+XRXKnooaC90iGC38Z+tyb12YYZs9wI9i/rQDZT/f2hxK4+atrdF
GpSbA5IVgCpb8PpWEpOiXqXG/6UHoLd/LYwgYWGCkOHWZZOsgE/9mO27Y4ijEd/3
Hn+Y6fe1VirUiTQrFdptib71WwPIKjxGfliLAkKIlwAF9iSmK6PjhWbfmuicVXEo
o55Q0FaiIwKXFzAylRjgU076bHvjqArBFkzKZ7LhVVvbV5DO3w94Xev0cq8LxcQP
C/rfV5vEHVaDA3Xrao1QYidcDukHSmkTueRMJeSSIlQ5CzOmkEkxTbCM060pGZE2
f01Xc/PLiS2DIP8CqwsHBfcS3zLLVs6cBxIb2LNl+QbHi2hQRVBb5QFTdPfZ4z4B
lD72HMLlzWp+j44Ek5jAovAZWG/rSGZtbjDpUHZDwF/HV5hW9keRBdkN2d2hSnqI
7K6ZrQpZccejr129CE3N06LUoKwSKbz4BznGcz2y/O9XNDv+9EfOt/nbUMWaunr8
qjjkw6rpH+14WkrJoK5rwkRTGE3+xBAfy5KT5jZDfPUpSX6gAPJWwyLQ1q4dTYxo
wrjNIzOo+FlXRtmXgeb1lZVg9A9xd8MmAmDPBKNkLiAqMFHn2+/HRgh0zmlKFFyw
sHfdF2ZfHG79zgjxtHVzHYQahA6/XZJBg7hp4w5Fn+lvnj4YO/3d2qSKr5Zl80NF
00geD9ubYStKkUvpgoonHJEpAHqCym6q/Gb2gLwAd3hNimQ+ykj1oIhsA8Jbqbfp
e5QGh+Dl+hEGXjEA45ih12BGXQ3HmMuKxsSzlkUKg4mGlmG2FnCw28VsPbEW2/xi
quuriTLgZA48ukdedj5uJe0nGBb1xYb1IT9STUFD9YvBNIONl9IhCb8yolOWbgDO
mzHfEq2ZTzH7SjkRU1Uxhzr98gKfHWogU4Nbflkj0+CIcWOAGq4f22zlPyncWLYx
LG1vrSlSsMRn2BdCXyKfM1ZJWGeEUv0ChObx969rBtQTbSmGq0EYGell8GfrilOG
r3zUU4hcEQI0qYNFXg5JEaPf1diJ+P8tWDoP+dPYeSc0K1aXU8q90hk0V1doQdGt
oh2zErT8J1zTjBFdzRzbl7EKM85T02hAmK8LOEPTavTJBNEgmiE6m4BK6EFWEnAG
Ka6KZoEN0uKqJWxSdSx4DhUYPEYQBjl/J+ratSEf7cKEQZafhUMVe2LPBrluYMqN
r7jX5dSXkyME1kH0SDsSDYUF5MD0A/KwwfTMIEOSbaXH4f1MD5RlS4AlQTfj21CS
e2dYvXY97xnhtRH/QDzn/w7SJ6gdgcSs/hs2V+ZSHUvT0knyt7zVMjVBnXrCuPnX
RjZi7AmsI/Jm16vdSHEsBYEcfMXkT7mtelWm9CIVbDxhkYv/U+N5xUpjfE0wp+qF
B/oFUdVkFsmRWK3iBKVs9bvGexxT0I+UWyAv/9JRJleGAGVrtPd1Pov+j13AFrx4
9b72ZWpTQue2McfEECdjfEgRuS09nMqiE/f13IkknCehB7Kq06K2aIUk/7HSq9DY
0xIsOWSd0s7o5PiXcGMykWIFIFUhWLZw8RfIiG4oI3Kp+YZ/Ta7+hKW/fe4NXDPH
OcaPTBj+nb/Dix47ebhd4JKtHPpbyJ14p8x+Pxi7i79JGJPdl/3SiawnVcrAqjqd
tUhm5ynVA3tBs/DPC+FQTVfWUaEDVCXRvWx5H8hV21eYDjB0x6hJjRuyZUV0ubGG
gyTY50D21PX+iy6Hr+SGyV28IPslQbZw2bUIwnqebl0pKXo5c4IotdzBi77maRrw
pgTkiGkbxWnZzbZLSmlFAUpMBU44VpJUmmW7ElCNzBkLOr2AebE6NeUJJXqo+A0t
yQE/U0hzXpiuv92dlXzZ3aaDE40jBgfRfphdrLeUpKuBdldT8Od5rccHdx14WBng
mfbmT/IhTB3FljkCcAhk02hjaMUcOCZZxJ/8RLa4Yn2C9Q354cSYjYhT9HCakO0E
XRZ7OqnOfkp8XBRCr5uqrapxYJ4F+SN04LqxypaX5tpC4c/0mPHjhLOinWemol5I
SSCTVnNLd0PK+cSgzUd5Ktbr1Xd+ehknkRIxjSsi93W1JjjgV9fw5ip6h0y8UIgl
0Hfb1QPFARifcY/0udwl6N6v/ENnvKXvuIzyD8TbN/xAJionx2UIYDSTuMrmzCgH
5KteXsW2ttfK4R3bOav7NMGX42nY+ETpHy/W7g4PyYKYGHiQywBujndQx95QZhCY
fmI/0KZziWgZmtd5hxgJRy0dL8dbYGx0oXL5e0YaFdEctSh7IGRDv13w1qgifXY0
Hi3oHFyvF6dsc0Dh9O1hAPEWbjwZkv+LgnmYo+ysLmVn/6h+TMMvHVTHIIBjKaxM
DtkLozSvhVLddzDZorZu2hvuv2oo7cCd8lxhA3vq5HHFWOSmTP1uaK30pPdA8am7
5EIsOKQDkLHLfAlczOCArTXgQswf79qH33Gkk49lgAwh6T85gBbpzQPj1v92cT8q
ONUShMxKDT1+E6dGk32z6RcpHMpaYCejpcFGSKXikfPPDieBMEEYl+c1EPzho4Q/
AnRfAylN/cMAIObR+Z1cbQoaCisRW+ZCkDMx9pCqmqe0qbzEstcW52it2uEpjbPK
cKOfBOdRcRNCD6vhGXXNoqIsV73pDlm87dVYhVpK2AQHn4hi6ArIcuNfKlWQniQg
k8psRdljPQ/vJKibNYfIzhOVxSwOfystosgulJ8LMMPUwXsoSo2Em6jQCnS1riNu
sH/pe3SPfyI7wQTt0yynyWkLGkVH/RO8KtLNvPoc2j2yHU8wUV/i/iUMHuwqmQYj
/aLv5ypDKSkFRy9/L1bAEy1KJqIRVOTnqsyP6zju5ySM6zTmPpnO88moPm9IS7cz
tCYCjMi0Ey8P5z0U3Yb4BGRPEKRbXXAgffbpXEY/o0+xnSokWumiEnTRdKEJKlcE
IAkXHtovwp5WOOu0fGEoHXwv8AuzR0307CqoycF6GltM6Wh1lnS5Xkd/oXl8O6yt
JfrD8DfCl5WrLO7sb8+bgNNeH8K7mo/XCXaIXQCimBeqEBKkopgYM255JPZBVCQP
ni+CALL0L+eYxyJJmH0Pu1lZRa2+MSskYZEh9zWFrx8eFHlgc5KZdtxqIZCIpOPm
QnCf10QhiKhKyH9pVIxNjA8nntOrA7yTpLZmm/apfDDVcYCSTBzgdUdKaKhHUhWW
AUexyg8B+xl08QpdUAvK3cTVjj+1M2qzegV2Q+8lPLkcGE+ZYenQJpVe/WCi8EUr
9FwA2D1sq0K4N8qw8qmofS1+f34mp/UXrmbhizcxAzaRvveO+Fq1ldp3fTr31ccx
3X2UgtrQ1sEqyDlUQhtpCwMT5XD2IBZGb8PelRSD/iNYqY+ABgu+9lxADlyCyH++
dG6kF3+gQKmu9cwpLnBm8AK9Vsg8FjpEJyTWp8IPAnqMR3l1TiMsay6JeLyjsbu6
PqQ5UPwAjDiAccmsdYUTbjLyn2ayXzVee1lyqbukdy1Tje5yj5NDqgOoNmIwJmFK
7pQkiABC4wBTFV5A8RdSUDe3p5+fucWri0kxH1I+86JPVVqcr/PVK2SFWoEAu0NL
zDEzTRWSLwlqrbGPXP0hvt01Dajc2ug0jYZKfGecXVJENXS7V+N0T1fHJiC0SNgl
6g3XUEOBKNSvzFunNLic9R0oiXZPHV8VKiaAoVNlOvDqIayo0A2fBasSBH+vtXlm
Q5vuUka9LXqASTaVRXuGTSm9mT4417M1skqfvkppEDvbpJplGK/TyVVPfU5kfegQ
KIs0uhEhKrNVy70I+AEJgwzFEpZc4/6UUUDEVun6AEsDm/ls7Y9ydhi2MvHejsCp
otJ+jyGV0f2C9moEgh3EbDzq553OTNNEW1P/ocwyCfOTVCE2UbXpOrcnqWofEG2R
m41srqYcItC4lJt+QacVs/haYdsLMQ7jR3Jgr9LK8uRkD9tzqD0Q0+8Rw+AanXrO
EoK08/n/9QUpa+cyh3LK3JPrksi5ANrRk0QYZzf9p7rj8E9F8OdB0xL5pgpMTtqe
E+9g9p7Zx/wAQfWnLyILlrD/cz0e2i+Ajl+DJ6AHS2p7hAEiJRhjawBh9Ok6gKlB
NgZKn4tpv2Tkct9ecmsIUP3B5PdA5t4c+gK19bEUKeiFdgIxyumDLFWdqte48VfA
NnvmV9UCpExACou0eD7WtT3ubdRC6aSnmIeO2qT7GFC6/gc5uwEFWHh9dEYXlm5b
7bfWIsS9gXvR/KlunA16vIvVPTurXZiFRCnTBfUcyCfc+vpoSKyzD4k1nEF3zR7U
bt3oEMJnLqaBzSQfMGxLVcsQ2mcA0y1gpcwvH5vOGuXWOGDGcUZal4d47AW1K8RF
SsyQLnqrv1QsKndgzjy+iuimYVWmS3D/GSeBB6jUe9V7sYlWRN0E1r7ZztWaEIc3
n2rYANf7suzrH0kmhTwchCGQcEcrpru40RlBCXRcEBEKToqrMKY2S87r9dlAXB1H
iUAUg0kiBmoPXcManJetIHkD1U6Wgak31ffMSIyeYN3AjvN0e/uyrAJRHQCAnTf/
vHrYL4ascEbGC7k+FjAzrp6VXVeHMqRb56Kw2GVN7Ligst9Cg9XoO+NDjYtxE9e5
8eEjNovAQKjhNn/r09Tdi17ugztjNLWoVImmrDLwuXvIAjgRzU60P+JJP7Ir03Lt
awNJzYe/Oz6QSIHOBSHfUJZ5RvWIbcRFja8n/SlAT1RuGCaHckhEyjdv2p6Zh4S2
z8O21dM56unpd4lyb3Hp1DTmOe8H5uBIJ/6WRCFNtie+gFuJHoILEJwok8MxcAwj
VGT3rgzac9GRVtBAPRz/lY1Moa+iHgNlfoeAccNGKwnHiV0YJwoyEaRu6LFZoyDx
YwJrBEpg2ORwktPv9eLtFGwOndDu2P+ckKc2ogYR3ohTIpl+1Ge1qPW0JJ3Kw6EW
gS647HA0SLWuBa4slUFjUzKITNQLLG9GF+xYVq6lFCeocaYlGMhAw7oMI5aizgSA
dPin/GnkfWGmVOwvUtaMbdoA3EUK9MRyvLKoumBNfHEQ0TuKEFtMc74NrPPCVe1D
i7KZcsvoEKrkIZCB7ht0psNNDwtiobBSekihbwb0h9NYEi5pGU6RNskTpfnnfHqZ
SEe/13uE5n/eMumC/hv/D7FS7HqfbSkS3VzsGnlZCenw2ghvoGS7Uq6WHpgWJDI2
6ia/eQCRjWa0WS3vNyck3OCiReX6STrbDaTj3K0tO4hg0LgPJUq+IiccONH6uqjQ
D3H7voW7M9mxfztqjuRJATBJM8nVyKOMfEEeApaWSJ7XywO3gIHvk+haV/6LKOyv
dxsahWSmuM8WtYSVwRWQZ+ixC6KneXCcDhSROtugdrZ/Pt7JtUSQXvBuymrNxakj
8lDjNVOTCtc/aIdhTP0myCU+xzXFHSgewiX/WbcwUDDnuv/OT4DnQxIBQy+51E7+
FMX2JURnuk1HkBbT4w2MqBaSH0tb+GSyAgHZUXOAYINGqHDX4e6iVdyPlJOOl8HV
Fp7dyUwyS4TGZr+XaTajNizgV3G7BU7HE2kKNgZCua7xRdwRcJVrkcCggWMwTM4H
UqVirraSd4eMirIxzY4OqM9NME0brrvHjhfYXOJ7UxSD1IgkKyXmwwXrMueT+vYx
ZvhTUl6oh7GFiDXXHmU/d/CjKAUleUgkhfUuM8JeLEtaFdHE8piAu9bFBOg/lwXm
pc3Qsv5lMf4KHteGUhqgHEJopNNtfm3Ycv97aMj3x8R8HBiFnqhEqnUr7edhjYEK
IV5rYIX8PDUBOFewR09u4PorLc6DFRu5S2+AGSNzB7pTBD1vPGQwVizfsQLCiXcN
yZ54u82pUj/B5dzl9Ibn5puPSb0UsIctBMRLDHSpnKAKUQJDHYaAIOLwa+SMXBEh
Sydk621B88lNxlg6rf/fmDtfVakJ2w1c8VYm/i43SnHg7tEHRLg22shyBoNB8Lx3
Cn0gQS0gTO7W78D4rhVH1IvnJmcQ3mbFyxmoMCCw9j2LLmD8k0O7q6e02vV+ZSf9
kjaH8UoHexby0K49Z+JuVS9iWhv3BESECWeboCHL3W+sm9m7K+yStGxtAu0NZDa4
xnlYr8IQ9H9BjqDuLeOTKfmELF2bj9O3Zktb55YjOJINbsEeA2Zhv0NF0f9t9XXu
1SRxwadcsL+lwHcdg3/k2L49iYTEgbAaR8WzZv0VoRS5h+ZoymH1cYq0QHQY5/8n
v1p3aFSvqLCoQWVpPP+M8RYEkWiYXzouuCRRj8ZPmgC/nC4BpJckvmiHdUrks6PJ
JZB8u5t6tKOtDNYDBNmH+2GcFcn2X8lJbg6SkvnB5997JVB0ENvCQsqQemsJSb4z
kkOnuczRCWIfSo/qTks/A+Y3opf+sKsI3fofuypEJM3j4eR9JWEMjR4WRk7XB7hA
bVd5wQc1pDQPe4a3WDbk4wxBGOVyRaxRm3MaLD9airDMI5rohFp4bBUANunypimc
892nOf35Dsl8BPC1elCpixh7nw6q22nov7JavFJS2iQ26Xjlz8Mk7p9B6s77nVjw
oX3Gb2IA3ZGOX3mizU80liT+K5KMlbuhA2eRTan64HrwgbuIueB+R7zxbi2GSexh
qbLmYK0pz7lQYqQ7qN1wVeG/uvAwNTgR6jh9iPKoEm1TaCJU7htO7Il90FBu8/+y
qS92I5DgwvhQLTZszr59h0CH2mjdXddCOjylKmgPWavqHbrZpbndmPRpRWaPyNt9
hXs+Z+3bfruP5vdZozgTiG2hhGrMxt2avW80WJNEwbCKMLXLpUwBJ7OvsHwhGBnR
zQ51RkQoIbXVPtGLnylQnxkhrUM9KHeP9Lx6/dufXl5StsOyouBeIcN/32BzmU2R
slJpUisi8ia9dM5ZC6c/ArbNaWnikLv2YnrZ2oMnN/BtpdDrCzCjDyXOGL1AdBsR
z6GhSFcM4EIJx4cUBaWAwC8zc3Mt+xaHwdoyMWj7YCk8JjPHb0A+5LyuCHCB/WZN
mEbIx2Pdxi4ZJ77Z+HRbD5aYTPtJ9iSzbDmomm/FmzsjjSO9JtPgwSXkRupqk5kI
TACLaWm73VpxewJk36vU1EZwb110y/iCkhBNMWlNcL2nOHGxDI5Gx+YycgAoG5Me
el3jFp2bSgE1aiU9ICITa//xmAeAr0Ipq9Z1QzrqyLlGEq166i54/5BOuTDgdgMR
5V38CdSDt+D33hsf1MM7qGQUyc24DMD8ztS2r7lgdrwb7oF7vmYAQXW22xUhqXJ8
rYu299rsfBBa+cwtcb1vkqMxK2eYfHxjzi/8Vu3J1PGNZCVWnLYEFeNcwGwlqV65
a6IiRfZFICUevEWYtHkqL9P6WzWdvSTAZoT2skw46uw6XCPqp+m9tqzpsKYxXFEr
IbR1kENdgIMXjcPrx7aVcOJtXhRUCEGDImjdh5Fi/KpbFp+O+FcGsp3skjVOFE8f
GrHdbJNzjjO52ZUOpmSOAh+rHeOloOiNZ5Zys79FBDsIA1jQ6CqDm5OomOvl96XK
EZq0bL2DQZVVFeJeJXog2G9qHKi4NJf0Nq3+lUIdSt4AdAEdBaGy+UWkhyMoRla+
8lQapq2v8SD6ovQowte4YoRfjRXPHxmaqQn8zv/1EtNuSwXTQK0RuG69q8A1Jgzi
vOFJwzQ+fxB6ACPFs42AkJkMRx+yDsLPOeE8vJVAIjADZ4Tde53gdEU3Tr+lXdQY
6dPdjUFhUQX4TCo4xTqIWQSUulJbzCS7sKu1+ZY1uveWY7YNHJNBaglNT1/H8vX7
1Cx+w5VZVX/VeRJXcZIEtlzSeO5/4KyZltsJ23Llchwovvn4wpIuokHrupOn+SHB
CQr+2rzlyFNdKI0R4uDSyhdvId2Z7ATSmGx+/RockSDAM3+SsI3VvjshKIfCADU6
t09b5p6CV66Wa9ioBbGRHgvI2Pu/8vKildPmiNpKZ9SCzsLvpVzhREDUlzFZGUUD
nR9rzTGk6EO/1pEwitetPlpFCFVAksAITIRiPPzmRpm46dYzLzRn7l9AGqwNVpLh
cbjF2Bw50l9xHZ5raPkg4fgdZ87o3KdesFYsNvrr4R6I7RovJn1vXZCaxORDX/10
Uqeanlm9U5ac3boUB3leehmtAYrLoVVMn0WZpbhJNR2N9UW5lDhHoV9w02y2fFP0
MOsPM517WEwWXInzbLa4//Fbcx+NnjU4xU6rHo3PkTLuPgnzKCBtwIzWIx+JXEoh
RlMaUe6tB1aqjYdgcgH6K33+btZmJcwIQ0ZMAhP0EqNt3aO7gwsocvJnRIQpsxKb
JxI/IDMrTnYmZpn9ptB1+FEjPS+gwXmhgwCyZabKLLdqzaJ/Y2lKXc6GiCP4pL0x
NoWQEQdRS1XWYtEDm06x1TEMu3D/kQwh4vHvo+NY7kJzUIjAYQo15uDhJUc63yik
g3Gps1+0De48rlJ38YgzCyeWYXQ1ad6ZXy5M1UhvVIMwD/oASvPwZkJTvWId7fX/
qEqNxYKj9dmWS7xikpsKLdvjgWCvo7ECJBeAWrG2Y8iPlP0tux8f7QpDdEb1g6O2
sWTkEPVM+1vpJ+1hbkqxqHv5m4I6inHBREGq+ffRooZjUdxazqUP9Wwa480PF+j6
s6tlYUXiTW1CkUutwYHC23KGgDmRK4Izzfp0cYMYfI57ncfVQSfLpCWzHs9IlKd5
AB5H9rBjdY+uvaNA52GaXvC4GSlXDDk8hebbHqWeEcdW25WLoy5ggb3xDJ3JPyH5
6BtLtH1J9kZsQ9AImtUVxZ44PQurtdYdr7X/yl8alAzwaSNdL2p01Fff40u3PhUY
OoWxSaw7EINVFtiedmDRdPmoFwLfnSSzvlGpr1bb7xBW1l9da8GZT6eWMMjAxlTC
B5CYbNuVueu3HfVxduAkRr8zEL1s0cSFIxA5f40kVanmD7ccT3bDGvJcsoSmYCKH
wa2/7KIFB+SDQhBjW3vKNQcF3wGTsVjKdM63VPxADH1vpK651PD+LFzGK6bZbcqj
cgfYO612iP/DJpnFPBXNhf+4kiR19rUXuRS3Xby+4dUWrEkw1lqtvcW8Tldeij1h
9F98B2Vwh7L7q/xne6+gI0h5RXCzuah9ndkWuPoSrPpOls3v7gcNwZZqGNPohop2
0uAcx4UP5heYXwG6KMOChC7SuIlBAOPXPT+px4vUJx7AmgEi0iM4Zn2gnM+KZ7TD
j3ByrWah9NrHouD6jqUPM7ZV9SARRNNIdr3Le+G4tiD0jsuYg29d+H+FGK5EW9Dx
OxB+C8C669pwPm1q6FRravKhZEDByoeeqhDgWIDtFleNt6Mh6GoPJ0p7rZndGmyU
zaKVFUq4Fep+3AZ9ubVfwpP3hXk+nNFCi5Ip8ObgRoQZd0abUBCdQav4OufgoPvQ
tT2JEl7Gmu2VEPzc74tJfF24PEf5Bb7usYSLpyNJ16DSqT2Ynz1HeqYvN47uoymf
Njjg56lMHeKLbdU+RkhUm7LG5o1jrW8/z02EOQigYtJ6v3n0UtQjAm+kMPZGJeWL
HVMma7Omnx156F724XFTbCQ3A+h0wV26djVpZLRFehJlPcenQ/3qMtpm16i3tW5D
zvpr9VqsRSUC5a7vUkifWqsudKT6M2TYvrl/p/gjU1nSEeG+6pKSXFqahrF/i46m
cT0npsmPSKg6lXWsazVs+moIH9Q4epE4KQdOVIpJl3TF5jswF4rz6aqaVk4SkvCy
ys3aXVbP6ql1qB7vpcqXqnVjjJX4fLo0SrtxXe0xnTF9LHXEQgxk8ts3Sht8MEM5
o59P1hEH4jYSRNl2uk5tx3Td1BZQlBELtiyFqskPoqbO08d5vDP7HhLLz70wq8ET
OPzqqjBlJsmKk8Z+/4zapvnr1g4lNndsK7Hz5ojdH/nKRRjbN/7iocjDyhZu1254
yBGPZCWMT7n8u2y7DHng2qreqAsTi0u1BQdVW4BcNF4E2iOb+S2+mUtNSlZzBI4g
H9qHfNE9YH46SY+lQBk3serbxNOO5BmgmBNxG4zLoNCkh6RGiDhSjBBOarf6uSSk
qwYWlrFWeMfOPQNkCG5FyuRlFyClV2ZRayvA4voe01UgEk6qa48yPCy6gGiQpZEp
DG9ioIGVoU06Vhs8zbluRFOXj+raQUPjvUwNLchmHzM85Rh079L/36wzAIegwd63
b3O48JsRkcnKg8RSGStS9/b7Oz2tFTUqlO5eD4xffO21wPFNT5j1asilvhQchDw7
ohOzjIeJCpoJFJ3uqE2/EIV8rSZFGdxG2HCObtmasllpbA0N+2q+oXPEexLfd7MG
QZIGRvOlO0y8hktqwit5DYL99clSB66A9ELeJfrd4f46rENT4Ghdzl9AAIBQA+nT
2dUVwjBs+2NvqBl8amSIOBua6L3oIm+qMYe8o/2XDi93dkeL1HHFdiSaJjqPvIAo
p8hEm+X1zvetg06qONv7NDVQTwE2SpCXpPUgQBpE2IrH+Ww+7EiEu82dzsPRsb/4
M6RJ/sWCQu2vbcP6P3Ixhcy9V0tIZlURKZOs1gnhIkEkuQPeqNreK3SJ5VtqYMQx
FX/7SlAQmoRE+zhaP3Cuelxr9fDYhPNLmnwr0mBYFataUC+hyu8TiDsU+5qBIzLj
qu3/onS5wp4h13BSDh4m+02J2WKDkB5Zp5vi/PrBqpL1CZgyhlmhPAjdd/bJgg7W
IdsMqmZ2MjqUwt4vsiEUeX2/0CvW3sG1iT+Eoigob1owXhMcVmotJ8t8BCggEifZ
xea6pCTeC1RyKc4v9lIsPPRbONJFGbtiLnFZII6SndQI3IvTBB/6l2J7VmuYdCqN
3R3dePo3m1ZV9uCcay8s/6fBXT3EamiGlb1jFKn6xt9zizbRVU6FtNDWnlvRbmYl
hACe4XGuoxe7/yWbQLJp53E/A0LeOk82oDXlFBY9kvtesd9pgmImV7WU8KPvkljn
9IpORQ73q2YxAEtx+V6dGIcGdqtNIRX++O6IolQsYH9UfDk9fAjuPOD9tBYpEvR3
daiMZP5S9vFFpcS9rz2hGHroecHlb00nweDPxUiENDDM2KCi5jWDHfiOAuQ0s04M
PwRtL5Eur8yLHhdUv4M63V/67Vd7IrLrt5v8C+Ly9b3lmxKQFmaMemnwcrOD0U6B
HZZw0cBAsAIt1nowomt4Ty6ZDx6f1Myr+jMyrOIrwBtVKd84P+agO14irUGsVfss
Pgbbl5j7bKBiz5FaaLoT0tYLIdqjAazd3w/BcaX7XcW9QrWYWq0eG3kGQq7KHKse
Dtq6qhHU7gpGtOjyNHl6SknisnieWPZHCjTCzeUsoPynjNJ/UF+IdrQAXFIDdRnQ
CZGytxpvOI2GIwR+zxTta7ZPKCeMyUMt6FSAIBhp/AkEHd5nfLC83LKza6ZLT8gQ
3enUWPVkuyHE6u1UFQBnkcrDkS750VV5kDNezWsdcLhMtSXtpxEROtljzh1ZUm/9
a1r7KFYzGFEgI6zviUjycKYlcLuDjKG8uhSN+GS6Ny+RiqhmLwBGlZHdB3YbLJMc
3hYteucY456gT5YebgG9yybI56pWV+ijDkcr+s1ng6NJy72VzOXfgmrJZdybkWUt
EGElyb0eJ8WBrFIKB5hz5mrrVFNvKPePXVqmi/QDtJ7xbpXZRaEQXOj9TmNcGiaH
5VzhN6oKKvtY0qxuzb0wPaqfB/Bw7WHaBFfn0+3YDoPOVo0uLSpc1ehepfJ1ANdc
slsAWTIZKT+eVB30pnTzWY5HRlNWhmUA9ZQfakMx+z48HUnSAsBNy8C4E1T4j/D2
SffRh3PXT4XlCsSvf3QCtIo8909oQNZaQj6+xtNfvXgd20ton5iDp9/b4bRjmk62
NBVJZzls5SR1p1ledppuEf+jJxxEKu34rrBJdQN0m9gxWqCteQYKPaWDZuzAo9JG
pmYzloZkp5z9pKbVldoTSMyYLpxPHTeatp87qt779VF2fUAl+GVU2Sy3ojhbiwFo
ZcXftAmwgCnVBYWXxOJ7pn8ZQNct8zhzrvHeMio1Y43kkkKjofD3HyWlx6Pqhi2i
29YiDMN2yN6cffRXYX06DLDXO2zW1jqEBdelYGGCKw9nPni7GfBtALb6ny5jQEVd
JFObssNBjrY7NY8tcjBascBMTeiFwY6yzXLhMtFvG39JIMlTwFIZybwpvBJeHb+7
sch+Eog0GmXxQ0d0NARnCefTphlyzoQmjbieM9Lk28vpUvHKG4aCFJhRxqg5/cER
TAgdqMkWbZMhka6va2CTSRZfpjjaXqQ3W8X7Ke99T8hn0Zinc0Opy+USjoo25/Nr
V7twY98XF6fyGMjH8YKUTnQYddKdrqKKEtqRLCO0r784DanvhOT1HT50z9sI3USa
V1+w6hImYQ9n2/Dw3I9J8vMtQIebpom8XKiVDZ0r7rnaSnIw7llhsniOh/jJ0aMc
CURu1WFUHLOd0XK+MsDu4ndHLkB6GU2d1vb2hFjfb98Z/Wb3nW5rCM3/v1PG/wZG
C9R6yA7xoGvngUngNd5DLMxlGA/h84G5ARavpxtJ3IF88nuuLCkwC9IUxZWylrJh
MkElv33FbfqZiJl1ufcRwDA2Z69rdQovnlpedNaBkcFYzcZiA3McL5UIe1j2IOM1
DMiXqaZwX3JPIFSLWnWjsio5/ro1NRRIfutO0K+INFkHvrJp1MhkkwhA0BZ7RwyQ
QB6Up01X38gA0vmVtuH/W7YKOidT4qV7Jqf4yYcNwhUu+B9aOVOGBrcvTIMH3hb4
P/kCsjmkh5g0l9BTyQQqxGX0KqBiJ+6CTS8hormbieBZlXM5k0FkWWtiYJl2hoxo
c7iAE9DdyVKPdrX/QCxUg2PVHe0F52QSxuRis+gtGLIRVlrD31CprdUWPw7uXX+F
hMg6RTP8U5Gk6BsFA/JZW9ZkPbaOjJe0pcDvuS7hMygwyZ8Cex4tYo+Fw6Va8eLd
2NquzgTyzDOZiV8pi1Z7SDKMPPQaKD2nGhN0jy4zoaZ3Vq6JEUjG/fFijQAwa7T2
YTpJZRwQxsIZmPXQz5RXzkSPh5tYZYQWIg3Gp4I184w7vtZbXbHDcoPPEtEhKt/n
FEdHzN7fasDglbUBMP0l2TzY4pxymMtZZc6msZ+ErHz8dbm5p09f0clBswcz5A2Q
5utcsXT/yi5SrO7QLxsy/orJZw1j2/gRrREgSA4pt74u8+Pgl2z27/dVg14tq/EV
TqgpFIW03Dg9oRtBFSTa2gCDKQNrim7EV0ofuUS3Pg6ZaPREvLO8smxLwBMGy22h
i4LKSr0nriQRQQlFOrkeQmt5HlsYPYBA0XVsMrBX8p4coDan93OZm8uWnuHvMYmd
Hpu47QGtIrbqvtNhYJ46ta1gEuAmmlU8tpEynz+iagFn+tJjruA6OYBCyuCk4WTu
4Dw7jcOS9kJBniikETG5aZy6lC7CJdVd2u2oxp6J1OHtzwfq3yYUV/VyeUNkMKuE
/ySZnJ3b3p70RzhMKaaUgyT7BxaibFORryPYScBBhjsqOjp3YJiEpZtCcznu9WTB
gLK2wGISW11+8z4jy0GoeeHh0nWVSmOFhXXDoegmj6J+nN++7JaAz2WDcMIBvdmJ
bj8qlSCLVwacd1NbDnXR6ExNbf0z3ziGBaMnWHE0xPmyyHVzIVxW2bGPPikIzqBt
fMIRNu2kbNmbLsSV8uLaKp4o/pDW3NMNvF8Gyr2wtIrPZSTSMEcsB3ywwcZC7gDY
zzJFVLNbG1cN52vaai7JJ8G1EkE2HMcrpp3RIAl70a8CDRjx27aHrw5n13zrRyTi
PVZQnPp1CbDwOTNO7/AtoRzTivU0w8VD8C+Mq73pxx2H70CndqWY3CalOlLmbVCw
ThA/IZUH7zq3yRlN49CZEUus+uupxppIHGNLkiitT/r8ahLZACPYH8W16o0Z75ST
Pxg+Bv7axnxaRSAag8pkjH5EkBbHzAWDthZwhpmBTG0YdkY4JFW6nlcj66YOsKQL
SvnQtkudill9xnaKTyhy6mdk33s5HR9QDq4/TH0d0O4fzA2uBinD7bfAL0Ls+Jt0
Gr85SkzX5oke6ib92m0RRurm1zAAe/4VpMuVSVNtPkl85sAKSdk/D3uNjpJUU19H
bJu3Vi6NUUbY/7MCluiuIQxllB6o5gdNH3Q833jbQyCHBnhL4TTCrfN2RlCatn6x
tWhogRnbaupW6I4073D3TG0i6U7p7hSRTzQO/kh+AZcIQ57NHVwPVvOMjyZ95hAC
MXWChbCN9FqmsC+sVd4lWCZsYF7MOP5UfCvxN5e25QhWsEyyI52b+JC3Jb36UqWH
viZCLZtHrZRiMaGROzWcgGZrKZXSalbWQ3pB+6EU9W4tq3J7L7bfCvAUOlNSpFuS
76mhA0LIAVzpUt35pDeDeIZWyJ1tfisre8gmXm3t1KvXrgR4qiNgh8jtTGzIgCMU
PLQYz9tXCsbNupexcOQQi/Ah2FDOc5ghrIcKRo69I/8eVwGZmul76fofTEfby/py
1AEjLjO3NLI2baXcm1tO/1KQHe/MqKtCE7Rjoud1mDJ5WQkouhNpedIhZ8sqaweo
rbIlGkGisytVALFRvBb6x4ER1T4yBRNhWGYz4cxzytFkBeUaJ7ezadDBDVxwDq1t
0SlcpZrvVB5mznbbFg1xjI7xLJicySMoJejjJw36hYQYRzhokvcQoS0aRFGxOL+G
/mrMcB3eDC7fxiGGwZTFR+1INKYRe9qeXt/h9X2JgyKS5UaQY0T6qiU+ZP+kT8pr
1B8ulg780Y2iOmw2myoX7ofUijIXM73gQZj70cL0bbylpjdk6YwwQT/8ZU4a34q8
yAufDwlCmwkfANfFHuB6D3hMHBxC66Av00rGZdcGv/igfCvcj4y/acmjC0cJ8GH5
S7l9fcCNCt4pZ1X7DTu0vqtInM3VVa7k1LGsoFUsylizr8qbZe93dmnOGwVL15Fl
jrFGumrzpdJffpEAyDsVtaCj7+2JL8GLJGe49NJzKPdbD5Z3cX7qaBWrsKK1GWrL
DAVngIKOghSdKaZbLMZEj4mG2BBIxfHlfETpBILGJqwcQsTnUwppxvMfSz9+ha78
BjvQhMML/WOvSNTy9x2DFIi01e6XLr9o6GfFM55irYkIjm97E+bTcbIu5zbKJMIJ
lby+su5Br4SZIws+D/LZrcLvWRh59T4rv8gLbz/c08erNX87KOhs2fXh5YarblRq
cQeb+pZyCjjfPdmXYe+HmdkT3uK0dASEGUhnCQO+nlGjS7pOMfuKB08j4y6DGWNj
CAjSWXNLWniziSn4E5iMePwX0UB1BGtF66KD9L/SRcB2+JcXK+xo0eFNsn4HEjnW
BwhckrK1KDOvyhUpMy2zvybUOq9+QdR0aQvjvI28b7sQGLzsfZiaRhuY5TfA5U6h
Enl5DY3aQ3aMPVitOerH+A1dYlwzZL7I79ZzDtSJ5kZONxckyhNZ2c4sNeRelasp
eztNT6rncKsuYFr7z2IYgee8vyBh8IGWMmkLPeNdthuDyLrnR40f8IRF/ys2QttO
pcSxlKYU9lbZ+8rGPL/grpMuM7Q/N2p6r3qyiPUd5Xuz2YVqparYkoGSLYa/YZoh
QiL/IRDtP0fpKpiI2Ha/5FHG/jxDS6g8ozdjJJsPxqX7rVBdkHBNkx8S1mKQXzEU
2vm28MVTYL0G6pFLWpwU2sA8EbjtUss6lEDtLlO61FMI1sNpk2otvJDpEISDIUkb
/eJSniOrkQG6J7NDX7eLqpRDp6HPp9R6jfq0oC3jaiXgAg0hVAmf/Hlov5slPX+T
L1e48Xun1rzZvbHplZUGRv+9+j8gx7gVF9Qss5KNRcGXpR/ONY9+OAgndtcp/M7T
qtCelMOYw9IOsrBTDtHgWthGpFshsDmcDGHlk8WNKz2GA6sm6KYI8dZSR2rVmoQ6
QAhEO9dVyNBmMc+lj8Xsy5yDgNPmN5+1L7OQc/b2vvU8dafMQQiw17JDzJf6bOJx
5uRAZMDR3++eczz9uyIxFmfU4e4V7WqgHzzyfvjaeBjy9yX4iTdL/riz5CSJNO7s
yqiSe72POiXqr+PngwLtttOQ5YMnF/duyGZ3DFM+t1FNtWi05Hu4tJsQHrmTZrje
yyl4M+sBW9MjqSUDwgXlH30xZvXB4SUTOI1ro7mmFADsMU92xfg3Yfy+lU72kNcY
yYEZwsv3G/+QzUMJjyqZSd+MVA2niajkdNLqBWF6hr8tI71EoXnBrCJkDzTjwB6Y
DnzpnR9R3m4OXNHAyYfo2LobcmFlR51cY9lJNBhYbT+4f8U/CySHji92TDqd6brl
QXCV32uxap7AqO1Zc6o85oPY6Gl66JMxlKdEl1ShW98LtYWqjEKlI3ENRIqSTw1o
6baenE6Phx8u04tbUFLMk5NdCRCJ3c/f3paQXBHuwnlhhLl8XajOfophvBlmWrhQ
mnZziCvD0DHnt7+vQ8YG2HnOmTArvSSS+SFqcGYkbkYXcYECDp+rsj5ePPZ/Kx/F
mH9+1p2RM4mlBGebK9B47JD0PdlooPGbbzMNvxh3GoNWWayPTnXNkluoRm7lHsEA
DvRBI7JO9KLTcMabkphIYDz9GXYgVn3TFvTPH0NHvlIREa1cEuugLeuUJ1Eo+6Vl
1372UFrz5gh/K7Ua7ePT9dsZYBAAy8PiD+MZCeW7VAYmpmEGh/3a9DidgqNBr0Q9
H7MvxQj9SCY3ZZHuX4phU9k+NQvVExM/pbz9JOuCg3YpqcbyhSbKHoyCwm75i0hp
6ajPvAjGiW95ZgauMV8hOn0Z6MImrmicfLBsAb9KVasi8uDV7tndHXqoiKNdJPxx
+tfGOb90gscrsCOpIJMLauwdtQmJxpLd0IzsoXY49MeNfQNge96G2+tEDckjMfW/
leT0WQAt3mxjIp2SAw/RrNcfmUbyf0gby68dNMghZbOGyFydcjY27zAjTqHkw+Ze
nYcmJYHV5FtJ+5hYEMjNQzsk8k3AWuuQ0KfEdgvDf6ReeXZ9K/CM1ksgaP+iVNGk
ZZ9Y9Lz8J8mc6oCHZeQclQRS1l8uYMIGc7ogAtKonEtb2AxWU8JZm0ucStIWmamM
7WTRJ6wuVeMxrEs8ix4Uuc9pwNIe6cOP4jRUdftzpmPKgdyl5sa8BkjsnTGCYnkN
gAMkoExVpmYWIeYby8GXCEXpRV/125efrrZkbWE/UTOLrm/GPhyJnqMZlUYUaECE
8VbEwdyigQgnjPT3P4Y3QKGY5zikng6M3KvtkX9DdXFGB+hYfjaJk0PnQ136EKFx
wnbuLXwroIMC78NlZtXfUVdIzhtuyzg2sMcBDRNgfOKZSA93UpqaeXQd/wAaQI5A
8m1EfSdgKZWWrJbU65QUzGidmWUuwBJqW+WlBVbDfYxDoVJPxZm+3V+uVXKLFShn
QWYHvu8zOZiEYbTdSGYsHrWIfM2XuychQsa8nJueRY+CKMxJzCYUYu1imzmgw1/v
aClbCk+eAXa2ouPuMYk6ydqZ5EPpFu2RacAXUz/nQlMHS2keN8an/BlRDUQ136qd
w88R+a+1cEhEGDG4eELh7wwhdKRwi0hwY3bVMy9Vs77Io5lI3us/pHpHiHj67kAN
yovffY6zE1eZ3e2FJDJeQfW2rEDr369Nz6ONDFby3c+mBGviSHlrfdWsYbiZ8Blw
bP9m6Yrx4vTZ8gihgPfwOBNXbFAgHKQbYdDul2lnxuN7uE4qtYfuM5zr+Dtc3UG9
XEfUAdhHOt/rlsmM8UWddBHqp9hOILcdqkUsXmbIR6+7DMzW8ZAByxBvR9pk1CUm
iukbW4APzkeAa9TV9XsGhtDR9811hO5qK4DEhQB/grZvpdYZKDNlHDDhndtHoHRV
RfT/r/gEPjcD9NN8c5hnrPZ61698L5GQVQvhAc/lSP9WNW21IYbbdWZj5R017ZJj
3kI0vZJVltjQ7GvFZ1OSEuNnej8C2QbFZ/LGJpeI7WCBYt22ycCFfxtLCT6gUZKi
l6KlLyR7sAcQCYGmwM6RPRruchAWhwAHT2+YR7cGgpPOH9P/u1+kz+gYUVRIC5+w
J/YmggyUQQOz73evS6jYhZzO+jdBetKjS8NNpGoJck11UWAjCa7NxiZQcmoV7GaA
0FI07Ie6+lg59n63wliGK67oMSMbtM7cJH85NOpFzgLNQskEgoxxW3NEyQtaBE6O
6njOIIAi86SYstk4GkCNrKKT42/Aznis3wz1NA3YGMFkdtaVc+7HL8tDS7yQfTWl
uQfqxq8NeL8J/FQ0zsaWH2WEil7PW4ypQmvHcEYJGLxWeCGlIqD/KWAd9Wa7CCtb
yi0JafhJ97lUqG02qpHC1/dTOIJtTolv5tdin2vrypriHXd3hKrsL2T4uAhOf0Ib
gMR5KC8HeV/kqolgNzy1D3IgTuvm9Nw8thoL7PLhkA/EXn5jbVGIQHxBKKkLZj0H
yWwZp98TusktHvOvdAxvGaTqUAMCJopLQTy//FXzaHoe2w4z1NV9bnmRHoChkWDX
a1r+zlMskBqw7+U455Ci2+aX8bKhP/0HeD/vkbvC5J4/OKA5d6oqCZ0i2RcMVCwK
gGR3telFrfF9HiI7j8u1gQM8fhsGa08KN5tMXdWcor+Bi6adklR4LmJp5scZ0lbH
nZLVF6wSkXt3fbx8ENekRaa4NbUbqUsuf3cUPR/NWaXrMS8pysGPL+BM5TRS/ThJ
26017n6kbda6sYfWNkhtxz3PcT3sN1avGnVtQs8mqolmShBNwwRB29sMLhHzg9Wc
1pvDCTFGD06j/N4m356I/M0DRFYq6hyhmLE5Bmf5aJUewjeS0ZUMo/oyqASXjHeQ
K9nyHjqjyUu0eJ9SNezU+aHl3ICnQbQTsXHGCW5z+b216kWx45Ebi4W05riq+hJC
DXg2h6/odxa2fshL16wH7kj63wqGTvbZtG1OlqFPxWIPUATcfiT02MKP0jP8Hz2M
JEGJiB7ILyEbySnRs0AUxS+L4/ssjBN84kqXdr0+Ry6s5XrdoZuAmCvj3mQG60sh
UA2/JUtlcePC6r1HJTxE73V4UsOUFnxn6B7jXWAxB7j5y1Dt0Ssdp+RN/9+nmupp
aQb33RmxV5BjypAwqgZoI4anoi8rYlZlDE6ZCFUzoHp/RB2NrQ9dEjB04g420HHL
R+VzEp0xjcirx0u/BQ/rCvGT+b0AIGyj1wbyHrlMIxwJmkdDL3AHk3OgSFJl/iD0
YIDtqhrKQU8xEq+wCeFim8kdQJbQ3HFxUR1GQNv+iIZRh87hd6JmNewx15qjiqlX
AFiKzXjuvBUMBVifhnCJVquximmwpV00N3AaS95cclBO5KruQSN7KdETan7ow2Ht
50GTyxUygjNDaoEq3uT2jIIYkgMRMj12gxOjjJauHw7RaKZlD/kB22S0ZAz49Cs0
klragLIotAA+rgEELm+0LGt1k8CcNAMIUIgtkBbovrFE8Yr+SavreWNkclbERdA5
IKGEWIertFEDfiqTTZpJyVdiGH2phoaz7Oj6AiE/oKkB8LZqh1Iuw3+F+HRCGlOg
/BS7FXOwGvv9+KucJacgw4FTXesQu7fd8vMB62ieO9qkVdBzr8TpBnS4Zl5OtXeA
q+MG0VFrFUK0Y/LCuIbEjKDKibenz4ELuELZG/REAEUyMETeQKhpp9tXnt+hnTSG
d/YA7KG1are1rpv+JHSfZ6hcmIRKOOI0UYkAoR1GO5ca1onyNQ/ybzBsVXjPjHBW
E+VtGIhh77SYEUs8iVGBygSezX7prWpX6IU8XUDRfX0pP3EfRqbPBCxNWZntBsgA
bPULlEsO/+lKDfGB8UpOQhqCFsL/zg9DnAGpMGpZlLxbnm0CwlHJnLKDZXvE9fEQ
Ysccgg67hMZkgKedG+iQW9YTOHHT8VaDaUc1C2bpea51zEe9Wlys3PsUy+NFC2RC
m8wxvr/3/Fh6mqYAlsi6wPWeWxgaYWwm9xgSGjlgFa/G4dcIkenpUq+zVgjT0uj7
foJxslTy+EsLZ2CNn98mLDpReAITEvreLgB6YFoQOamfexLrveI7jIdrMWt9nyml
Q5BnCxQT95PvtOyVhMxxjYadpVXbLNwpG3dpBXU5kMkWvr2BykxBqQ5JkO/3eoa3
36UnIaUPVnOYU0OfnPvtK+Slci3uJ14Om955sID4Vklz3Cj7aoQfxfyeuw37yvC2
cBROp9WQrOXXrbeHFJVICJEWyKqnLgMxRcV/3FZhFIpklqsMEKT+KCXArQcLT80x
S45MZl4+8ggSCC4+11iY3p9yvHj+X9809ZTPGjD1ksnHOxljk2XkdYR/J6LSvYHu
y1UE40d15DDGbvOGWY1T3Psm+/CshE2P1MVI1H5RUHUGCQXvdCUJHVnmEVCZQrwC
drCN4C12tutj4nxPexQp2tDuWJcRrffM8AXGhhkaYU0TqaiUsaLafx9t7C1+KF8+
ZlT1Hqb8jq8hGWa2M6T5R02BGnrE/rpdCLPysuc95njyxOkHg06RmLcQMNhC1GJe
DFutQTwCpkJM/wMc2T103ykDDU7ES2I54+igYKjpaDwZgHuqTUp4CeHuM0POCxul
1Ebbe4/ucheZKRYQIP2hacUrNh2YMWrmNI+Gg3+0EqOEKmwSHRxu6JKVp6Gz8KCD
qYHltAHvwEW6443Wg7qhNHjB+EcPaT+hyAKUIaZ0Hvwi4HZg7q2Jzm/reCIm8BQX
LVlNgP+tumzo0kpA1fXt9/xImXzcOhNX6JNyb3WwFUhZHXYu6rPzpekjkfTStCHn
3sYA3UsfZRU6jZJYm4zjhvN9ECOPSfdo47nKltTdHspv0T54B1c5bXrY7LVp2FDv
uowRQe+X6ePl6Tohw9mSb1SkMD2pkVOfIyBUvV65GUtufRQl/kbqnBzkhzy+HQPc
RCOLBFc7kZJXCCa+fUITxa855jAcYLo0amDyHbAO0Gg4prtxOnsrhnK6bPezFBWU
UQPjAifoYPOPzCHbQ1U1epuo+5/TB04T/+EeKMbfq8L5BwDqjqVic3swGxjdc5op
612c3f1Z3uokINRFkBrprl+ad+x2/TJNfwCK7V2KwcKdO0rnXyLqvABuydTteUnP
r2m7k6Aennnsum4ClL+VzVpNyTY1/L9q828CYOPqHjEy6U2rsiWK+SlWefnsRlms
yGmPHNn7uuJrqF+tinAzYnJcXJhaZf01LV2zmZauil3mTWhHwGTWDdonGzD/4c/Q
k3ihQfow9UMYW1A0Mg3rS3hK1nF2s9c8LLzo3jR44Xw6Nbzivqbtog9R0yKM1rMz
4nkha3WOOpvWQYlpRkl0mdaspBpDr0WL+9fivDx8u9oACe3IiRqQLuX+Obz63Xp6
Cll33ItTk5Sy5+gYLIXnptNJs5zuLJdfUe5PxUCg7qF3CFA6dHpVIDovMHgQivaw
Mgu8lCjnRF0b8w/7XH834kvvd16ZH729QBmfLYqkWDKVnCojPl1b1C6JqRKvq8Eo
wk46RrEtNYHbEDS3tH5/z3Yc8+UzyH5fDUoA0sp4SCajY7YhyloL2Vm+d25YiLqi
uJ/47d+dTDd9sdn5aVYzXeEUeTpFsxhB8/O9fCJtGs77CCfYHOcfM9befblewXxM
c1VR+9oDhGl3rjWHOn3kSgR6V5UT5vKHBTMGKljIKrVKzVLkKbwOEN0C6Uujyp6M
tT4ySnGn7V02sRHQSDqPY6VfRGTY+ur/LKyF1rYq4gr0yZpTea89zjOxbnho+NWn
RwpVwVPNLV4/oA+hNSCgOWTF2vLLSsMTDtv2io4J1v8EfjHV8DjNHPxrIbVTnVo4
AsrcR+o3e383o9IEJOYUai7dtA6OCzHMjVXn/bWdijh8cXyOhvQca33larMGeazP
EkUeLuiIlh/+SL7KmQJKWqFlS7SnNcQYhJjgfHE983My7MvhOYFQbG9GLNaMtOOt
wGVq2z2LUmcJPBCqcbUKn8UNWYQMspI/+zrc59FsQMkjdTy6EvU0ICSUWR6AszJM
0TEe2q1is5PSYCTGVPzWcs8spRajl4fISXw5mZ62IKkdA6qBpgZMY7616R70qmwc
ohr2szmDxgy5BuwdyJ1EaEDmG9wOiKfzvQyEUl4tlauuBfN6wVWxg/pLjxgjsPIe
FZXZ7jGwic2swN+wsxlIY6tom8q/cZHyyJjnX2SxsyWG5rZjSYOpfrVdEbE9gBqw
HNexQY5OXnfupVMgqDvCdANiLD2UD7SnSodtS9miDT5AW6TgWGlblcujmCwKiCtp
9xpZgylP8pvNk3bWj/35QVxbt6M8a16GEAEyXuIDDy/pPq8MJBp7uIemV0fKiU/L
GOnJXQxPSlIpW92lqCCXlT6FGzQfi1AHS4ye5ojO80IH9F+Zl3JWtDvKwSa440G9
tlhzxFjLH1DPo/nIRKX4CZnFf9qkvi9Huo7/L/k8+HIgJk7e/cIbwd3YIkGibAp0
EmKox1NJtqWzN2Yh7toFZYlNoRes7Z++DcssRBL4y7pHSZdsJRf3q3u3PEwGjdhK
N5fW9RyeT7aGUi4Wblt4XU17+6B1pD/IWTjXcjvTIhlgW4uGWK26YJFTzL4VgovK
UXclHFrptCkC8TlrXdswGfu1qMA1HQqnO+1xN28wxlkS8lDakHu5bgXOAjNlOHna
WgVcyksqmWqwbBexbTORcEt9hS4qfXbHOA9MFsVUeDXVC6xCMeVncxHkoJ45sgYW
6+Ib+xRQmjza+8zX/sVOT6Gr+ekG2wu1Dt8/4W6bCs863lwbmRjiHjpy6yqTLPob
BXYF5WVHyhzlLj+VF7venSh15b7SHxo/NEesqJ4sHaQvmvQ6RXeVD6U1YjpgI/lv
AV+gMlsItvsmOzeBcwL/MsVG73tYgeMVwnLJBSw2JsIPKZKlM+hATzXkXLcIkimk
mElIBXLY0N2D55drEKTWy6W2D0h9c5KODtbR8+MKUVgNIAQcNuxRxZsI0DXc3grX
BlXlZi8arKraNOx+v7NMClZiS2t5unoYaKCT9UHN+Ci+jTGHzoKX3T6p61K49IFz
3zqDJocSFBNGz/QFlJC0gUpv9/9WvE6L1oLM6o+RYPur0rjlt2eZseg0cGujqgBN
Bj60DOk2kGykE5hniS6sTmay6m47nbMo3yXIe+N2Rw1MZLUmWHmyxU6XZ3FB5qvA
LWFiqRK/kjtl6UkdbkRtHbMycGhInbV3Q0l4Dfpo5J1VP/0ACRALhWCicnepuLzz
EBKp2kOVEb4BmAJutVabv4aZ8X8Q/RsIINWgV2Ex0BRzJf83t2L3VmQ2D81f19sS
0fugWfIWfMiNwHyo/HoLdZhxvsLmcLEhEbwC1DLgNTIymLS/cJ7YrSmPs+pIJc8K
4ilvEk24bgCSwy2zxNX/J0EIqP3gajmz5yMERjRwz/T4VwzppVJbUnn6bgnl0g5a
ZilBfqRMMbGF+9vfPvOLIJbrBcyiUO2jNKkrONwx/Y5omqQ4nKvOppk+8OSxRiBC
0frvWNgPdO4q/6fnK94Ahf8MquoAhILZ/ZTQ+1BJR7YdFvB23yQSfxBqiNPYEbMM
q/HBQqN3EXqM805lGriviy9a/1CS8T2GYphBuCSG+Icmk0KjUWPD2Rb9Kn+0kR/W
jXQon7f7a7JI8M7NuqrhNhcN+zU4cMcgzYrwHJB/zCi2RV4MD1Olf3Rk+Pf4h1wl
3meXi/7k3xmZHF91P2FvQ3wK3ph9hnX5iQt5OK82o3P3vu2uOa9MMUlhQ09rtYBz
Hdgr4tGsxnHcW/8AH61vQtT5UZgsYHCNpJIfZ+N2qg9xrBobHCQ+pBNtNM32ase/
9tFx/t3tKuOIR9mzpnSEXdmkPk4KsM3Uhh3dCM0X8+CV1BGew5iwGPE/qabgKUgc
jdQx0iDF7XkapGZvpiFJ3O1AsbTO4bKrJUncHSuHaCbY5oig8b0u9pcsYTnQKDa6
6y6JXHijpcxdG4MDl2Tkiz2mWZueJMuaTFgqAmfBpTHDVvjK0YSksbXNLvNcfDI+
p1X5YCzIXRyer8s4Pn4YtKOe/YvIHA3x+g40ETVHrkNC2VjGtQ2rytTuD6B4kFY8
JJTERmKDo9iSqD0QIfiGa9Xr7fl6K+CtkOdZddaxtnbn5ZCOmB3D8WiDrM+IUT7p
iBLieCrR2wLeYFzlhfsih8b0bD/6HzL62OMd3ECrwwkcj69AO+PP7ciXjIDWlnOj
vkkTeo+wdddFXKtOtoycDLDj2XO1eF1hFjthXKjKSRktAzPRAaPbQJcaGeaNrgle
iXgcnofw/R/g/1xN7ZQtIvNreekm1zAISgJdkQLyoppd2ilCy5MX13QChDo6EVFF
UKks/+GLEoFtovvdPhw9IkfOpgcJpCEPVTV1aXoKsVn4zp7IBfmL4U7Qu5oJ1KD+
Bp50Tgt/QqqBzRUE63/TLStor4Mp/O3/YduhQKXw3cMLKjMzZyNccJp+IRBH0ClH
CwOkHQTleHvK1UaUb5Sh4OQdKM1cjxYFFhgcj+vr4KLZUz++xdpycO1XU0XG3HSl
5wPbs7AnLCjMl2L6E6WoLlkA0onLyHjXrinuXBW9M3rzEmifZnKBAd5v6TAfAq2M
wyoeeTJaeA0vgey+uNKgoSh7d5bp9HjQx7BpLfklhPH8kPTjThWBNU0bxSCUxHib
61PeYCg/XffYnVmY61OtsjDf06fi+AAoQo1gw9dlyGv7o6zd/tww5kSgScGWwp6H
r0zCf998vJxUQmcreCR4f144yqL18nE6NCKVdSsrNwQtJMKxmpuKlHzcnOlJj46e
e+5SYhC5Dz3d6MU20WIU9QnR1MBCze3qS6egTkUZpsggpoQUusyPTxSNn0HMG3LQ
3QYTo/fTKrtviy4hpfto6iMgCxsrmb2a1I/pPguhK4svsmTDiZ4bjfTwTs9jAwF9
KnEAzAGnIbB6T1Ol6cRJjWfYVU7qhJgnkh2zvqZv61ZsSKltr7rbpV7IxK32fbs/
xp+lkje+5KmJjOkx/8bixwS6jDtPW1JiN9kFCl4Gs+yanXiAopi6hIMmPaISymz4
7uW/4GmCcV0AvHmfefhatFXrattJkOej/uia7dUpImnjiwn2Ir4/ANlZNVHSIHYr
gxSx9vIk3tim6fYyH4xB9Byf3a3kkYSfpYwotLzYh5nHWhURl38SibhV0E1O9Gpi
zYe4Lc0H+zP8+Tdhm0OPfxluSmyom3SDRdu+lp+A4VFpbsyD/0YNV4gSwuRIGC2j
aKAvRSJb7HzRn2LmfmUWXBOrZ091Jcb1qhkxrTmqj1EARGL/TQ4ZaEJQbEVBe3z7
6cFqLEWU61FuM/BQQiN+TloH1/dBU0l98QAGC1PjE5K+//sYXSD2xAthAItBw+F0
cbpyC6Wo7V2Ga1DLXxiOj/MQtSAhsVCN7PmI11Nvsio5Hq4bIO1OaHDJMoaGJdB3
g01GDhr9MApU5tGT7xb66fEGY+L9dsx1XF+4yWElJyKm8y6RF6Ie3e+FHSY/wiob
JPJbqFVhwF8T8p1aD9qokPL7zSr8G86I5Gywdwj1crb32R5BvZbeI689Z8Uz+cQ7
fzsh8Fhll69dodlIucYcgRPyLnw8FJudflNnbR853LoibD3+CZYBvRjhrkauJb/j
SQj4HVTZIuLK/r0XE17X4CX7wDtGP71GK3VS9tz8FdBrVCfmgNmDfMZFIoSIoBYD
Era8I3YZJuKCcefWiCKlLdsDtbGlIWUTrz/22ZJ+l7Luh2EjjI/qNEPi9xyAEBgq
+mr0slfrjDILcIIfYNlIQlT3Y4f2gCF/8+7ul64AmPfY/4g1k5u62xxHvgIG2iOg
az/gb1epy+JiWNSNQ1Z5/kVfSdKAe7GwK7FmMUUVfVtp3HU0lBxn7liBR/PYqKtC
JfXeXcy7HJZcskZOjVfiWYKrKRZM2adbywMmHvCbii66ZLrcRYSsXDxg4Y6rKnpm
ckGn7x5wqtyFhl78TrVvkNO2vdPfHPw0m1PuCLzmpusmpR4nSUk8P8Vc191D+OQO
LmKSUSLrddUVkszm/dQlgn4PL2iHmPnRpvZAwl07PT7oRUhpUYRtE0ejSrJ7SxOb
++/kl3zKSWXbSkaT6H8PPWCF4U/EM/WWOdXeyqhuAvZf72Gmy/MiU3/obNlk0Nwl
FSex0ZVslYUHpBJDKTtNrdVscpqwKrNpZHh4ZxiCu/hMpkHm7SwAqbUSIXXmcaq/
h7W2wzr42VogjURxAOdeJoyLRx+urJFUcHXMNT25zTVSv+cYXcz8vubDMQZlSoAS
avMIByBkN+uyw8LQVRrQTk/wLVbw1FqbWUP4voRLRZaN8y2pxYIy5Ojh0QEVuW00
+vnr8Z/1iN2SNrkNi/WgfP44qL1amzmjYSqI9W0aImtlHxa4KpewatgMY4M9ZhL3
kS6fod0jfT2aEDq4Q25fIcRCFQuC+8MjG1fg84zjKHOH0OC8NDbB31jrnPIodHSL
6k+3ATVmwyFSM1gFIyRMvVikGUJLrl/zckwhZ9d9F/ZZHW3lLB8CcucuLL/o2WLg
HlZAXXs2h03udTcQWILYAhbUcKmpM0dPs0m2HFwsSaQVP/1WL4Fb5HPvydgVyEfG
81bnq7dXtNqG5wz5OGBi+Gv0/9ikjXwNKxJfCV42pjp446smUn9jMw8dvLpqqzHn
5bAkuAieiVmvN+JWSI6CFNNTlzEmL1+THuwkNt3d0ESy3v8qrU1f+YCB0K9QIxss
wJMvlQ8IJjB+Hj9yAr0FcdALcURbFCyvA+wEqcPTcqPzuULOsaayOO6cKHorXvKL
k/XA/utCCsHzPCOwTKcDagWPylzU88qxfacwRdLMM91BJtWHITfYmIquCqnd6Yqy
ktmvM5d0dXMaFe2XfL0AL3oTiX0/r+XdOJHkDw5Q9SXewECWqfsHcXDr9WvQqZPr
KZyvnPmJxF0OsIUiw63y5QNJsLjOip/cftCNGeB374vh/zCFpAcCcooAG2EcXQ6Z
I2RkJTO2FA6f9eLbz1OHNDTSWFcIOo7b8P/wZg+HLwiHL3xnQbSU8b3E08IB+48o
fkc3Vtyjr0vCqa3IO8o6a6bXKUa0+ZHU7nxtaR59xoQkwjoj07+uXT1psXr6+H/I
byaROtj8ooLn3v+szfjA8dP8QGp40wlaqbXrZVR2DGpOmiREuECc24vKDoMqoo31
aVmgQQBK2W55eKXcXPnDfvXOfUxkXSwO9GG/2dWDUYFLWEnig2dx8bSRrz8OVYTz
jR6lVtGNPORnUdzkgPnfW0tcZ1JWCLsQvs589wMncgITJoanWiBeCjJ1/4zdxTpc
c9HGHOJZQ1HQ2Hjb9hUBEolhYmch4LtkzFHqo1LWjO/ZCm8SNWYXF191afz/BeGi
My+UL9siCFvPKv5Zl/s3ujkP3cxzsWCDLRnyM7Ypy7vOhFenUePk75V2Ji0x14fv
sL9ouWH1hvDHHAPPFGiVMRRcnjnmAp9DIN0qw9lTkV26uNbB1WhXg5VI36L7DGrt
BTVMwdTgBEpaGeRTpbbgmAA6TdDcZzyroc5EkZFiEJZdkI/+GUj0ADR3mW0hSCBJ
bSdhzy+XNiGSw7jTo3MgGSX+IYMVGz8wSiSx3Ly6PGzNYvhQFRW4HhXP2dlAC8pz
rnOsqNmaNUxiNVH5Cqun/6yhQDXZl9JPz8TtDEIvZM49D+QpSO1xuOAroRMpMKrp
uFUWE5vhD1t9eIyHfIhGMBaJUscUJF9nggRSfp1ZBmSSIMoNEjt/l2blRK70kHdg
ys/eE/8fgPQxzpPaTqmwVUKDceTRpD9lpr4zx/dB/nubDjLMR2a0Qh2VKXJrxuK0
W8a29ZhNfNC6rCXUDd9TFiHvA8DWMMVF1fZ7Pyc42nEJH+nf+sXPnLA9U4dedylv
MeTkExfNXvVD4iXcGuOcbVsknlcaMWHpAqBTks2RjfI19BLIiuQMK3/9sZKyPo4A
7sYcU3Wn22YseH8Z/7Opt5xhAMJOoXSw9P/LMnscJ7erpWXNeIH9meDrEDQiFxru
Y/56k6j2bpT9MqXqfLz0aKAjTkJ+DigHoj0Hh6wtaMmX9mxYWkln2yspCcy9GSEN
jMo2+xpehHDKGbiAlybNvqBCewOal+SR5xHga8DCZD/TKkSB3tdLUvwkYcfCfNqm
Ylpr8O1Ufmf0ZD3ps15VGfR0rffF+XxokDqg8VcQzYUk+/omFfAA4pV0wpf7oKp8
j88hekYH9RFW5fxRKtICf9LX0EaRPX70BqBdW6GW0dpLcnyIL91+NU9WsgqMHSUV
HPFCQvPyr6ZUUQSJwdnahBOxB9nIb1+6okJweGoeDnnRDGr5+xvD60GnEyOe9rlI
cS6m7++2u6G9iLA5OFNAp6E6k6+OPwPA+BRz0/VLkiWtO4g1OOI2cmvWHUpdJc6v
pWxwcIRL0pmKGovUa42ElSQocHSMm0TF2EnhBBmbvcSYG6axjS3I6d2/7bvbwzt2
7m11EFR0DK2Ex6I3AJUAzK9V8tBzBAyQjYtW3RWDoLN6ZDCSZ5r47PdIWdUyIx/g
IYx77mIkt6LP9Bw8OdSZJ0hoNWd3j290ZlAyNQMRYt5Eo1OaxEj5m21+HeqSPj7l
E8A0pYtka3bLgnJjM3wF5oYVS4mTuIuXIEgfVETMNbQQDxmmFUsMj2NaA5AkIbAi
c6CcHBqq/WiyLtrPWUQEHg6W8uySGWuLo1s81jGC1CuaiLcyOjKbLgF2Z9zSEj7N
4g7WO86jA1RqWLlwNtfPiCDNe8J+JHCADOEd86prTV8rEzvEwee7SFgG/etyf41y
jD8ZORAf1Hnx6Kajr41p5Psl9zH13GjwSy+J5HmLHnyMmdkOawry7r0wrZi8J/kK
tXDNxW1hBDqB/qDQCP15eiaEd5BmfyDl1xJPLVkCqaSDJGIolN+C+L8g+kUcfRho
3tw2aMdYJp68VRG80GmIfFB0QX8IhxupEW2mrOQtiSZZA8eH0G+73BR18Y5870it
2ASr08wMS+sMxZd/zdlzV2LefrftxhVTUKTS+AQnkGzoDa6XT14AGFzKa+28qugg
QV5UNxPh3QwDVX5WLk3NCMUwErI+KM+lo4yglOOi2xObJtqcdHA0eKMZHJo1wu3X
SCcnfoFbVKUa+eHNP+lkA1IMIkaKKOs9CydPu4PeraG1mS+AgiONw3T4fMm/6GW+
icQvaqSXkaqdRotjlW+jDbE+ct/kJ7ZvChQIKECLoRZrafVTNU5bTL7EuSUCOAgy
nTbQPIt4I/fcXeJ189ql3aAI9JcwX2WFomjk9TnY9yhzHpN4fy/11PXbHZBGQ8Tc
rEG/K/ySeFpnQPLqphPUhFFUMMgtOZr7g3nnWPQ/4+PeHVgu5+prfCY+731a/Cub
8ycnbyYYnHUO6rYd6NheZ3WELpMIuTERQ1H34eV9n4dkOzCueUwhL7qe2Icb3B/M
Jo4Hl6QxHHCDZuTfoLyE/Lbg2tnGrzwrJ1syhsSxrG8eCRwcA+JgpBhsS6tYN2Fo
G4tXNaQR12GFNjDYaYhgEpqENy1PzFyboC19/JT0UnDn+0oyQEB0P1htXTzBZkho
GpOQ5/5pcjMZBPqXm1qOebJNWkMCpy5tQnPl5oyXkCow+2IZg4lrw8kVcgTC8QWg
ZzO77jXo02QoU7k62Z7OTsid6oPb7vly2PsfoXCqArFNd2gTG2sNDTvAWFsRWNgJ
PQ2ubj4Z8yuw2Udjx7/T6+AuwxmM1sMI3y6ig8LGC+5NVzkRkbmW7B7PRKOLHkeL
I4LdoiKJVqUY0EXwTtddff6+TvO7lSqZJI+EXGdL0RoGdGF7O1QCN+/s0VSklAaa
StWXfj2dvhqRCIjjZFMrv6tkWrjIgIdJtyrDlfW8/WcrAAwv315XHDq93Oq9fQtv
QWJBZ+3KpSaKuu/buFwfrIBiwBcT+9SGmO7VOrXqq5PKF92jHPlygtb2QzB/uOyC
7zqspMklVW3rF4pICeQgm5Vn1DIBVltCF4vrQQ5lAIf1oD2YxPzZ4eCneL/gfDKt
TyX7pm8V6SuchRU5f39aObYXvQGlFLIHRzNWsrLx6wgh4usGOZ5apvk89vbwzMdX
GhBO0YBrihGy/+Fdo6r82jWwLU5mMk0n4ttukXt9SfIv7pBaZROecX90do/61LI9
All7oTMT2sagZekpNazTjROdZVEf+jFA/sgUUUD2KnzGv3ixDpP66cRfMGLAutwx
wjsxDu+156o+o8v8z3cC3gEiL8nxltcbMNw79SWZ9XTK2hTUBRFejOA0fEJ4vBhW
AZF3wbKPFcXCpIzRGNaPH4Sj+6oIILnqF5aWhlBE6G48xSqceSZtGnhT8naUR6iR
G20n1vuRmg3pGxZg0qn1lc2S9HfC7i0aVdyM9WUZgh5xpUkUyeq/f1Ih867HDZG9
zo1QcX10H3TeFmvebBsc1iWM3NoiUoWLSkgv/VR5C65RSg3/z+C+O6LIt72Bhay7
Mt2fFdGUH+T47zTQx9znQ14mbT97wepiPDu8Taq0NbmOcUtAEgChzZdFpzpehKtm
XlyazSMQr4Y1ydc1cGr2MAsOKVfb4yTIDA7yJnxlSuS8rmzgIqmRUr7a2YAUNWSc
VYR+aM1w89cU9BLZptk3rbRe8Pg39Rky74TiJ9JrcUt5yrE6rW02LdX0RrJQcyGs
IXKHSAC1iWRYHlEVFvgj9pd4ceIV+qIkoeV+l0+/4aF3vgQiRUUNDahPguPEjhg2
HAe59YkiVT+c3tq+5+tVhIkmVRKIiTqS8F48IqI5GaTCnvCnfwnUhDHkALkchKmQ
T4tLq7vJGR3dI0klKGNX+JVnIHfX76SwalowE4SRzww3Q2uGSjZhfa+Oofc4zAuS
ngRViVIUf9HgUw14Z6KO5JlhsxyBVeUZsBGP1z70z3sxILoFpsaeEKpKSQpuy6k8
NcQANO6xagLGtET4VWWdO0Hvp+hMnGfHCDB8xJi7bZOhYlnxmybyIE0y/uODwSGC
o8STifr6vgA2ctlDnKLoJq9dhBGZMM/lZDgRcckFn+wnL87Smgp+7GF2eZdB+gfA
+X6C2bOZfvKyi8nKyx4DoV8a8yUAdhwAHh5/Yy3d+bpHnLanhKucIzfpjCXdGaga
S3SkOuQBI3gVxqOYRxmgvKPC1yCLW355CzB5YliP5oheHyI8O3otKaqRj+amn7ZT
zEwSVbbfLKOq6zMkZo2aI6pdDBNwf5zjxnAd5gqtcaUvWOXe1rQMC0GMeHgXrSgW
LBFbYXlmOuprscHo2GFQTw1AMxUUvac8e5sA763pMPweabk6CYG6M3TdP3kqAOio
NKPdbEO78a7dQKb1Vuaxsswx6S3B+LuTQTYRY4MLfQ2y8UkZ1ZoPdHtkVGMLyWAp
319kTuqOeF2fcNYrdyf45xG6JT9uymtuywf2EQkni+zzZUGGX7y7Hrq2WzJQuJz6
EsAlMiXmeCh1OId7ZYtBLxZHrmiIZVgxSUNkz24DGQsPNJ6va8AennjA2UrwiNWM
L8fx/FhAkMZQUeyblXIeFZfnFLdKv1i/VQ+xeBvB4guonWbP2KuL7oFlJ12FTsXY
3k9MJzY3eB/PglL+wD2JkQWumKMotPJiHYst1lMsAyNnT27djQDAYy781MiPHw1j
Yyookk67M6PUCwi1liTcxySHqL7iZ5FN64V7kr2TyhR+fP+oY74xQ9tTS4w+nji4
zkDdXUvtDR529MTtPP7JJgZm0W+HtZSSbdqEOC+LVwz1Fz2ek1CC5otL2O/TysFr
l4PKMDYwHMO4mq+GTy1pCsJpoUqLoU8evXVIhDREDdXnn6ft5WSpT5E0fydfXQ+n
elAnPoh7TNusfx4rAjKwFuQsyvYQL9Dc3pEA7bkNB/bVfnTYHkjVuoc7lzoXvZ2w
XqwXKIMVO16irFWQ1BW5IdAODepfjCXkInuwrnKsA3H3e1Zc7ubCK/vM5iA0IfmI
Ac3s1fbETEq9RHyZeslCsl1z1las/PuUlaxxQOFi0wUusBXjHCnFxhgfU77FZpV0
cKAu3/CgtgRoyapRxtnTZqjvuaWb7uWVs7Ppqhjc/gE08sJkRGJ5Q45XzfM3RXLr
dWKeAzDk8Bi+Hv8y188fw7B/HcUz/l/r/7oNjE5O2uEJUeAZ57r6w9bsBE9keBm+
vLQ+wPEZJ4JIB4SSqHg6fIjSsgasrjHmebRgjYTwn0lYYrqVFZxVAh86zKjjpn1L
y6SQ8UHozOV6I0MAgJs44S6ubv200FTF6YqWRWt1gOxeFfbSvHLyYX3an6GXP4Nj
sJ3igQPMiTZ4FFyxxtqPviYTmz/ur8D3TTI46mTkq6QeH3c4fHXzuY7s8e94ONwr
UCUlGG/5OaU4/BY0PIx7ng+13WEiG/iEF65WVjSgln0RuAUeH8fmgWe2AaOhaNG8
qqkgm4Jv3RkB7gx34jRxxooizF0aUe9BlOdcdY5EZZvccJkI/r/TL0TdiUxGTSJE
Ti27QPPPnLhQJL6W9MRkJZAsgpLpXg0+TWcNfYrfoDPaqtZnCQM3eAUSYZI3ZTBz
VCsky0nkLeCHl10DFnCK5V9rY2LvhuNqUR04ZwFGmvsiRLIyIwHQdINSEFvbm9d3
Ecpa7aHLo+bm6vr7z4DnQtpvLAV0Dg166Anra2/M2UpO8ynuZi8mvJx5rWPByUmW
8EqNJ3Gt9JrUxf4Wpy/ZSxo8oTo6pCLOgixrQ7K0q+MXYx9I4Nz8qWkPqmHY6hCO
zsCnLYItCsBKLLsP6oepwdL/yiWxbTfxzgvoEBZP2AhujUObl/yQPOmFa8KVTHfW
hJv5vFMqHk18PRJDz0gQy8ik8mXGiJt9AUHGwzBSFEDUp/ZgTiULh8N79wRwaSY6
bSVlYEfRxmfOhyUDAZs+1HaA8KJXBxiUv9OkHiUu35cBzxqPutYTK2hJRHVJyQ3r
H+IckJB580Km6L/0cHa871/242WTz7qwA8/NY/xZio7vLbCR2zagCsXrPsDoMUeh
+WaWrXOczw7K5PN2j8VDrdxw2sjOjRxueHbBLi3iVWL74DlpRB8qBbTrXKL+aB28
EdTgTVJEmOf/rJPWYqrZQl+ns1bQhF92mi234uJXM/GAjJOwNQNyQPXzpVsvJpb1
gd5svbLdohA0twVORNDNd2O4SeDjwmc53QzarMb1rr2+wXXid5J+0AXgB6S21+Ui
6Fqt0X15a2u0jG437w0nqEj+l8EjwlNSq6aVNKR0siVQm6Xv1a0DgoNlSKUqDI3o
keDtdaaJCy7Xh2AaIRysgOatWu/W4FpCA2958pDzmU6Y+iet6EyZvROQbVhObakU
6U46lF4Sfh7krXJQUwJ9S3nca23neQUWIWjhH2bO7fgiAsGjCfVCq/8MY43YUGzO
6slmW9pW4ud4M9Awfqgl0WIwaV9qLYyGxm3O6ThCEpn8HctpGL/y76+sbpb6DJwd
uSEn94v/62fnuQ+53ba6V+Tbz6IdYnYLcyRuPemidtsY/5s7NbdeBHcdO4Rt15pC
+zrks4LXY/7EvDpMKqtHP7A5U8prCyDq1S6NHwW/HYUWxSjAm7IWsQ6MKgF3MuIR
dIm8Pqjq30sBqbCOxppNg0Rbvqtv1ysozStebyhhwGOCYsPZHPKkGaQckReElRFH
yANrVTqQeUSts9JF1pmklnVqFBXNyScFCQwAn+FzPWLyn0HF+8U6vtdI4RBmLAye
kyvzcx4PPGDAmEkLaJOy5rPMCRcc0sOmZvg1ikzWBGZ9+zESrErHMyyrubfReAad
G86xIdE369SJQCA6VtQXr9x0gae4qHR3jxneUmWmWfhmvsR0uYjwIKqEIHBIrICS
9ry+o2iJ0i9ZCIpwK3E6cTYXmeWf9fBhLox5PQv4rou5cgoOKdrk2k2NaWjtOtnF
Q8ifwYS5LZK8RSPX6WLKusoa5rgyvfnofx9X8bPaVxXtEqB8cqyKlik1X5Gdscbr
Z0ycHf/3CQNAi3qxuxKP8HbWBYNwiDYrQUSuCUcKpmebMZbnYhbZMB5F3jBtPlrS
5IuLutkcOhj6UI0MJtcKI8lgarXm1S8Fa5JUU7S5SDbuc9ueG+4DEfezKTs2ns6X
eJVnzic4MkOao+UPNi7b7906tXA+uyOxwD2t2NOiAAqtRinq3a5nSHUwzYfXfcS8
P/WhhhGslbwZlv2VWFnMeyz40iToKroWI6wVCQFFkYrzu/edV0vwjHqhTDKtpO9r
Oji07mhAuxmKt62RdfEB2jRoI0qT7wre3RfAPPrrOC8YcpFCgzDUH/izUXXJvbwU
camXZK6pQlcZYMmDWeEsl8BHiMONaTZHlcDQv324Vjg+wOL53Gq5Htc2calNhBvB
XySeqdnlRFR3nJRi9C3Wy3o4jzNPfFAOYx4yQrFQSd+wNgPTdFzpTBrgEgt+Hhk+
/S0M++Ds6xy/XWCXlQmqVtIbY5WQPZepCJSOdLw0JFCKlYa6F6HGHszyE+i9RfCH
FMMXWLBdJU3hYYKonyZorAzXwl55buIvNNi6wAhrsJhPSeDAFqr2Tw1YcSxkcnZM
5FzfWw06GPMqKHlbB2MWEblsNUob07SKd1+cKDrH43mRizDsuKLx1H0D6uMpG/dN
A08kLARIy3U1bZWGbRbZx/gWsHlzeav9LUBxzQXKb5D6Mk34bNCCw+r1bq1W0wtj
mW5xHJfz3FF3vF5JEOvTRXkUrxnttupGXv6KZ+Eh/lOdSXztM+O2TyrwSZikcsen
dvJd6MJ3PxoT9uqKDTmM5E8do0BQ1RVNIlOacOba+XfCMMlOa6Fwsohluid2593v
dyIB9bjY3bU3AfVMGraaRbBlkk4S3QhEtoiJZmJnJ7w0EaK6c23zYp6DgCbOVi7n
0iuXN6SIesby9uiyONdsOuX3jUYDSCXUc6kQnFQugIZdo8bgjLE+Tt+JEY3TRLky
vSX83sMHDPVH2xwb0lXqUoWpw6xolX1kKmmRFxM6V18JpFMTVn4oCwDBIuDEEaAA
CyVfBkK3CXgWreLxfIJzz1pbMUVPryg/B2DtWCOonB/YYRBmcjKXnng2UMpM28Ui
M1uPWzcI1WrspK4fem05q/HXjkU3myPR/eNtej0jiUYYCe+T6spAxrqEBc1KYevI
meMzuitgt/gnwMtXEcjg1/V5dgv+rBXOsEPgX7kJImZD3E+J9OiDI/7k0Kfgjf/r
pgwWBBLTLVAYx2Q7LHC1vXnY0mPjfo1SXH/xB+cfTeTcWPBlcDstdzw6mQ19QGM6
VkM1S+P9i54OZgAs7W70jFrDv2JbBGNVUe7IWCTfDvYuzkGiXbig7BP89oB9od+a
wzJzi/npuA4vMMoN9ztyNe2dp51i4TGgD6IVHTp9y6kRs32llKgnnjJPXOHVnezS
ee8hZjTHKWfiDvDo4zxBJDLweALyDyqp3zfDfEgvHo+gajxhQ6c9q2Q3kCC5s1fh
5UxPuG8Naca9aNLms3IBG+VgB2OYxKiVwzqQk+rAtFJTGhyid/u/wHu2DkI87TwE
gHRWR+gFghfwAdHnWSYRLNT+micVaVtYFRqIC2phK6szUSlvEhNWR5dyzhIh1ID0
oRGGpB9RX4ppAblltE7Iilk/0Whp7V6SPtCVKI3A0vzHd15gscXz3g4ntIJUi4C6
mealaMQXJxjmQ8F4GeSAA2tFhhyBue2g70NXkvUtVSTaP0pTIgLsiI4BcGuZCuSS
kVOI5tdXFFu+BHC41ONZQxZU94df3HTBsREKLa0lXQopsArN0eUbtSB52WVVK9ny
7Oi2uG633JQPPkhYmwZW8rD3TuqrnVwGyAMh2+9M9+ENBuwoyL+8u/IuO5NebKrw
7tdeu6alde1vrGAs+rxYCPYswk2xlxiKDIV3H0cru8lk/BxOSAtd9K2c2Cfkwo7g
FovYPbS90OUej5HMQXvLEFf3xDsDB7RN0gy/dhXsjsT47dg6d/RaURguz8OVuuuO
AHmU310kawMzKuspPUYGlTKkH+6RYiWLYaQIgXAa/M91BJa0MFxpPP2igqF3RYWN
7qs2o5xWGTJ0TBh/DzTm6Nuw2w73kg2gN1lEGcBSS3IgPaRwxhkUvyShSqdhPpzW
lgu9hzLTT0ON3Ay3AmSUeAp2xA9jhdHc8nWVp9dxp0Jj/eSW5Acr7uhbsKSV9mxf
ONwJlmCw220nj/X1WGbkDdEqIk0j2ICV25jGFdAiYjgsIw40tkQOJb9Ij2Dqo6Bd
286eqwVDo/S2aikDl+/3Qhm4t5uYEk8La4csbdE+rheMT6o+QGxCsoXLZlCH4KEc
liM8U3U5y96t/YTeINnTCk/OeoFkGeR/gajv/W+bei4Fb1MooAJlWZfncWn8s/ue
oNpUVFICsmiYYl91lXBIrwjqQmkc2DvrUHsg2iZwkLQ4u2gGPxod835ajdWl0990
7bOw4RWLVbQTV8pJdP7X3XVNPqLI5MdKsKTXINLGYYgWbGFLd3Q1S6suzhfFU88Y
p/hyx5gHIKXdqvvs/G9FeKh92qGXUsoX6Emp24ix6Smcz0lCaq8mRtT0CYsYXzvL
thP+u7rs+FVElx0RbA2O97pmhpAWiKhcEWp087Msi19T4obIBoaa7Lta42t96bUy
un7Ejy+Xv8FYgmHHVNJ2F2cuTh8y3D3Nsqw3NRIlMBjDzMzdbfw+XcyZpHfeyEe5
sLAkjArRoCGvZYJohS0xZCk/mLrr8BzSaS8n7VuIII0x6od/9NuMcE228A1UDfDP
SEz7Q7UV4+8maT9jlVkg/xQJRYzf+bSzchN0JxfpzbcJsA49kjRpmb6qWWLqcHpj
dxAxbkVEmkLvmrBOhXaWN6EOHSlBeGe+IFMGCp7Tqh2bpNI/ClgD77xbkKu0JJnS
g7b2JarBLWGjOYGTbhZUyx6Dl5/bprwW4EbBUxHMKXZPTL98IhhJcBUcBaDO//Vj
41gqYCbbVPxQHnr0SbkEgqQNCHORxWjrs6yifhJq4ltq3dqfnwF/tdLl6HiG8lmg
HeCsRPx8GeVUlEdl+O+Rlw2AmGkTWcUkMIqvq2CMLhvAdHY86kiFrwEgt1ULWAWh
q9BvtfsoLkfnXrZjrJ+/wresiKS7F1TVO/CXkMPpXiP4ON+ezBVjWovs5AxJo27u
o5R8N6YYyDbeMlFU+qjdjyLt3XXQ0YTdhahIb672aC1EiswNW1255YAFHx/M/DHf
U+Dh9e1n+eBfb3LYNdrEVE8zQxAYaPNLbsYwBu2Z1ghMi4R6QeRW30PbIBT62kvq
CrTci5OfOw+za8DVxhiM14ye/d7UghCDNNMPCZVS23LhyIXhpL2IBZUbda0+ZQSR
nJh/8kmdXXe7eRDJ24bhTodnyp9Qw8AR3tGKj360pjPoaucjbT47iDnN0YOp2P1N
09bOB+iWvXKzGNFOwgq7/NgVf00KfkK61qLI73SdiuoEyN2iiTsi8go5qRxgONOM
3nwz8Z4XMHT9Pm5bcGu71TBxU+9hqjKfJ2GQb/cb+sNeiazV2syp7exiqnn8b11N
o14lZAPWRjECX0tQk+v/Q4+gchWPWQ+a9tvu4nCGWTm/fudXPZPukfxX9cSxbGDL
R4+KIExxJbDBhacvq1BaVwsRMhy68zcv+d5NUpp4fTBBiPPyywTbvAtftKhOKPrC
1vviZdOVvEJI8XJoJGHIdrX0Vvb4hzl8PLLUvCvJs+u11f+gZbdtXsicX4w3l5s1
AzA1NOzhMm7mKFEdAZN5dG0O16uiUHypj/wlK5zVua3L1cm+YRNzNhvEEkoaB4IE
efqP1k4rLKwPuQRYryMfBLEqZvMhPypxGGumfJqtozVlsLVLusN2O1ZNsjstRNZz
vcXAv/ch74x8Kq5hKxR2laKkdtw/tyjv/2Ldex6VXZ9ABZW6ULanuei//p1GwCRb
2/hWjaKE2yEafH0floZF8k+onb7nKslF7oQZlLOIaMibiD2OzWLmwT5LjznyqEuT
c6Wj38BVgdb51/Zw7l4GawfnCq6wPZflfgi9uTaW3gLS3QY9ODwPvqDB+zPHR2e4
oc1onJO71CSuu0QUrrZ+LiE3MEjideM7/qPAuGr3an0AL/15hmEGow4Vh3ssJ/2J
gKPvbVfdlGxWqoduSecz0iKDEIjhF4mGB2v3LPH58GpglwzCG+QmGdgVO619I9a0
9bHheZv1IpEHGY2q8wgzi/oNKZeyI/Hpj+OHq1symG824QLKDcgHWDG1NBTR8btW
vx1YFt6MrPlqJLpkAUKwGMw+2He7GIsVxb07znztSFu+d63q3I+7/GqyiodM/zkQ
79eOunbxzuG/D5B/0z2T/u7cipEuJveTzG3zMOjFYh/JD8clbOmXjCRSElxjJbU/
mZ86zJ0aUIV7+SRvsro7gHiqB1B0zfF5VwgVZi11HaZwL05tYXq6D93hozdR6fnj
FYfFf8IbmanNBu694VKqEsAfky3p8Ur2QO0TBTzqlDu+c3FjNGh10sujOK1fKOrM
yp2qSEqT+Xv8SB3z+p2CuDr+zDPuF886BgTHHnxRP+/8xlK6htzbrl41Y5wBwbOR
4AaVM/uDCILZAdQeo/dH0b1U0QgDIg12Vlj2SEl0XewnSMkiQxuqSmvoGzXqf67i
vvoTn0WzICVrbV/PJpjBzMnRxRzBA6ictUdtXRHQPW3pELtifBLNkNqK7dEqB017
iDnrh2wumRSzCP6rnxkYmkRpQrGNzfNnZY3MX5jRvGp29Vzo4zX+1MKJ6Vq+Odj5
SVosgtk/aAHNIAK1w6fUp7YiMC42xFnKEt44F04s/+Y+yNVfhJ8O1IKQLNyIS3zJ
oxd+IgW7B5keXGN0vhfXLE5Fl/hgGrq/Bmoiy1xAf5yH78iTMZDPPwkJFxH4Hp5Z
e/0GcXh0KjsSS4XGo+3aRbRKh8OZLWPNnujd4Cg1u+CwIeM0B2rCLT3hUYM32mfo
wiipPwLVSr7nYQLcPpnrGMfE/ue17NCCbEk9+KTliBgR1hhnEQBKJFEYOZ5K4KE1
porQIBmOeZVlPfOnV69uqEWBXa1DBG6WswBq1DILVAd3BSkBJ5oYmpFrFeBZIh8R
0Jh1SqAhoj06hILA08Qzb0HlRMFSNPWntI+smjDuf9j6D5/nyVXUVUGHYvH2o+Mb
qdy4ajv4bzlZYZa0N8QYsrKm9FzeqZwWDWqTdIZCRMZfKJeB9EJjq8YdzZh6vpBb
SCR2vE68I/JmgC4XTDdzX+3AJIAJGiKqvEdI2gOeQrp/WrnYeucnkDL0jtD2Ri7d
H3KwcH6K4NGF8KJtDudbPlit+jFlrv958VIfhMwFwcWCoucbiSWqzY9sdhvBmhT9
RO/8VaXAd7IqF7JAQjNcG437Cvz/Cx2lO7iSNetgCjE5qtgQWdZ1l8sf40tPlT2Q
si+saut2kqpHkUi8nCEZscnwTCbx/cc/uBny9i2NL+rt3o/nBbfG1GXZ6NxD/gQ1
2x5tBmz4oWLOnVYSHZjHE7SOGfZFJbZP150WIlxwlAqHJSbJadgq+oWZPnCATfep
k6uQH3G1lVDZUy+r/+w0Zq9fb7vsaR06fvB2XDsZ5mmIVPvL2YYMpPloJ0gEsEOi
PsZvc6sq/0uHkROBkO4XLO12134csJTfAJAwv4gcvMirSxjnddEKg8T6F/thAM5F
Uiugn/MIxetCBjmo0E05u5iss+O1UT2UsVeBkUVZbvQZl8EysnIEHeMVpJS+99pY
Nsu2f3Ud8k3ZzBmO8oGApjTz48Qrhm/3XMfHGNkh8GFPmVBiUkxIA0YqPmoLYFKP
RmY8W9tj7mf8v8X2N93VNapV4DruLs1PGaLALpbynevysfd+7MEcXJyn79dOLKn3
tPvLs+6COY/ZK16xRTPiq2gEajyij9VYQA+YeB4IP6P4AU60aemDj2bQET2/2bBA
i1UeZxuUvTXqqdIGgiv/p1HFNWWuWQw43b+HTvibJLngc5KrX+DUDFGSnzDRNj4c
mCaFdE0Tky37yz4EDNOJ37/n34rncgtfmYsQtAgB+B7WVgiJ/1TfHCadVh9iUJM/
zashogYg77hIOVveeNgzg+qcPLRD59GScJjEZ6kxPaRvXdGoF2pfmbE6jFZlUWUZ
XKUeSZTxevmtRj4uXdRBhmIIcQUP/07fTRHyHw3udh0gF3nkRwYn+ULeZjKXgkgs
XJSLmK+zDJ1L8Ne+VIhhNcew1d339JMVXDeM3qfO0R5uXO9mOAJozKzmdOvj6L5T
ahEayMiipMVnxLYmbNDyabMpXFugLeTUaMzkTs/g+541spT+updUsU5sYik2rRnc
5+GmMFiuKqpqd4tHpgh6+5xh7er24doXtQpckqhXbNmCG+FxvL8R3S9dhE0szA99
ZDGFGOqv3WPQ1mcCmaxks5MaKMmKNBIontXRKeRCATkCQaC1Y61hexP40xWaQlJj
0QJ+HaSeds8Ogs0ps5v/QSL5atqG77Lx5xoHgDH2O983PMGWYGY74y/7vdyMi7iB
uQ+BCBZGRZUTdhPEB8vaBGKbSg8Qtgl3JCnfwp5n0oQin5kFL0JWcO6VAbx/6OxR
QT0v/vRjpMAf1eSLBkC2K/+aWDOdbPuUauOSiE9PHr65Dh9PsBOJ8mI24JrnpBHZ
CMZyEv85jwoqrLYjS3F1tBB0pWVumjRTiejX3+wsWYnUPqCEE8mu4iLWODo5lEs1
sdENmWBGHNjzldzzxy7OhdsyMGUGneoHpRllbTrLFW/Tl2tx1iSuQ98QBEWX+L1H
vRTN+MaH8bby2/+uKVVkOcg6QhlP9TYLQvtcDxIE7AmI0DJfkg7t9Xy73y38NHax
Bwk+D1cS3RB+Tj8uzYXDbFQREv8KK0nw+QXyFuCKr0mhMocl9SNECYTY32/yi6dX
mKgaphW5cx+g+ArnDeUVNaC84OwwqQee9U9ghCvECp5ttdXr7KA2lDtVXXqEQ12/
wYQqg0ftgpBy6Q+0KEYeeJ3PEGH63QzQ/czkh+WiRAPl5AcxLNV/ahLT97EAXV/P
lWAYgp1ZzFh7I6ZUuN8QsUVKVMenK764Be/CkgLD665WXGR4dngOt9Voyxx2tCOT
ks4qizSaDIfzZIPXU/9rOF4i7cQu21+WQp03IXA/dHI+ndU1S+kLD1UTzpOjWLu0
iu1iAumTykZwuqy27iWX7Ww/YKn9y+iitazkIlhCdG12l7eeGxTRiguc3xUBYkXq
OwKL6AoaNqgFD0wExj50mCFqRNezCTJUxkniPqHq+NVbmI9mfKeCWPQbPgpT3mfN
15dRtxGb25V/ySXtIA3vaXV5euXq6lLEpAhLv4pGyq3xpSsB0JpzxAY+rveUZ1HR
Dqiqy0S4/4MI9lHod3uLhbkHJxl7CzdiUiCk3+jtjuVrn9Srr8Pk8+OhGPzKu3qJ
w2NPMj73th2lTLUrplgdBEONtMIWf8t/SIOqw/bqn6+E0JOYTK26R+aKKGAstFXI
bLX9+cgmViSmDkTssmK6iT9HpdVT8YxvMKvM5tUiQm4uTIazAnrkvMxOdYMiUkK4
NDr1xsb42pzTyCWBlwOI4goWgMU15mzvfvZgMxLpk4dZl/PKvZt+jQLhNvX8IAg1
LEXmZH0XmV1KfRziqFMU7AdbtxAknoJxMn5TB2wc2KZMh6KN28+WtaiHandD/XTe
JjMrxKVcZBuwCfe3ZHrZdCG0H0MUFqUo9Oavh7ncSpMa6d84oBKciDcX+XQqtaLg
ko/HUaiFFuiVV+z97HxdvIaHBoAwossaLp6GSTX0KiFr5PGjN0uQ4/aRpSrTi1o2
5T015Qbag+pj6da0rS+IOMk0ypsUM+w4h5Rcy/5I5F2fcZFROZ9KAUn/GqQ1D2rE
yCCZnyGt8FDC786sRViA9pK0vlnf9V2lmP/am7ByCjCCtzAbsTQ4P2kbRdd4wXNi
JuK62xk1V4CtexCCHeZGafWGk5rvx0qZMELM5OwuWwDNmgT1YbFTSgnU2aTrrfWK
hyCogIXEnmsFYxHtEUg0gqh20zBFRry+l/eaK6/eOjRxxE1FdEKNXZwq+IJTmdZm
O85cCp3eVPdw0iIMyofukYzOb4gO432mMBHcPNd76bes8iMYGQR1Ahsc7J/GEpAz
2T+glsO9uIRS2y5Ws6Rm1jvOOcFTddI/oKUgwiA8ZF6dSjzgOTEOCi6dMRyQq8hc
4CIaeYZLrObGa0p7IphwPotXpd9jdaxC4lZ+i1xnscaR48S94UUv0xNsYT8lkrnk
hHvsSxpNcSr4ysCLjEb4lVO7HZ5meetpERL94NyY3azlnz2lyhJ9dEfAJpCgVCNO
Hw46mM3TtAYRGTV1MnqxDRAa1vSgCOblgEr9NGqGLPzCGObSTqPjx/fI97emrY45
3bSHhKdGvfPhHXgMev8eFmLf5grjWZrZdIgCMvs+AW8Hdenqt5QEJOLIqwjFsyTm
8jaCFxTPj4TB0QE2b4p8K3SL3DUyRqTHPsbBivPQLtpSGIWs7exaBlZl+0/LRAbz
fD9WG2LmDAzarjXwWPUvcJPXqMtsUjXS1vokjIGJ/Glo7DAgD/QPpBEGeHeRfYFx
uFkqPtNGTPmKStw+7L7xlhfaT3FysgRG6NJfChs51Nh63ovoP6ilINhvdQmro5ne
2oP0gY9btfvAGZCbUqfEutFmKtpKApndlqWpi+tPQIEOgZIewl9BSh526YSpmOnk
xW1kyujAOP9RpwM1TWG/YrnK8NcHktOFLGl8f00lUVDDMLD6gPS4PhzzIAPMQrBc
sXetZ87g6BPn1Q6xKZtXVzqqMsJo4cA3qTLijMN/WVD2JGI8vgzi2Te816GYidJu
qMdiO8DefgC6/hKpf3i6Cac62IfjcIXTPJhr69oU0yfZBeMl2eHCtsOGXRejXtEy
c+H/JJXX6dUOGQyCIGrUBFLlYbonae9TzJJc0nhvS0oeuw3lzImpp26HJyuY+6Q9
E5mo5oAN724M+9AIYCLtEzRQq3hGuZ2WmGydlF9aJJR8Cpntmto1EnKIg+diUzOR
MSFyv3OdFM8Yy2cA4p4H7LgK7kKPHW6owdtvIqHvw/MT8wOgErj0PUuFAxdlAvwr
VwA1hPvFGGoMwizRWsY+GbbT0TKqj1gdSISYvhBjHwkIFwHOht4cYaySJ5yyZROD
TQLMkqMQtZuoVrQC/CrMpqU5ibEtiULd9b5FZkD2mEngepRcj/BQEArjReaLkKIS
hRv1NUdxtz5VAWbwLSjBgp0VNEQrEVmJLCoYqPnVDxLakUgALO23WYN4UatqtTDg
OnW7RyjfaR0LUI8cLaPO7GYaj58IWSNirH34AcWmRaVkUQuyqxsjdqVWz9sogZxh
k736TFzyD+3sX9+5otCtF82rEPonJhMB7D5iHc8MKmTOEdAqphhY0CxaiFJIrXj5
5+U0Tl2xUJ1nYwa14N2OValcD/bF2KPtgpKAULHgudgRumEEkuh0mF4SbXOBWnvh
C3PheflpzFj57kLEDfecB7ZTJsWkBXtKEF842hPB6C7+coJDRwYkOlHaHGI3yQkX
RuH7dT0xf0S2TS0BEw9IpzFw4uNPnMLIB4tR8IaTjvYu59hy9oXq/RgJ6P3L0roe
lTvCyCT4HtpNyyaq+JC3Phj23eS1iuOInlKUYE3iCeM56XKzbi+JhYkbDnrFknH/
pwVqZQL5C3fUtIKpiq+OOgD+c+ynuzSUBI4lfvcRw4M4WeZC5h30jczHZSpez7OX
tXeve9O7UsXlQaPE6gBqCgcewMg2mx/z3ME4TQR5R5aDCc+SUW6gudJBt9DU4zZJ
B74S4osbOQD+C3bPvNjk+pgjTPctS+HdcUQJBRg6QFUOF0gtQOo3TLg/AL78x/Op
scezbqnWuIt/n6jDxjBpVIZ8pTdNn9O3PPusbuClvOV37B0QoixKOviYFd0aWfnO
09bPZ8Szo5/3RXpsnBbLCUIhdFscHFEn8LV1mggbBTDdTIMk9ftu4mUIPil/Ahgi
2RlABhdMcC7v02mdoMgR42jjgyYoJbpji9U35zaHUTiia620jUGYiz55SfGqg3Rf
2gzhrE2SB93voxnGNQvhoai1FpIc7UWtKVnb9aVWFP3Q4/0H6SpWryFGfXYngoBa
fiElk9N9kWxkXBJAVuE70McqWiqjWC5mUsLd4IGzVFbvH78YSziTCD+/ko9PkfXy
SOxgR7AT9waqJ1mAXSkhW9soHnLmGt+5Fn5MunoG2mShosqRWH3EKpV7sebcQaU7
5jhXC1wU6TVC3TqkmAEjLYRLwgXFn1x2kNV+AD+3pc3dmOFG6kbA9JhVLhnSwWqY
XIhRdLtKOy0rRx54776zNkxIg+N9ISp+6v70Kj46jtqRQQnVrg3fW/HlqaxIXlwc
pv5mQTKLSslzrqKspGpVPsQJgBxCa+Gim25RL8yNxYnR3yqbLPxdrEUp/gfsCKM5
zXdchenUt1LM2nUxAbAu3w3TEpiYl9lJ2k09VcslpCOv3XKU1zjo23DB8cRQ1W8u
neT8MChgPg1B9uiWFm0/cJXH09mbQt2dp+P+A6d4CzqJ3rXnPvwVnLdEWcxqtcwV
bfmpqSh75wZofA8o0V6z3lA5q15r37EqkOCrR1EzQpO1ir2mXjE05lU4dW7m3vOg
5ZDBPYq+vf1NHjK0HHjtzdCavAjSphfcuGfmL7WmjYaAtOVNFOyCzrXg79WUIqHx
zuISRmfQY5/e6vnbjzpRazOFC6xvmx0sCjJIfdavgMlEyOJv5qZFgEayy1El1g1C
CleVf7Dy5qiND4Pmw+bHs/MeK3jLVeh8I0ifRgLEqP6L2ykTZ5zOSDoNqyipVJHr
LZj9nmT41BF0xv+41dmr9AB1RueUaaZ+aYX/alINCXoLZIl5TJJkKiCMx1UPKcDO
uBEPqQbfHBMifJbviNgpVsJ6GHztVbQElDpsntERiLq86WokaB4Qlym/gzE3ElRy
UHwCOj8Z6zwo0+odtpAsBm1Bhf17lhK7XDqeU4fVteznC2WJjtfaCvLHNIDxR+mn
+H7VQfcL7R9CGgbM+7QZZOthJqMYjoOEbd22VDSfeQnFhftZ5AV2KSAeK4Myfi3R
Q+JaMvTaUi3/eSj8q0i09h34gEpiQAFSr3glDhhe6TnPJlBQuscQ1hW82qbH28YH
0+8JdgJObpKMXNwRjwhFync/ZRjnAkFP8lgjKHpJHaXvCVH34ijfRsvXiroNh4wr
sMBuF1mb/l4Mdaeq6lbObTkMf0yyPNQcYlQlIqbKmQFyLmRg1Q8KycccsXfGH3M6
RPTd41VaA29ghtRW7VBaSwrU7ODmsWgMUAhyU+SVCLRauPGL8+ETAChJ0fwnyGA0
DIZR/4KvW8eyc5PMa7KZhO2odFtdjcyMiH3JdmGlgJQkPXtHLRonsjMEiocO7gsI
IgLgSv6wnjV54/6hsMk35bhPkb2QxedCJRVCrL/aMOwFUUgAboDtH1gmMnZRuO2n
+BucPVzDUN9gXx2XKGCPPYlz/LMoGZgrONLFEfRUMfntj7XdgJDAUwwOJM0cq9Du
19WRg3h0K/PFm5PT8I0bUAoD/Cd1kA5idVzijQu8uTwKo7sSaVRW+fmtjDzmRk74
De5oeLN+kDc+AU2gLq2KinywIufHEtgsHbjvsSJ4f11L5swLuP3lBoATDb4Kxl+D
Fq31KgLHRypXGXtx1zvt4+onCGlJdL61He6roIJ1MRW5zdzp8Y3zWXXLmiSgY83s
NqZmjZnGuuMy9FIiylTQBazfeNJKtPFyYD9Vb8f9cnfdyvVw+C9XhROSCRCfmpU9
cT+0HCx/RuyZb5Yk8/2h+Xv4cIvdbNstBl3dVSEO3K0+FC1grEV6eSaMzwksddGp
sdT9e6Z0qOAovg0i3y7UIe3TQBO6wfN7rjK9pGny6Gvr3t8o10Nk+II929HfoHO3
OUZLmA4ElseOhQep7lWEqhQpH11cOV8FCGOIeJfFXBindNL9sSmPDdpIIQkP3xuH
99CzkNncaK+BcO/6lGZvfwAHiYJ+Qa2qVlNmRGF9LFUfO1LLHVtYm8lV7SN3I/0I
p1smzViFFYBI1U8ztDhKO+iYo8dXpmatQyLUVEKPDU2qcYTPCeQGrZI2QGt9QYiW
lb5Xz46iyMzfpZs83scDSpqQkNi9xVMFxhP+vX15oB+UXP3K0tIMODW8evKVFRNT
yihDbTuCJD7fdLpbfM/xIH12Vx3r9raNzZpyGPNAkw7qMNTLWxseSDR0WyVnPLr0
QdmOhIUJsLnWOYQOKT7FtR++zCEUdaG9HoLFhDKd00jSDxLb1NZeKzAAO4Eo+3U4
itWUpMFAu3pmFE9MR/lSmkjA7tKMdJLESACUA8ZGC9JTQJyD11APoVtjr+FAd1IP
py8o38RwY8wvCMwJcJC+5vtp5VVNLoaboRcXEVkQ7PMor7HIgESRYsvzxLO10U5t
7e3h2qwVDiY7iPi1kwSho7ifCp2P7BcpAWWDTQZGEkXyGx5nKX2jP/pxUT1tMtR/
YsHYyoteOFmGOMOEYiDgwUYjkz9O1pTr4FegMVScZNtu93kNaGEHss6/mjeYHiM3
rIVahMy9B230HLjZx5zNjizhEi/7nyHWqzEvSTOUTYB6a+0wyIDPBIwQbgywiuU5
ZNpib8n99pz0LgMYhIcGGsLg52boE2ZNiJtS6LDa1/bmMD/GPSB4WDcdAJ4jJHEv
nXYQb2qgUFRd3tuFKTOpb0QvvqfyPZj5Lr8RGf9dN6fORUS6wH0ceK4NOmWfks66
TQSYdwgphLa7PlxucdqxEqEYzvxHbbkwLGM//+aGQ+OpjshTmPMLiZyj2uFmEKug
WiInuLqjuMWfJhLNVj99Dt95iJIj2gxC1K0KLkceP/M1ilERTMrRQsuu0uPv8Ssn
lBAxcL9hyJq+ZwDEjqYzVgRNcjCAf2gYiJbw4w5j6yJU2XvdduFuDqJJ52d5PIOX
24Uqnb2KNVAva8UjzeOn2ZQWOz7f5iCumoydXhsf+YtlYtJpWPt4twu9jnLHnB6e
h1ZtUMhVFDzaqChecXDGbImEQQmTDudrP9409yr+iB2EVNWRNLiQrxda7lHNi6Sa
Q2+uCqMjTUrk2UUNr/48g7zWfOjIcb1z+MYTfjkOUy8yOUm9QZ90h2mSwQABrHAA
HBeu6+5r+FIbyzVRa2AgbJIot1Pvu6n7rabeYTVC12+RFFjWHlkNPxhDdmj8PSQK
O+qMzORlQSDvhf2aS0rJUQ==
`protect end_protected