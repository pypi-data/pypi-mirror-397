`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
I5JJnrdmdIVaCewvA2Wm2rQAOEaynP/rksWXhWeRXk1Hiv9MuBSy0NLrHmKsRxXi
Hqc9AGHUztmoF2eeTqZahmY3VKtAE5IuB+os9nqm9zWqfnRay7udiSr4yrQOmdca
xtSHRO/OwKpCe/4DDvslI+gNwdnIb3WVGb20S+in1Ca7la5uscYpqsjzoFu+6J+s
CPDBTdvQrKhv2kb6VViqaBR6L61VDu8Yc2n8+siiZ8rQa6ahvnQDfRauAHRyvrAm
ojbEeKV/NNtQ2tcNEby9XpRi8e9BpibfHwM5lKA06EP7VycIHMYTzXALEncfrcIq
axtPH24ayAM0Ja97BNtNFVZSKnFsT2Lbi6S7hci734EBKkfd/NKbwvx5D73/cEPZ
gTATSvLu18lysRaoEke8BDbXkVBMRw643ewFRd0liwPBQR1o99FSWekd3Gp4T/ZS
Ig84AxfblOufHno6onUEf6FB2jNF405HcVDz2fNB1C6Lzxnb+WbwfYl+VtGwdozx
7m4LPD2wKD6MdZf18wgNvsk4YrwLHmWRmtnebI7Mbir1IabWA2JrUyW8Nye6XPBW
7WBXwIFE2VS78CrzJUDFmomFFB2jeRJQHFF5G+d3WcKajx4b7ibXM3cGEDUBikll
YVwr6aqsE1vYh88N/zvNjCv9FpVD+4KKZHOs7nsLnupK1igxRseENK1t/PtZ345r
Puey6F7OBNX/SmfoxpNPesaQvigt+opfx4+T8wzhs4uk1mc6s6pB+APFc9o9xcRD
bBiGohGpiHcqoKTcCfNXeP7vi9zwj1dJ67mhCFe1ahq3BbBCLfsxm8oNSX/2ZNuY
jTxwi2NZ87peMcXR6cI787nLIZ22JumFEhLIKVBPgWkdnfWzdkTGQuv4n0X0LrXI
5XWJBQf52OixxMunwSCg6kcmNOyE+vl5yh8Me84ojAitenYEUja1P0OBHeJHzU5m
gFuyIgRQmQo13Ndf05TcPI0RkOC/JM2OSigknBzMDDrRfpQY5ze0kjazNK0PBs9z
/P4oocQlkldncvNAC29cmdr4pZiRffwzZpR1WKFKpMFmLSfWvCpWurVgFjUZQa/f
ouL3rPC163ve2qUmi/xv582K7RZM+yzcny9q5ECLc1EQyWmU+NevA8+92Cq+IvnT
y+DqReRV2a5Y6/QZlZ3LiUbOr4FeZ7qCmio2IaoeILYUXBxI2DQlcVLtlxt1FGh+
nLCo1GxVD2NHtzazv95slUS3Q1yM55zwCXM8AVPrfiOalzhJL/2Z4AtOJa31Ijff
CD+GjQgEPQvH15fXpmRb4b/qKZUhMCJa9OI5/nkKCTvgXrK73nrRkFhvYsygK1zQ
wovJskWAqSueR1Xbks0DN1G5SjdZEGJU5E93QGJ1OSWqVbw/nCfMhm9qzrXxVoA5
YPUUQf6o9bw6A69+mnWB2GgWKMSFWWbQOxECznhE/SgmhYRq3hbxnufgx2CCPSVR
OoVIWrb3WYqQoCj8mnGtsaDp/y2Bd9WfaQ6rQWbH05cA2H4pYc1xKjAmyz1iPIku
OH+67nEE3IqDmTpICVfLN6nf7C1CK6uYVgytNMwnsq+sdbd/kyfHTNawl7ReaDfQ
U/704HZv3TjK6INH9IhEqBH/Dzq3+b1FtDd6hibqUyxcyK1nbM4XQP3+LzbahG3X
jP1aR69GH5z0yWrhAspIyKbqouyUKOLNa2wwx2uwhDJ/NRsEQ1Oxt0eG+wjZjXjt
ImnEF+TkrZF4Uggqj9BV1pm56mj+GcwknncxjefRpYal3xgrOJQSm5IaDHfKKZVp
ruTyfPD/RcNugcjR5E9JNYbBzHBWj9UJevj2x4QMS3TM3kq7+7379xxbZ9SeimDZ
7HVOXyTtSvETnT8C7L2RCeRaaIHR5C0vV8sTPNBH1W3cuDdSCOA+qRaXAzxr/NOa
Cn4Z0zzG0WFTlEx7FUhWHjVfzx8qEXsb4gJ5kEWFX/XdxCs8cXjj+YNme4Qz3syQ
ZTDitRjwsXxudbwjQw2L15Fp73s8rFWg9P1JOOGXO7+W0zHGNprXXGWZZ9+RuJXO
Umrkx5AAT0JMxTIlwhj4Jg3PC+VdVhblyrDzfWqsDpimW7T+ZlzGFBiJe7qZRVuY
S2xTVmCMdQaiEGyZtpGW9kRYiJT54cuHve8hbyFrT2g=
`protect end_protected