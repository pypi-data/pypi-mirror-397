`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzUf4aF5bC3IgM/qW5fkpB+/qknhIJ/vFdXfo0jO/Nqf5
3sM936qPSOaBgSER0wnJ5HSx8r9ZgtoQV3ERrRsSJoEDf45ivMuj+I6kVtDnIzVG
MI3u+joUT2XFW9ENShCbfJKtf6yv7NOLaG7L5YJZv1LNHSSyuV2EcwHP1uKEjv8j
CVZwKzpOerVZgBan3ACiTN4Hm5ieZGaQ5cQIlj39bLs6Wu0fxCMhmlYYFSQZFq5H
j1dkwcw+UHCmJGkBBt6GN70e0267p6Un2F97SWq5gGkZCzGiHSvPWrGDQRxg52Hm
zjkIYeWOIeVu4g1KjjDv1cZ0b6nUuDA/3RenqFRpkws/zJuvWNNObgQMPKydjf4C
uSTo0iYZLotzaIKsVrTTbGMZjFFEYQ+MhdBYpsp3CzpDyDYAVOkjfR6WBDTHq6il
JwlIWAWnZiv3wkUNbiQSrzwD89a4hmYFC8wa+pK8bNheJQaGqgUNoPms2X1AR1Kq
34viK6qgdICJep04el2hg+AORiQuw8f5C/z2cxBo61xsvwYtbnnX+0gqR6urlrwr
SILmnIBVYUJm7pksxxe2jRqJPsvErKqsNo3Q+hyt5oDAWuZ/syIS0FWLMtJ3/MrS
+vFo19EFjEDuD2oHYk/5Rxq041VD5cMPHa+3ItE69P9nNqDFOm1z0353z9essPnr
mdS0pdgXZobcjbd8gvx6u+IktICyGcygpzRLvH9Q3wmgxMijJWgUa/Av8AaJlQvI
0CpXe6PAPrN7lsrwAaNSlgWLTuR0nWCmiYILi1re+LmE4PotuQMp/MdVsZC2UKdM
ekkoRraHxVKsTnlYSMSfP0sN4KZevkRW3TYcTWl3JDp1krHaW0VIvlB9UGU7nnZ1
rkqW23uLDiA2h4VsfLDR0KDyq0lQ7gyz5krb6dX6Ux4H/RpOAPjfLgMZ0vHW+Pyn
afTXrL6DNEoVNujNZCUWazKr6o+cB6xAdc5XtkooOOpTXzBG2VTprpZmwUDhdH+T
1vUaX4xwU/SqDNCFPqhhMJhi58hFs6YDbCMyyyKAxJ2GlCEhplXfuqMrCmlWJN8V
URwxQ0NiiJQrXiEtn0JZuTOSgxhHrkSZ9kC9qUEf4wLJjujPxrZxmuWlAuNJpQLn
5zYDcUpYhAKYoMvYVT0T8UcY0tmWRrB9wxMVWjHHkkKRbJoauByyA2SZTfKGBX8a
J/fq0AlkWG9QE8eGD65lngOgLMKpTuwJwyh8xKYpxQ74ClV7WYgjzBvY6yUqgB7P
Ssn/VoPzXrtuBk7DZtU9snC5PwBQLYwzQFcgmCgcbKMgzN2qa61ROQ8sTOsODQQX
IdKc1Jqjrv0wUa31URzdV5fsDf2v7jAB5AKyTvjzDvvQPMONFK7Cd/aGvqzmJOI+
4P6BrJPGH3V3x7Owk95RWnnxz2GePTrsxUC2dx60N3GiwbFGM/nKkaf0r2a+GOMP
1hHL9zwdT0Mtknj2TLL4AMQ2IhH2HUYKfBpxiAj/MJGCprcfy+u47kZKVa9CPKf8
eJwLSlUQ2CYwzK2qbdZS/kLoiE2FMeDkvLgoro30UNgwjQrmW2U6MNj6bXPcgeJY
BEFMsLquhHGc8HWUloiAUC1n++D9CNoICBprMV1+rhQKl8KguPwPkTvclBKBdysF
AXUhvA3bhYfzPZAjspJWgvnFhOKCwVHs0WjUKRMC2jr7mVbpGA2tAxpPsIqS/5lJ
sW6f1gg0blARuMdUskiH03xpGt8AxAV3I1pgENbJ8EOSm/RJq9Y0uIdt8qogTqiU
YAafLBvMoXVSKryZ6SUnXrPrbZ5fds7kI+hSQ+D59BMR+lh00FdM8gKkSojC3WWk
r/iaJvc5oELh2QfHQ6gCO/HoMYES4QfHB9CudGWa18aYeIux5++y84e15FHCvrVd
fwMDDo1Y+JQK3MvFsS0iZ4233SLjynpovFx7t5gqmvzj7nez6XDqcYEv1QVcxpmM
ju0x59IroV6vvlFBhzsjLnDVVv/sAAqCiUwFXinYsCGjE8uINCWu8RhoM+tS0WyJ
c3XBFMVCRCgqCrFH/m9HblWRoPgFeKtrn7S/fgJ12huRsIVQ2DcNLtPq8nmftYTO
JeI0qLXGtGHC+cZXw3QJ7hbRkiynyGb94LACa3uwVPFsKm1i/AMJTVAfGRyyhC88
J5qZ8LjJqXO8vqVdF1fxSyBZwfEcW9n6VISmz+bzJDlxHwLSTT5DBiD1HPmn09yL
X3u6y8Osxw9Wp1am/nQz0UaHO42krq3lL5oEXlV0QW2lrR1N387wMaAy0iVycj73
G4q4sf9b2eUQL0i3pgH5cQ0XIEJw4+vBb2kdfjsqPQOoAg84gUlZhcMuWdM6pwVb
uDO+1KPRWtx5yBjrALi5RJ1AB+esQakJkbv0jz3lPc+foC7HimFE1gedkUHTqzbZ
0/pQ/PN7qr5OdqkuLO5RpVMZoO2SyspuwVuL8Ny651cPYyZnZPNcrmMq7v5JhKxW
xQ0c7HDmSN1pIa80rHMOpK5LTntx8Y3x7o+N77FxI8PRJ+ozJ55PG1KRx3R8nsu7
6nygOUU1KgugxEHvRpz1lD6LELkM/ZQKb0kq2wHaYE7tgD3KoKKdN/zFg53tEECX
aiV0tB0QwGK4XBiGdvCUgDwfGJuAIrMl8c5ZRJuch3cH3amu57QX6n3iXJySjP/q
IupxTLqetSlUAj2lqj90UJDtypi+YcDvZMCmH2bOofuqrscrXqLWu+jAw/sVcVnf
G8Zse7hyoUHj2bdzonk7DSLUPR8M8WoFbYbWahx7v6TskkqXk2RudZMXB1HJU5l7
Kt7TUuZslXOKwjVuMQv/3nlVR7lENT03tDwn9ElGPeVIREPZpiXbE/7PrcCHflAw
mz+pjlHB2fWi2pmeMh8yqKg8fiLygOROYgSu5bdhI27qmOgmeY3/4lNr50swtwv3
x8skVx14W7fZlLbA2248io9FOp+X8qiUQDC8PCfyKeqsD8nfei7nd2oo+GXLGaxG
HhOGFkcr327j7bwh+yAwuGXRCD49vEq0Lc7duQ/dAPXN6U65K8V07h5HwPAXkL6q
g94BYJZFQGSPR2YcADuKvuEQS7wMvokzgOXOkfUKabeNqCIuBHKic8uiquRMr0iy
uZgxkWZIYfYiIK21YxdNGFn3rMC1EU9Jldf8jm1O8hTFGaMclw543gqvUHjE00KO
GPk7Iqsv4k5Dv3zg3W62SZiWR0Php1mlELRWnU6bpSZUMQ+eotKXDTD7apUsMWYL
opZNr9uGVKA21/scSel9oh0aUF5qydqx/yMF6ZseUUzOCqsDAh5bX5BZwMPVhzX8
AF9GcQSpx6VdmMkin7xr8cxrZilw3NcZTJJ4bSo0bRTdV/TA6vEC2P+653gBFPe4
rA5Zav9NGkzIWM+6LNo1lbxfsUzKFyu8aIw27PEMv0WVSImAiafKqVRfayiO2XpQ
gEoxgB7gdjQYTsZSrEQ6DuJ6BFxk4hZugD33peRaLrgqg3vF98kl1XTKZ7RZ/cX8
tUYCQmyhBxGAkJdfrv1EATZ/nzRODILzP5RAmaaEH3KoE73wdB8mglscBUCxLSvG
rjxyh7nn8E6W5VTpsrwRSzaqrm7kS5IjZ5rtCrbcBxDcXZfiDjpKzOVO1dIVSWrm
cghKAPvQBkB7yWKndON9kOpx0J940kl9FyiAC+sF4mWRE3ezXCXnCQb03hbcKyxj
XuNKS0KaYOMBCUVFfYDXoFIrqOTI931ahZf6VvLEXblF8aKAIcpftoaLUDHeqnAj
/gApDnN9VoVCBCdvdDYbPtUjrTSHyptrmeLJHsnYUghvIAnrlIa/00WR7Jj7tlk+
ee6mhUWC793WofHS7Ib0hPULonvRLKoOYxjc6U6UqlOJN3iLayLRJJIIV9xvQtkw
f0zBJZwHcI9XzVX5h7/N7QEp8/IDyWVVcUhAgQggkJEqK9MnoyQ/kKudfWnU0XmN
mezSPyrFcbP2altIsQ2+jo48nu2wExh1E3xpA8LJ81S8F3IBm47XgIsgZVd/APeM
RmDiMMdcc6il2yCZodQNKoM3h7rALNd2epIxEuGBoN5zVmWVJkcgOqunMQjYLUj1
zyLg2f2ud7Z6CbfkzHWjx99D4mQlXKmRKk6a5r+BQ8QklYNALuguobmHGmwQj9JU
oWjHTIh23FzeNv/51Q2xu1ABXvu1DYHjEwVSmqiM2faKukJmyTTXQzzwprxpoJad
BryhliBDCE9Zj3Ho1Gp7QDxe/g4MkCp6rntoKLDvtbykZbdCnUV7dyZAhb/a5U0s
xyf0GnxOOyf+HqOryyfFn6mAO14f/Fy4VLC3SbF4DtPNNA9XTBOPt+3aDF6hJfcx
YQywDAJq4D+uq/zmC9oBqioV1YvUv/t23ToyGLUv7ZZRBgb74XjhIEAklQLNsY0/
LvTauvoBtNmVCWH8uhXCdX0GXrCvq2iqWTt8kqD205e30NZ6KeIlaVhAqBjNdE4a
+N8cDhF/g4c0sMmnlwXarNOU3BKc5c3KmX9MH0QhFXu8wC2vzJdJmqf4KM8PCdNj
hX1/WJvKyHQJu5Tf4BOw/MC/2s8VwPk0neMn1hDdx3qGdq9tpd0sMmjNezhSZJ/g
DkP7TIn2VZvo00by0lYFy5w5UANNbKvrNa85p5XYhAdamaRdHbiBgLSpk2F2i7rw
Md+XR6KlV/fBJr3x024wLlF2cACUNlEe+F8y8RkjiBam87OQwk1Umy2vCkHbFRXA
riZ5RrFvVeapowpOEtIOcVHyiUaImyMLBwSJiGYLO+UeWpJzXeKcRS10JFw8PLSY
uRQPTeNG+0VzKPYg+y2hjsrAi55y8JoaI4fzqrz8Ki5fkuE5ReEa55XNJ7MHgF1E
8Ni5FBC+tejZPy9FH0v+M1UHtAfGka94dgx+RqKIKcWlC6umFjtWXu+tDFm4oTuZ
H3oqIfNR/oMSCdw5rlpjNuexrvcQP+QzuV7AGtny+KkGGbNuognkrSe9cKpkY+w1
5OqNGF5VkAn6DaB4PjVRpsWziM6ZfYLPFJbRIfijnQMfOqYXhFPyi8PZHHmvNm8N
G/wIg+WAdKmikMZD53G1CxHbujBOXa29OVDpdhDTtxR5Z5d3bXZKG6Fbo/G1BqXe
aFvncl/LYydWBcgBUvIxwXB12lt6NrLZ8QhwPw17rGtEXYicinLga3+YLEl/uZu5
YXz2XrfszhqDM/ijq4DM9i7WbS30Kaeg2RzdtSd6P4a7ek4yZ1YZLm6xf1xYchhn
V8xxknyzqWPEMDC/iFNqnzKC/Yip3Ee+xWYLUXGaQVc6FmMX7ui99CUbKrcJfCcH
rVgHiZrx8uqJznPJVOUmdNdSulJMgNq8sLmgqb4Mqg/LOUFj9iGhdZ3uAqqoncev
FwKUqoetNOpGKQT1/xF26nBPAgzhZQaVXP7H+zRyrbTxxb/FnLM0rdqpIQBlYUw3
BRZUkA8CssW8VEzKw1vTmuI7algQ1pterXz4hFoZ2rFAUR8iQnrRArbhGkE5ktee
7bi0uzZQxoxQbxzCbMG9I4BD5kub7aFzouKXP6kAiOD7S9fE3nqCckC4dics1Rd7
3rLEOLxWeU0fRy43dPKNz8L17Q5fTTisHgCshyycdY7iTxPMiL4P4A+0NJY0afup
l5jElzmzBbcY8RbFRVsIHkst+NERBCcXqN9uIyFssC5vMEQHALAYEOrZMGhbxPQB
zpd1pNlwOdwof52mV+gb+BNG5ZGBSjquHwfWzHn3EOr5tUnzdhDrmLiJmxhFWFUG
2yO5W1a4yYxzNCubifwnHFUgCEPsCkLxLdrwG+QnplTGpY3FE0grfXtbephb+57X
Hp9mklu9G4nuxVX+oMhRtR6zkjWIAF04DqCAqsRh0x9+c2MFIEsN7mMJ7fbxk680
HqPZKDv9LB/4OUS0N4h05jeigOTtXFChnUKWmRogGWdleGPOIeiwXONbuiPtF+FD
NHUjprJGCvp8z1vDXRMSCpcbo/kSuD8EYBdb2mR5Fg48QIj+wNrmiFklXiAe4g3X
9d4NJxrIB1jyPreiekVRTGi+Me133M5ifsUhflRDNxmVm+Dc866WfLTCKSi1TjSV
shlkM5WSZAiRka5wIlOePzPOiTJki0I+iur4ZUSwo3h9fW5jWwPVndyPTlVfTD53
d22GvgkaG8ajyWxA6EzgVEiZCfW9TTuPV3RmqQr8voHHIM87lnV8UjRNN67eCMgV
6Q4Hj800cYzedjElHWsKNvWc+6lWTsQBbQqmf46ljUEzNixV3c5Wjbkr5E3e2NdJ
Lahi3aTYuh12ToFmzisXY8bwSNr/FNKtkphSvp/lcolR8u9CeBNfcIhgMC2yyree
wh2UOwKCk3lWUyTDHZkkTNJGZza4P6uA04gvgZAS10M8nIojNV/pgE542yZjxFgr
cpgMK+eyTBBJDlnpZuurJ5gQCv41iaEwzX0YWyVrLy+lShteDy5dyy8jkMMFi2cI
xWf45w8dlN+p206QHpusZnvGUz5twR3TAnGjgd3OFIHQVQZyyeTTVvnfdnR6nzH2
g4l6t0f4SLHplPB1TZZ6E3FYfnnLSzENHUmlk+8bftJUNPtYXrvrXAlMsRbDNqUL
xwTJkzO+gVEf0e1umHowWNaicXWF/C8F5nJh8RhLt44y4yP+Tcjph+VC32KAKZXk
1OMhjtEUJms1M5BlsGQkCC9apMhSEesgVlLN+yFxd51OUPCdnXGTSOmFdN2fkowL
5R0IyckCLFKBtWZF5Sf8eahrRb3yeEDITP92nXClyiTDrcc6EftGLxsFEkGcgofP
DyAEZSuIwmymZDQjjbGfR7uTQfWPvZPUT1vF0+WBaA2vv85u8j9nsSccsVvJIB1o
u1zq+gjalfouGWyNum/md0u73OsfUyc8ZMKfEadrn6z8APi3Tr1/xHxUtjtxoZrb
eSvLINZogZ7xHYT5yCsLulx7g26ZZXvagWrhFYsmveBijlcFZ6PrKK0T1EA9u4Ex
yJwX4ha//UkDtDjhjF7NHAb7tS03y8+atpJXaSWrzUs+oZdoqhcD7f+JXcMheCnI
a9j6KAS/NTaFjWSAT8o3X6FBJrc4lnCwDu574PMRTzrk6rjKzzM5dFoqTneTL7y7
KZIqaHncC9ETWY4vf5YFhQk4etxMRqONCz1Nu/ZK4/rvRp+WgDAj78kEMTFKoqTT
urc2UpTLrWJi7FL753EC4MCftiVpDNmiRRXwDuQSmt1nQQE4/6/A8wtJUhC60Kn+
83kbocQu8bZsoK8vPHC1Ws0nQf4X9T5mPo7hpkUBo3O6Zu8+Wb9UGf04Io0mzqqU
Kcy/O2rl0/bvuBwCPfmZbmw+30qsfszem7x7ZOXfb4t1XFTxvpb2RwQLDUis+3nL
omuFH+g8l92EDzxJnlROfU2mKg6eQRKULAPbS5VD4Ps2+dTzyAZO13mcvXWNbNa7
OhABN8HlkV9Srac23AW71LtHzkDv6IRJ0IoquzktxtCQxQHWrSDCKw7LH3x2rlp6
KRcR8cO/HcxeXbMKyy3WBse8QthOVlKM7R+tZP23WlylSsvmTrV0W8GDhp6SljUX
V1yb6oNLbxAmFFfGRePYz3Gme12PcYrG1uy+HrAjvQoBpYlvOyXcLfN2Rc6WK+kf
Ry0OWuBemKAxbU9UVjPRkUn3knhiuBFHk/77iktVjFy8Ow+GlZwflgld97REw0bm
TuY1efsL0R7MZBC2pzYt231EEwRCgPcBfUkJc2+xaZQaLpjGDC/rmLUnNRu5Zn5D
Mu6qOdKtyGIBEUEnjBJIJ5Q3WHV2BSdn+sarLxmhLdXIULkDW2UA6VJ9asuHH/4P
ICIIR2P9DMPH2ytJt543GwrBeR97nLAIXj/sRYI2YuM0YQZshfK3oESv2NIQuJTr
r0gystIEqxHA6soUoaDVsBzma5L3qAjsPrazI8PFPQHK3Cbyzi28iOpCqYAFQSb6
jmrRZwzx81lh2JqjGKt4/bJmfvS4YM3Ec11TobrfeIjWHrn1Vp3/irK6DusIvmhR
nKf6B+nzFV4jsPMNx6HgkK292zQqNu4XtB6zwt5z4LZk1xdtLVgMYToHaz/fYa4a
Xf3xBQEeunix29+l+spAtFacfgM0p5877NGSb2Y0s0n4HaXy5X9n8qxG1GI6FwzL
j2pueJz1HFg3VdKMuzFed4Dr3Z4fsWhL9zHPFcbbDX7yQvZx00PjIsAOK9KZj+op
mp0z0Cb9JthADcKQH0m25u9aHTkXzyKETd999lC8M17ucPKa0Zli5/MyyByvxuu5
SyvpkWoPUUk4WhTkbgG2iP/0tgPvD9jMCL5t9Fx7zuBOdb6fe6gBFqMdbO7812pe
+GKyIGIFZ5Nl6B8U0XSJzwj7UygF9F4TPPIC0U301LbJzR/CXE67C6GZVfdw8qa+
Ve+31tCPR1hfkNN789WRGqb1bL1QV5TqSbaNq1QhhnmrKHbSMk32TIdVflv7VNEI
JOJZXRKh38z09Qzk3onYB2V7BSV63FGRmPYBeLx3c0cBk55DMGHZOl6cxHmxuFYf
qrl9XtNHgRHms4KkIVuerU1SMX8nxUScRfVmwLDPjKtOhZZCMahJ2n1UQVtnYvrC
GZS6+b+l7QAzjyR7r6LS5wSYsRfBwDN8gYIt1UtFd2UXRDTKgiRbgloC4Bn9LORQ
D4/LPITiNtG5EHckj+N2QIhciYy4Bxd/JlpyrmSkEchphhldiR6BQTqZBQWCS5P9
PJrtqw08utv4R6eBdQkwFl2hk4glx3h10mDLM5SpeWMT14tSpa/fIzNEeWcR8Ei3
I1voP5NceIQ8eA+XumdTO7RxrrIDHYHfN2ne5EeXMQBjicLAdNb2VLS+aXML65ez
tqlt6F8Z6DPFaNO4ZZKEDPZi1ArlQVZJt92vZ88lbo/JFz76CIfVQ8vWj3ugHExV
gEsKlppsH81aIT8RDoVl5O8mVrMyoQjPulYt2xLuYrGYpnNMSHJY06KvSyDe2xlJ
jS8fjBdhLgOd9MkmKNwarGATb+pHL8xdT5ZG2+SIZ4npHr4JmQNLRDb6DDW7m2T6
MO+B7ZQnzk++LanK/HbCLgHVvr+ODVF/bBu/EUMGq2uLasAAajk0pJ3jP4vFjTkl
0mJ2wc0HG2C3QRoEcrELGfkCVTr+TJGpRGXmmkVxrXCfCC3K9L9/21HYqJQKNz1H
xE9pK3cOjiO5Wp8hRTdWJtoiTwzbwn6eL8FXi0kEzazLH8MwBo8HOEK+0wRgE2Ia
exqi5DFlTLQyL3fe7xQSZq39SJc+8vJNBu2PI7jSoZBQK8J7Pm78LxEOWkJoLQT4
M4sUFJPZMU/Hy/mjomjVGiO0peCgYh2f+hgEVCPKNu1AwhmtTXaOXogv6ECAQVuF
l/Fya2lGkbc7iT7qA4E0wtnuhe6rXEvmwt/tTjq0HSiOx7BYpbjyW5r09MBT9btz
wPxitbotNvnZRjCKVd/v4oSgoN4l4A/BvIA0SWiZeZuV0NjsEOYDdd6ntGu+JHqr
hNKiZPTHq2v/fm5UaM08JjQe8bPu+PTN+wkKThNSh12hxVrWlDovUX7iYWR7ts3/
jq9mapyhIlmJ0BjGcnzWerubrjpPPK+CzNim6Qt0XjVuhVXDH2O2cB96+EMS3WtL
dkovWu4/SyybB2E+eR8p00ofxgJaTfbeC1ellXngp/pBYmuzBxJdq3CceYF6CRr0
lCuJcrlm7jnzsN0bi8VL5O1mf2kQFARbyZoW+To4sBy0ZVTMHfTsaePufW4HrMMe
0ctz4lugI3q9iaRU5zF8qx21+T+XmRqk9qQ8DBA0C45N3THyJCTWNHV95mMtHZhY
rfnhnHKO5cs83/q55xEfLI79UneYtLN4Wed+jCbZhfXD6GCUTPWy/Bf5OOqsnte0
GwczioKzl1ehzpSMbfyPk801/NJOQ/kAWbgT/5ky4UwrvnvV6Onj2Aqv9Ya02HR3
Gy3jxOgCkx+uuMvTXjPZY/sCWRSNuWYXfnJ46CbI/iAA907Exv2GB9kSypwG42t6
7TfAXstVaEwNEq3HTdT7CjvsFFdlZIsHpp5yoeNjXcH0YGyRp9+LKbO6womWHfHs
sQUAJcOJvOLrEy82z+Z7+gcBE0XJ750hND4UVoRmFyvpm99JkTuJzE+rDjaIvqn5
rSQ4C4Xe17otsxotsu+3QPtTv1AqKNDL9leBCbLWaqjXf7/DCN/VF7kHtrL72jpf
zMzsQk9YG0WuGcW7Ph3/KT6fgItADDegoW1Yn1ZajiCZyickYn95j1IJxrOC0GPh
rDywkP3K8krB+OHVVO/Ye7ZJ+y9jOLraCbna8NLmW6NeMIZN+EoIU7KoXpdSy3MI
Qt+WYI/4+jI5K+qjIKqHmVXJgGZyx6n+IpiXkM4ZOee6VI1EXiE3TibkRyuTjnxh
+6Ckfmw1RQLDE1YHBStOEXKAWPZMzu9cdlgDM91WJDS1V/gjOWkzoe5Io1deic5X
y58rggdMLx5K7tLcxnWiet/lMEWE5pOaf1/PpyCjvmOJWB4491eTmA3hDfoMskUg
OFtTjDJMJd2agugcJRhS1pMLB4DCfmtyZrcAY8xczWyYb0JRs1Bg1qsJvZHFgedO
jUf3FdLRKlNQI5VHrEVzWSLXqc6kfAE1/EfBLI2cfBzGtJxT7lg2YzXeJczNWMzZ
IUp1ysKlFy9if6V/ws3HwI+RD0tsO7GDbthUJw5ZAkJieckQpBAO10f/sbCmvZ+4
c/xg6nekqr+5uaWgIrE/LFez3kSnH/PlpzY8xzaIv7VMfaaP756lCpoFu3DiDoLG
ZKtx68RTri+btmmsupOVHISpxdFPm/GCkR2rAR3j6BoshCp5bHPko2uzYW4okHA6
HtI1oM9/srLYCFWedmkbmNDxAD4t+U1zUc5r9w8TktVMkwKcnzDJhizPIf5MN6nC
QqYgkPV/MV6sMO5pH5+9bdsnrE72C2uozVFC3JDl6gO9mEjoL3W8ZTCIiaiCVqDC
onyQp6r5ValZ3cGObhxa9rzGtyytw7L5JMfARgKxuSpzYVkEb+aBg1f0+3mZVc5n
wEPYsBGHs63GOzoHKnOEa3j/eRWOCdM1u2xt4zFk4zlaniik2aTmIrGdYU2gfiWf
1JR+EQVlDrhAuUmeFJlJsdWkHMm52W7rE5a2JShueaXVu1HDRh/Gcmfl+5jJ+K7o
cJ29+h1+yHdntSdf0dVIoZnPxC/yiux/sX+EJenDWl68VfHTBnH9i1WjKdACztyh
a8gi2IeCvpoVoYbu0cdwNoIaUVfN3gakPKAQ1UO52wiQFbDurzMO8Xd7F9yZJ8Gn
NivcWMcJC/vT6HFZeQZNO8vVZh/Z0tqPlTk9fhKMwO2Z+Z+ctW8SbhNJzAQOv7XA
h2I2LLTf7bei9o/Fa2kDDhS3wqLUOjK1StfcpXUdneCBf6cvYSd4qCDKYzmgy6TY
SkXS7Mz5ZoLZ4RU5kQA8tbJVB6o6ojXRKKVLWKLqc0nlMZWr6/afFQisexyz1Sbw
LKBGJTFgQ7dQBekjCZwdJphajDt1KXSGN9LQeXP9YDPvCcBYTIPwf+rE7yyMWbk0
hiq8c2LrXx0Nr1VXgUOJiRGy2EohnVtI1UTpoJZf3tThWAvsQlkYQQ/ROKiFgrr2
FNKKobi1EcHuDwofZobFbKOB6abNCMg9kpNHM36v2Hy+kzkvRg3OdoSoQuwUX/yn
U4K0R6YNk9j3Gzk5M8stra62x4q/3a7XKlb1TKZua13hHEK651DCd4rxzy4Ir9h9
KbFbjFbMtLeNT4VIjbCsK3pZawS77lkpeTz/n6Uz8uKDJ1KXr40Nac+69SoctJ2s
QSfb7PsdedgxvZZhc9VB4lgdCwFvIx3OcX3Q6N1XhWEAh/Uxl9OpMNY1LG4J6mux
8vlRdZS4WpTk0rkoyQVAMjBxeL1tXOI6IDi3T3nhFkr8s5ZaIPMMwANzpVWb2kyS
ep2rFOtmYRtXo8oM9tduB/G2W22NWdbiMjNjeIZR/wDiZfAoF5eQ1eGZ3qpLsnul
WR29vCiR1WcA7QGnYxa9hD5aWJYO8eCkT3j/nGA8rkyKcJqiFC848JUdL5R+xah6
yY1qDzGkw+nWxkLQaxPd0zhQ+gp6dr3NZMedT1+QkHpRZq2j1qnVMgMMckRtSJfF
EN69mQSmu1D+xsksCP6PoR7Lzn41JXq8ZPytf1k2SedlHWI2tugfkfdYb6QmFuNL
4K5IZG1yWT7BujbKsuKXnjauSPmflZtLZHlDSxJQ33YWtN+ai1MiDAhzy7esqqFy
r8Qfq735GDbyvvVvCTvFsdT6CmzpHON1piMdKoHwhvsgvIEO8+6vuKuTj2fI9LAu
i3JlfOnek4E5nOxQXoO4BDrdVQUH/NwmueqlKMLBtXp3SOQiQDCAc8cjBDtS+MHa
Ff3WE4XxHytKl75HJ5Mt4OApaOYEn53q5onuSB6ToskrBZ0Qzcmy+kDKDxIeljp6
AaXjAOgTF+ZEadP/LtC4s6dQskvnJbLw0ZmW0KAgX6U+wp/cGDbauxk91+29g+1i
X5wMN3astD2pEZDGh5ok8vg7IF5OI2o5XfJoqxLmyRW3hLuz5MA7eY54FKG4iWPL
ZdblsGVV+r05edSa4JtctWiDHm/FSTLinoQI9hnNsCzio6RggWdpEKcNqZ3/seca
W7/xlBiHFv+cKfPniY+utjbb4RPSGQb0QfVUk+7lvJiR6TOpwm3mOpBxslXm/OXN
e2dsZ+VF6sE1WaeknE9rdl80NNrQVp3jWhORbrtvRlt1TJvmcj+GzE6NOBl0j8ME
sOkSraT5CfmJyKbYHQRxHODXq62NUKTkaB9npBRKjC1iNarfV8jabodgHVJan2CV
Sy+ok2IFPXlYI18IM/S+2a+MjiEu0lXm5rRZacZjyJ/bDZz2UgJFHftDqIdVVeJF
y6yKta9ZxlecXGsDHa+gozsXk++EW/F+2BAQI0onjVGtbMU/2is/DNZWWKbd6sWx
aKZA2xYWu1lya/8QXElHjikoR+s4jZYeO4fg6aVvDwu88izF1DIeYsyJXnJLBcdk
Z56XHhYicot+5MXp6J5Tfwr4QF2ZZkJiSZFr/A+c2w/UirX5af0jHOfZmCBhberz
yTVXebtxx6EW6lyRKXUXPzPAeUn944kNFlcJ1708Npe83Sz9wmK39ShJFL4eL2Zi
pV7rU/1+6uB8s1oKD1pTxskTULvH6+DiJ+3qhrTGJOJnpL0uXlNZ5BAPMDrFgx7M
Axho5PvDEELjok1yW1xqU/7nXu/I+U6yEWHmO+9dcp0RoLCtCcGWbXqwdPTxEQhN
2kqQgVPRizbkIlFukNrkUsiyHDkxikxfj19/NMgRFkAc+pSMQFtSXaYwIySRRDeO
xYqSdtRTBSa0fTGJ1sd3srxAbxUoHLad65us+JGGToPtk9PtMD6z6HMSG/7V+E0P
`protect end_protected