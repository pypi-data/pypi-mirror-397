`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQMy0Nic0oPYTT1PeBRgvHfGJPhS8cExN321l1A6dBUYa
fg1ulhR+nyDXSfvpLc/Mka2zDQSKm3Jah3SkEQj1ToM1Ps2LxH0whZFDHySGkCST
69TozQfaLYteiGye0t8QY3pA7wLjMBNGE9BrvfDykgilriIJ8yd+HvcJoR/xC1pK
NGWMzhD1FlE+t87SodsY7iGaSfs1gS/6VGUEIcsweEIso77YIsjPSzcUWDhuxKsb
ejGfanN11L086K2cfdibKvRhJ5oQakLKNNPg9h5uxthZkd+NqzwJ1ygAVvFEyUqW
P17NvtJ4XeFxmKGUMVRjtv9d5TDc0YGcQzIGyjY4mn9BLFSYlclvCmzQ9YNsHSH9
vRpIh4rKzDXW2RStbS229eKvCDNizC6bCa9Gepm+8bmsem/z2o89GhJ7ip2CCoa5
qnU9TyKKzSYLtCPXwNl8dTlZdQshIjmFViZQn/+0qE3Zu/XRBvqWA2d5xhSNE0Sv
eNKIQt1XUkdORF6KJZ7p5ioe7u0lyxdnyprco+XuEu3epliEczw2nvgVHaFmEOgF
RaFDaFhmVrq6+d4EYMG9/Uuh2ocdCw/jVl5DpHKEDv+rH0GplSgDhYR9+SyOjrOa
f5h6g6e+ZltOdJqjdU7oPMbSVnSu4FJEqnkzQ8CtGxquHRz67qr8Xr5fgW/gdEha
gtX5TnAfu53HAv9RiTGQsYexpNxvtov5btgBkywibSNh4+vAzP/lNIPFNJ/3RMSk
LABMOK8tSV+h7DhM2oab4XSVTV2DoJw47YwU1EAKgV4gHgTAOPd/CW4cM+80NUJx
G/zfQ4kb1AzY12iUVpABAgEJV4bFClWOG4ZdSsksVS9fw0b42gLl5a/ZynEBlzZa
Z6CiboQWZ0kl97OnmdeFPPm0/LJ0//Rq1bdrekB18FDLBzTn76JggpApGpAASh+j
OreisoJKqYyG94JEakxyfMp1ijz15RD/NgealulQglUNHUxIdlRKHZ9kPpK8HCYi
tbUq27CcfRQVzKgB/OOmT5L8sPm9OW1/FCOicPf7eZvwdlcDB9ybct+KFKpW4JzT
T+YKVGnCXGm+YYYurgFuB98HV/e3z1YSKlZ6tEf//Yjua4X5sXyQv9pun+WMJ3s9
4oqLDKuGAbOPkWjicKENX6CPJqHWb8LLSI2BKdxQNnRAVeJ/tWWu8JhHIXnM5/XL
miUKEkl8hD+DAagK0LKQVF6gf5Fu5MM2tmts7+hmsGrxUv7mpBU/okMDi7Qbhe8Q
o7qDEeuZOc45Ezs4gXH8sAHj78fXGOWGsjEQuYzEtfaCoCuTx8UMVujBN1DHGyyN
fRaHCbyEgF6y5N+gFin3Pek3D3db8ZMaVzwXJZ+dKiWzeWlmqsp1i5W0pLh84F0C
UL6Qmregqq5SZJrKOpsqcFyEn2mVVAM2ahrn5ZGWVLzFPd5ecJi3H8b24C3lckwJ
gtpKEZBmtX7ZDK4b3YWBGo+/USUDWEoKHet/wgfFqjrW1ZtMQt6WqK8zO9UQ3cBv
D3lMbTauF7zOnymFw+8sdaq4AGhw1AqFJMtDF9w+BV/78072h/ykqWezqq6YZbY3
2k5WTONPqMRnz3n4suvubZBR6DzAxSI1/OSDAVJ+VlQAPJAQFnQdilQwfcvMS1HV
bGAvhOntRWqG2w+/dhuHi1JUZXEBLG63dDoBMWGAHIJVONHBaWiLw2vYZMzjMIuu
+877LHKK/Lovw+4QMGXukyghQXsbsZxmmYBVT5NznCoGjZ8KuiNRaq0mxbLxPX1N
tado4hjcKiOG3Y/sfI1KMXv3upfehbbgTm0xiAn6G3GwfK33zGY4hKohP2/r3/7G
Ra6QHpmWPP5N45o0gTdhnWq3AbB+p8PFMTkwkrnki01keThGL2lzoOXjPEfopmig
/wC4FktRxyfgGJJbbFOkNdTCoJnIRKs7eB7nj1KfG6GX7SVGPndFb8rvSXnPWCv+
bWjK2Pi6TK3FfuMJnzd7cn/2b8ZVDiF+VjohiTYKBfZpASAkvEhhn3YLJHdTXsnX
mxXxn/4R5PtrW+Gf9965fXnF5TuApjlKSiwQdwNLGSN55HHBVjcxb3pPgP1uabK/
v603hF+o6cPA6+VPSHF8DmK6mAaLyYz00bRrvOt7bnhg5FMnhua6cK6v5g9Wy+S7
FbVp+csJZrDsbMxwZMJLfawNAIGzl5jHLhIL78nzvpVrXJx5o80NsdVcVRt5aPy7
SiBmtT1JpCKKAYt5KM6Y588MSPl2XOYESEba3ZtHCOM4KvOnqCHPcmoy9Wf1D66W
o371zO092MyRZ7k33NtCEUhnuiPqKweNxyEjzo1/N4B8wnGkW1skJ2npZrI4ObcL
66G06oYjb3O3phHFA0e9HMDRI+3PuWygQ14bDt3SyGUExy8kaN6z2TgRwELsDxkf
OySXjNmmsPJvSdQp9pyjJ2cAktxbiPZ2SXQ7d+JwY5qpJXilqQUUFRT8vx2w3NnW
RLAuy/x7tpoy0e+i3tHJ/1816oFY+5BvUSFZDJsJNNYo1LlXJOvBwXjmj9drRzoy
OI/9KTvCB5lRiuKAThGgUivO2QKyZ0UpXVixpOFZXWSQ6fUlEdKrY+Nexr24BoAE
5jWkyncgdmYutlGLkNzTQsYN9EtoQoELiwm+cmgPCV5qWvMh5YQn6qJg+fKaAJL7
EDP0Vmq/pD3OwU4XLZKQJpXPmpV61BofUMbArozBii6ygTar0qB2/VUZnp7fASa+
xeHKxQgmBKxzW9mul0+Gb/3u5R0kDv3+NBmslMpiDttTrqJl4isbU16KtaFBFOQr
39qUNlZLo66Ui5MBrO9Hf1UKhBWDnvx2KgAg/KsvPEtU2gqdpmYC1efbKYzZXv+b
11uh6CH1aYn0KpdHcFw8pbJ+3SAVg5xAi7AuO3JhE21htO0/3fLR5OZ9h4Jjy+dS
iBKkS9EF6+ha08SVTRTReyPOGaJ3KNicOf/xQoq9w3yKVPf5tjCXJWWSuWP698V+
B9N/D7j5dxqSaDt8aAZlItOrKVrdMDV5jXTeQXlXCyoWZGmAUFB4symIVu4Arh1t
cXAnFKEmh++98EoNAJhHFYLVYLzX+DQZBDwYU65Zi+QwIfhV0h78Da9kWVR+OtMq
uRQnBdbE3LhrnmpScomVeoBzIkTrVa4NlWCJvrTYnDZazLWmxW8fdHLZP8NSz9xW
uy6hY3Zcv4xhU7gN60XG+qbEmld5noaBFVOAmx523eQMnZ5C26hfz86q9Aa0YoKx
4v6n1W4+RGOqfikTxb0X3gtdRxpPoGeL7YGK0iBfk3BgzeZouR4gV9ELVhaWOlth
Du110Rr4ZP6WbFLAVze8pNucEq9W848FAK0YuM+LT0fKz+gHBgkhCePRWxXUHBO+
TfhyPwVF0nD/vhEfgOZz1G34NHHRzk+1hFEkZXVvQZKM/veztjtsJHNbiorOo8QT
PlxyVl9svNk0ciHaF4jEP9J6jAHFX8NBDs1ZhPjsDxTS1FmQ4Sw6yx9iwFyCbY66
kyOT9DS1JLOyp9A83ArqfKQozBix58BW/L/JwwIEZ/uhxii5ODasPY3ZdU57kHgT
bspZv+Mm5r8S4KlGJD+IUDJbxHQ38mcLQ/eGW5Pr9IJHd1Ea1axeB24WhZOd2bes
hej0nYq6FQfZXRvl880W1cnFXdxBDdrN/nSm91pnsBkFdK5jWIb7Zoe+fynH586u
EDMsGEoUAN9Rde9a0pncnNWl7844sSoNIJg758N5EreOI+W3pLHQPWYoI0wpsx7E
Z96F7yo8jbxWiQtrpG8Aj1+A5y+AVX5PF/iSKci097NEHFhwTqEWpWPWy5WkJA60
2FhXkCJ9berLiRF1zRq1XE6ceBCCw0H2zQ5IL3NrFghT20Z3iCsBPdUMdj4Xww0d
huhzMfI8GQFDsYVu6oIVgzFVZz682hitQS4LnWNQ0p92TdS8zlPt20jTKrtTpj7h
8h8J6ObXN8GGuXHGEQ/wheQiv5rZr/GsmkDZ4jf5y1L8dsUIFiO/k4geuI0IBDOk
pFpcTRjnNY045tAk9diJVBY0/+u+V/UoO4kW5OjtCs3tCNx0okpK0FUOcMA1rFGQ
nf+4NWYoWo6D+Zwo9QcA359NJIXmvZPSj2hfwlwc6q8V5LCz76ozv8gpDu9xrQ+F
CcYBMW2SF5WvDAfarDrzq3PMQ3C0fysrYvTv5BBWwRX/6Nd9i/k6pqeUWv3nNDi9
bT6R+4E2dWY2UpytWJzRjfb+COFGV7iCLh/fFb0egq4ZuOTEJ0O8A5Xk0UrbjgoR
OzZVy41TqmnbCXy618nVKcMu3oiX6kFIEzwz/uCnw9eXw4H3ZaTavt5s4JXud/Xj
JUpOdDUCWDQC9mYwR2icvyE4nUN35IMsiCspUB/hEX6eQbgWhQLf640ZMR57T7Sc
dS+Z+MKypJ3GQcY6IrGWW6B7rWIj4hFrM/VWQWX39if7FY+8Eq2OJ1KTSJFdzKY5
C0s/dg84GDW5RMcA4PofHuqDKI+t8qX6kk6QVw+cSieDZP8i+mtU+yGy/Le2jIA1
BmAm09ssgtCS/FClx83Yv2N/7N2JFQKuADqhWpGB9By8c7czvh5elMC5fXBtrHkF
EqZqIJmGFA3ZLFI0fdy583axG0e/FByCdyB8uDynEwHagB+OL43IBZUvXGkpG8Ls
eDzhtjaODT0HKs919MXCv5j/znW7MDrEObNxjHUfw0CMu9Y2CW7sAXSZ7Mbn7Frv
7CLZfoqMpQ9YmaO+dI7jOsLzKE2ilA8MocwgmUvYyBVjzFAEnLgKZfXPzAqr87EF
V5SbLIML92DmcVQ2agQArXNogvdY3Syz9VznUsWEAhewgcTCXlVgpTAXDkmGXFWo
QKM8ylKyLUmN1nKG/1dyj8zwMALgf6cELhMn1sNqVAjbChzW63Fv5XUdvmKnyk70
UrqxX8bWc+zNI+eDk+WgyFgcEZWGd0O/QVgZNtRYv4wpJvHGqEtbc/5dggS791Rg
QvGf3aRnUTREYnv4mbXictrIgpjPZllXhcBN2b7r2qc22gkM15FmvazpYuUDcBsj
K5sA2mhhX8A4yKZj1EVREleK07HqQ7DFl5A30VEZPzoITa32MO0mbInMYGLvn8V0
7g5uIgqM2gt1mm1rHbterw7vm+liZu1/Y5ANjI0a1xpSoWNzuUNsZuvRyHqZQbmm
M7jWSFkvCGh02aOR5A+YR85vN8K/XvicxMu1Dk7V2ax0qyhuYlDlGJmMQQuhY2Zx
dwb2j8RuFRE8G5IwXGxlrssm0d7hLThyUUYAlIG/CSCEAUT2IamNLZD+a/Emd8WW
aTJyz4mB0lar7djQq850hU+VvwZ4Y+7LFqrwaO7zHk1K3ZMzBBcprWEQxrxr9+Da
szO/wEOAwATIhH7Mg/hun3cjmjGPYQ6fi9a19Rx1SK7uNbU3zv8k0NjobkzNqOM2
7rssiNRl1Uze42gk5+KIbZ5SiDEq/0WSz4FsZszlwUR5VO6727ILakP69vzEEF7V
3uKQle7sRRojwWUHXan/51YODrBlsk7+ddbteaXkoYBME22+3BZ8DgnB4VWqRR/O
zeb23XVJ68s3uycHzzN5/1v5nNRiwdcWx35Wv6y5+Px4Tx5/QbZP9P6MYxG9vtqZ
OF/+DuUfDtBdBgWsouQA8VoOJenNGBCejSLXKNvsGEGq76l4vu7bGKAUU/mtj8nz
a6nVUzyzErUmQyU1ADx2v/7ddL6LkkOeiMDFQa7MCM4Y+2sCNprkWTzqol0udi8T
4dOGJBh4YSU8c5fppu2ar+gmJIBSDj6xUo33hcsIMVvcURHPF9cg/UDN24YsJ4U7
/mufqtR5qR9GbSzgrcjkI6qKmxgy5ga3V6Y7xkvtLeFzPdYH2wM3Y1c0cJg2UCco
Hs7+8dFW0OZa3TUOSpxtITjgBdGWiCDfYswh1PQo+kITj9/LHlHJTZ2P8uFlo29g
hrdze7w2fNP+W4GEkgKp6PDmhPK1FEmBRi0uOSzpypBAn07hBvVqKnKSxOmIldPm
tQJK8ftbxN7LrB51AqaVqG8lCxhh0Fxh41cQu2hFgFfUg4yJooiqwca0UoQhMgb6
R6n/Ukb5KDs1oV27HdUV2AEFI5RmDZQJpDtVytSjVJFXdVyPrX0Y1M84xwCUyWSi
vTPWhgKy1d9Fq8nPvPon3EvcMC0hIgcBnO9F93OKIvEZNz7CAGV6Vfg0pIAUfjxs
R4a5ytZWduYTWQuIIW0wb4HYPjBGyNs3pbFBswEtfL21lE/wKSVWuw5y5OUkqht0
lKR/4tAODmfCFEMSlr6bYjaaRKMMhty+zbzZjOsCkLaivVLxfW+FAmy7l0oHhPty
MAP+SD97iGmCR5OxSDQST4xfi8RJ0iYArmNIJdzz/3nGDFbqT8yndQLGLZrBDsMv
l3TJ9Kq/xqHP/WS9m79BJ2KHz17TQc/WuFK0gOLP0FLgG7uWmYBsIXb3h8x88Rxt
NIAaJq9oigOt4ktQEhxVHI4ITriZm1N6MIK2URhiwQnAA02sp1MCFn9wbs/Ck5va
0TCCCAoexsXuw45bjJEimHO4t9es4uxOXBXenqHCnK+SsCJLhscBvL5tOldhKXCE
a+KJ0Ne0yTDO0PXlS3gXGJM4yFvF1JdCcrW5QV9cFz7j0wpiIyloShYqtc3nG2tq
F9JP3DxX2yecImWqL1gZk7rSfOcHaBsOn6fRGvVN/F6KO+TNA7KMq0O42bPwnqvR
hLOQ2JQqdDjpKufhQ5qajd8Qvj/4uFrBscNThF/VLmULiOPCxur0/x22fL15Tfxl
GV57Xi735dlhnkNwmy7M6bbTzHFRL0RymZCeKtkLPgINtj8izN9mhDqls7j9TTuC
Ej/1TcKTZy5IR4oMBaQ1KewOr+GmA1a6lqAWNdTCChT1UhCVsWZq3WpZRjq8UjK2
IpT3PPm3njEPv7PSoVjArNt7zv2tYgwR4+qUwlJnpUuP5VSvzXQX4oQPIE4yHeQl
gKxDyZYXqq1TBOL9sKeGcrRDM6q0ALuIc+r5qHag58iZtnseMaWjGnLLmYH5GMyb
GdUzOdi6/rfwQubyMfliab7nwt9mC1IMYlp/rNN4PG7oIR7IGE0Jn2UObZmk6YnG
s90yByGx2kSktzXQuttYLDWCnsOUDnZ1v6vwQv+yyAmEF209lSHA/N65xBUhkMi4
olZasDTMyFLpcdjCyDAMRO8/bBQXQsxT88s+eiapqGsV0usxbZvapFaxHfEWSbVl
JZlpqnlwa2TpxpsSFIDOBjipsdhCglPeW+TCmsQ3fcKqG3TB96Jezm4OD4i2ySQS
I9RNdNSmc6XzYjulJVD8x7IByx7gYTredjJBn7bPUISVlmcSLifJZYf6OtIu+5t2
SRlbRxS7AdtYvc8AT2LmMBldF+Q8Pvh4nPc79XUoShYNkPwOlqrDZ7S0TQLSlNqx
hKcVAobPSYL2jRXdaUul0vQWhMicjvLZCmY9twHiDtUCYkw66ngv87ahfIhv16hc
2vydMzzjgX/iZa3ZXMQXIRiECL0uYunj4UOQ4LG8Ll2TOdlSOzIWbxOwQBJLLZ5U
loRoTOMHF6SSa8e4KzaruIRYWr4bsGNQarjAO8meqjtJBk9WvFFVijtac6ZeE0IV
Jsv12c2mvx/DK+zWAlsIxFoXSTRbsxo2o8s2w7bx/PUu5HAw8faTsgY4VuyWt3xc
zBSNuCmdnJw96d00qiwvjr/uoV5oc5sK0mFoBhg2sCLyQnNysOOE3fc2hxLrkW0i
ZF7vcQGOq7lGhxKemHim6us/jzVKD8s4XDsEOQ4z966OD/6Kg2YcTxBHbUclyga3
y4IzBl/ALg9pxTT4RQziI7b0RJhxx+qWB1U3M3n0NK6u+tbb++7uNfUPRpppdZ7/
+cIrz8Du+pVt/8KTlUXd5sQ7zvlgYJbK5hIoVOFJwYBnw1wFphfV2b+OTRDUcygm
opDg+YNDr9K/toYb9Pjggvo/cgO+oM8fThtfKvc0tkXKacgUARQtBVaoQh1SuzdV
DZiXrSuNRUGE1IoI+mGxjDzD7UHA97Og7IKwwh1D8KFbNLrjV4rZTPmGa+/6DP/d
2aDth3IaALDd2AWRvZNcUsDINAFpHAs0w1AtVd2uAImKky7NEcHiNr2rHziDJd+j
a5P1W+1EjOFeJlqmWIKIIJV5V2Ib82GvLxEv/r/1CyJQelTPokOR+ayGJ3Hmr67R
jmGtUGDYvjS5BPNvfblj3qLjV6WAsKftvOJoGXwibkpdu9HUK4gvGqkiSOnAe7H6
YcsKSpcUH0UNpZ/85MH4EqqL8HbnXBf+/yz5dBycTQPDAYDpwXAmuZuoFCao3p7d
ZEH3VdYcenB79lF9QF4XSVUHxaxV9cWf8SlALI+ZQISBZ8usHuUjRoyfYHHDQL0F
fO5WucNbFbTGP2jCudS425wQS9wjnmBGbbSifZWyiujtJICRhljwe4yy9T90idXP
+2Gy9DzcLDWtNdegqo2fTMCVRUgCmpVlQS7+BAnBHI/B1bYhI7oPv/EdBEJNE+dM
PkAHXLyUKJm9J9P2ndqElJfIWiu2iRaf4FRyiZ3hCxFzGOwJOujNw122l5miTXfQ
Jnd/JnrQjoeRB70aPlK9fDt24+cJ99TxQ1jkBmr0oNxwQns2418P2PdH27jwOPpR
KqJi9pi/8gN/uGrlaSgasBEjaBmO0x3tM02785nyIxqrr9GNzWL0VTMluzDckhbX
tbNd+LsmHhMxxv4UK11ZR1+F8aV9jdNypwOdvdn8lwWGywDUvUJUmvrrHNkVTNRu
7m9VJgAj5YCfLKBB00yeB5hRZuyWMrlpKAc3dCr8wog+ui7MykVByQpFBu94gdxu
x3CwTzc4mKsfUYw1jUzP1rt5C64YTVSt5aPTj7s9VeHSZ5FyYE3DyKRuoxoEIB9l
iyKSNGF38dv8NrfIttQZotI4XkfrXOEUA1A1PQSmPK4SYqd6ghvFMFyMYPVUjcvr
ROcm5IGgdZ5BuYl21fSTCJ+NnLVkgdgtaM6/4DUHUKa5A2xV+VCUh6BodHcwRvkw
L+hJ7XBWdxsvOZ+8epxChIAbM85WCOl4g02525WZjY8RiodTUoXPb/Lrj2DTBqMQ
suM9rz60zlwv3K4QsRkAEx4j+HR0UEWjl9KVQyxvLj+9AvILVGHrkcCNf7JxOenK
EdWtQDC85cZkEa6lPU3WYGPT/p4du1Sq+aYllMLqzECxmc0CxQcZA2CCV3iVR8FR
H0txzV3p/ET8ku3+O7qRnFUjxoXT629fafciY515MKNf4/n1rCFa6kLenp4l01n1
RzIdl6k24BmQkD+QS2720Sc7DgvOHgmI9Xq8lp/ezjZCmvu2H9E7lwFQZYHjU/J0
gImTFN5Mvib09/DyzVdLV42mWKi9dj2+25Sc+PEwUCABwDPSyrqHLPG+uhwRNdwA
hqt3ucEXMFPmI6z6Gy2BibPP/jkIO+8KAUQRbCfkITbPUIykJxixtbmZvJC4tguB
tDdya9/2IbS7RtT+P16t/6jhX6ZJ8GLDXPu3z3B2QLWO6GnMScuzQF3ZyKY4ctG9
dwjw02ISvOHLaGoK/qaERAKpfFz8kZVG4pOgDFYBVW0UISIHlvgUvzUI5ADtNBpg
4j8oF+nJiRYzFBbj0XzlHqKYcZwIZuKirIDpthSYKNByLJLIZjC2mvbFliqVUeE/
r2sNw1/e4y864qs9Os+TmC/rCVS0pHXeZDOkczvIRDTL9FmEUkpFWXpKLvt1vBWK
q6h6VrTcZpM5hIYdV6nOP6weqvyh5PmrFWKTS5VZQnjUtvt46YoS5tqhjsERMe3P
r72320MfT+o8XHL6mEITininCpR8/cuoNDdV/sSztcyetTRUQhn2uEcv4hegrqoF
2WFncTTx+DMKhBF+SPPMN6abGSUe8RikRJEKspAn2ECuohdpv+LXRLoTv7znufB3
1gklY0d649tPJKaVcPezI+qJiyqwjdcD65s4aoEcEkfirhpiJhHSP/ekRVJ8xqJ2
Ygzyaa4aUn5a5om10B7pHGGul6hTraQZP1ZztkuLIonGyNmsnuL5wIbUVjmQBmg4
4iA/xi+/mqOwji4HusgLKOXuW1YRfehKvOklxrtn/EnbK0+G+2tJLFzw8oKGMLhN
jsYRH8WSNMu5ycsn7gjHCZQTQr9SU8NP3Tf4kpQRwZwZpP3ipz20D721xbTpon5p
KigylIzR7vtpskVNBZK+Ixdu4LHyoWx49UEICczFpV9D13CD2LBxJHV5k4Mq9no1
2UsPYNDwJo0bU9JZVzW0dwnxxPCwkJBuD/izaB9sWyA7/GUUjnuxCDM8LaKzdfdl
jC1IikLItiZT/39130GXwqVdVqdwkv0kSgtFGgxMpKFslMycncvij/ro8v2p/510
vDikBeHj4S34dcxBG1O57OWTGyS/ccfBj2ZhGiAuXatCnk1n9bP+dMPWIwBPoQDV
c6wrbh1UBjA8nZkLEQVIkio3AJ6mZ5hO3FzVgN4vn+RX0HOfBa4g5mkHBeApFqDD
T2cNzy4dzLfO2U6xUDOp9TtrHcvYKaU3lwBdAoEZ4IIhvIAHYMMN5SwNRoTSUiJA
auHLmj8kJW6gciRPAj7HYZ3lnI/RzHNX0CgDyCsPbnnNACYprneWNJLEN+nvnCeL
wX3TVXjL9WkGI3dFj+B5VAJ/IMSYhRkbDunfBLmdmbfopoSAHxhCzO13vU6kw/uG
PyfW6hPGYFx8tW47r45y4kWuElAzeXpJxUcrFNTh1T+HhFIeE79tjgEAXfP85RsV
92+UWkiG9DB7lvr1wzs/PIKZ6zqxSW2tNcSW2rdiuowkPlmAaTmZ0naARItmIh7O
x/HPOTwcCNXptFAOzf4e0DjTrpfpA8fDlRtn1l/fv32xt+ewzkqO7wY0G1zbLAf4
741mUf72tKFT+vCYHDOQHRCGWzc22mYwwmnKiVUWVCdZzRzLVCing4I4biYieg/J
GJUr49+zEcgV+KDm7F3A8oJ2OtwD67YNgQxQh81nBSwxEbhxFuhK/iNN24fT4nIP
JV2tNuCyQqfnYaF9dVCD6NczoEZC9EBYXxeptZKY6Z08lgQfIoRLyR4BK7BxV5GA
82mJ37np7UzZyc6ikoPDriNOdx/cwSNyimCRmU3iWqo=
`protect end_protected