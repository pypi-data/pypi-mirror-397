`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
Hm0rc5KfjNwPmEU/4qyz3a24v0RsApmt9Lh8xZtRWaoplTDANXLXMeiO7lc+sVMT
NVgoNAdWa19bgg6pdGxB93/sUU9Zq8SadqSTVOOo11zxmcbGzdtG4V1nJmupMnlZ
kyu4+BQBITz/vkqTXrx1tjbDyTbvq4JrMpwpovokOI5yjkd2fp6mv64DzZ+HIppa
sAu/5dly8w4K57QMWB11AcnYQPTWYeQNbw2RLaEPLgUMa9bPbkyfmITJ9f6p/xvM
1ZG0KQzAJQGj2tIgge4U+JinkPsctGl3waJPNdkKN73OEHKvxVJ/6DI11uBiJH9G
y6fHJUfDuknE5HP+ev7hjeVEyLWpJRYOH3RDgl5sJoX5NaB2zWAh7h7Z/nyUiVcl
n6clMUomMgn/ogyMp3uYEA0/fz3Otk+izsBrGDE5z4XWoBDjEwHWJXhV3qVffT4K
oiarl0F4Nt9XHAw+esl9yo6DOjkNu0NhBYoiDbJvzzSyjTmo/VYDY0afGu0VUKZG
eqj0d0tzvITZGXGlbDC8Li36V8AnIVzN3iZ2JPRWTF44g7MxZebvOditczr6VAh2
dlrgHen8CWyzEicMILbJHnw7Qn2g44W4s/+s9gQy1Qpf611drsVHPbKv0nvf5hrP
gm84Q26mTXAOy4tTZpDaejty3uTKcSOMiQLbIiz+P7HB57usVoNqy4o/p5QwrbP5
Jj4rzHUwMOAeSSxMoCJ6UWxriERWthfHFeXBYzuwbf/GFnR8arxMr2UyWNpDkyY3
+gzAVFKcteoYnVyoDKjGDCntXWMXSFOl890/jgdCG/6vULC5CDypf3Awx6jOVUKA
fDEKZTf8OczwUKOacwduu9ISuEeuDgJ53zhHeIEE9b/6F0z9WW8DTXsYBaCmA1v/
d2Z49n+e5G8E3DM8xPBSRyn3Iu2ywnFnTSt5yhcszrfUJ7geLdNc7uI2gYVlkgjQ
kjX4tJ8YOc+0d809poTf3dk0QOC0m1lBhnUmxulpyM7tm71AIvjISYYVQg7dMWt9
DEJZApY8s3q7FaEBSv6TYVRgmCA+kACdr8Pm1ztqQ/XBSP3fKhTlDDVXqs+XGF1a
qziAAvCyivdVYI7Nll2I4bENIpf1alGnwGWXGUF5gUM/GXY+Fbg+S6i3k+amcn6o
hRy2HrwUVcNUUpPpEKE0B9w7X4T2W43GY99pt35r5jsofCfyFYHcWWCIqJo06toU
MplaF3AnsVwLQi8yeWfFyvfutghpwnu0ScEBB3x6cSErAZswp59mO7816crjcjMT
T3NieeRvnUECwdMrRQ7v0bbciWsKhTjVAEtZ/MrObNT1Pxsp1hk/RmzuWndgaz1w
RU5Wvp/rdpFRT/5QLiHHiKXe2MjW6UZKqdvYhn3BrbFlcgY6AYXO3NYmKo9xxs5/
2/U1Jwk7BZTAtgZltrFF8qpytJyGtdqsPgrHCJg39SUceAaGcyPP0HGfV3hC+63+
yHbjclTY8Lum036nYptQjrRojumj79qqU3ubi95Eyx5q5pmyZZ2nTnkCUYsRjb7u
hwUWHEIdcnFScHq+NmmM+Q/j/ROYJabfFhI/VMMXEcgHAadejTDnu5Jx0VEjiVJ6
K6MIUn+obtH0FKnH946pu4Zfqa4zdRpG97ZLWWvUD2YutB48vucFQg3NaW6POxUI
XFykfQptUI2zmZUv/IFpgtsw+IOkdXuN9QoGT+h583WW98I6F/4TQdEjJotvUVFC
0UhHDef9Eo0FZtJKnWLiPA7NxOKE2WtVGtMiRdi1pj6gt7xaqDs6Cfiir6Bc4Q11
IZ8nU9fNjYDRDZPiFNAKnz1OGjNAec3A2Y7KxR/Duy3dUfeHkM9Bl5JBoVJMHqD6
Yt1TN9eqQdRPXuO8pGvPi15zXdQw1I6oMMqN38/d6rim0s8ae0DZP/OjK26DSEdt
ekaAbnudHq1bNowTKlSthZ/xiVSi+REyRf7o0tJNtsU8gduc2aZk+yuct4tBVzx6
soeqyEOtvdx5Pa/bcr2kUDp2aMvAj1Ai36D+imdREONbBqA8ZYE7gNNxwdZEDG3i
LpcwW8BucUc6A/CLLi0JCP8iJ76adUITMwBEpC4Sx/nUzwjM4gzDm9XW9M119JGf
5izmditpklqSWhvwcBnDyCsK44mHsywpk21SZDQE8+BIKAboV97YQyDZ81xboeL2
iYzxXptii/0zTnE07hpIexlwUpBwb94IGD7u/WELbbHdqDX2W2WkkQBxTlVVxSDI
N2KX0kLEQFnWdvuEqqIVfiCHx/B5kDPhF78Qcw6dEtASe97DUrKtquHYV+u8RTtA
VX0BWM8vskSu9cEQRRCOYxgvLTNbJOEtNZtH/qRN7E8QnbD9w9rlgw9wSkaOLMDa
Bp3wih2ZmKfjwKxR6SygewnX2/5ZNlAdM8gy2F1nD7HjprbhD/ZKFgL5esn1h5M5
sOMHv92Q+FBI/SrGS+ssUFm4NnqAw6CFO4QkCmb+2RI/gYL6hBco23oCpON/i14y
7mEeHX5qaJ4Vs7EzejkgOv8xjZ+00o2P6AXC01DMfOYgebDjYlPaT6cYWCz+d1T3
DHYaKXbQnxqe5xYTgM75cRr1ou8DTCdMGGcV9UAQBdF44yqZ6p55m6WSP/do7KEW
ud4wuH7wDKiiHLbe+Uoj9EAu4KZgBvOE3RW+itRoWM9MEcjGezFvt2QBj+YCtmFe
4vbg0cgqbP/ooj1PMjuEDaXA0YXxXx3wzWwnq6w9m43vZU19LkZJZpEVPBc3pTBF
1jQz1nr5jeke8hhcb8YHv839+ZzAD2e3q8IKIRY3zs2za0AbiLu5E/4Bwv9t/N3E
FiixDrekzB4+adQG57xCxFeXKry9z4e3S5pNRCUxgQLwVoXYk+sdsWn9VNHXG2Af
4RikptHaLtuubfl/MParUigejuw3Wo8979Qp6W2xM98IGSsb5ClbQS8k6XySvwIw
RlZ+m8h4BPv/zRy5+VZ7eLTtcIKBWtCGNltSx/2VFmfTKu9DEk526eFre36pnYEu
QPyA8atk1wkpdJ8jyTxecYmHN+Sw+JnvagbMJi4Py/HvEG9+wFIlUsJzkaMbREXi
LLZFlZyv8fz14NYuWzvU+BhrhgROlzhkRd4WLLi+FPG4MVXehximV5Y7WP1wiYyf
qxzkQchxmKYaz/YiyXwoLMxy0EsmKa2PTAUIsobyevhfZgm6JpnMl8bZKYGfjyvy
jx1Msp3zekJ1tCQaMGzvTbltLPOCTU++U6ocwWCGoid4gM5QNyrOtQD7jcom1uLY
bTYF90pWLDgC8KwQOhvbLugJxK+/XEVrt7ZCZssbo+lM4rtoeSku3h/HcDxBzK+s
2AFWJkFqtz1C77ZEeXQwrdawr/3Uw1Di/gtFlehGVLikhIIKWTTxKVEZSsh7YpR6
ruWU7y0k4IW0EzZo5B4HPR7+tyBPvZXjS+JFIoxVLQdnYbZiWnU7hkDUoKRLPclg
GUHhhNehLSRLio4NSLT/OFl/VvQrNpd056SucTamzEpgJrmGr159wMOnQdeXug1x
QTsKw7R18LdqCx6liG1cZgyX7ayQ1qR4M7XaDgi7BveVoFB00RIt3rrfVHzzb5QG
8T9AkQBk618JSwmn/cpXtMbJbn0Ku2/tFu/DdhjGzocK9ch7W1K2WQ5yoequNKAi
uR2Y7QMWk/tzHnPMlyDnRpN7dECnnlphqA860gnoN//cvH1ThLyRRZnCjgyKRzra
5r8z4UpmhLJLMwdGOWoH34z8oxLVM3GgZcNfFMe2f9LDfMZZmEl+ZWB/kvy7Ti5S
ShxEONjhEh+7msf85jXFwD3iqq0gcIgrKSw9Rzdu7gZcpB8hACGyo5uNpV1x3EdM
tzWMZchMZ47oJ1HwGKsTu2LTjLScuJzh5e+5SJSAg+opuMaPd1Ec233YrnM0OYwt
DIOv9XqpvU4DnA3Qs956Ip51wuMp/WtJx57iKO/CfrrLX+7GRft0O0S08RPyCpEB
7PXi7ZMK7gnywhNgbhfRrGxGEx6TF60LNdgYjUC+fyN3ynZoTJtVbfmsblQ1TgqO
cDK3yiubHf+FpWUiBhG8YGDh39Kztb9QxO1SU5ZVA0Xq/brT525myPqm5KZWJknt
M4RUJAaPteiP1CFjPo3Ur02YIkxXwQm9hqLi9abGGCTDEnwdXooCht5cte3wGlRn
l2eqRsNkkYtRMPlccAD7uUDaq/xgD2fUXePb/hMOAQUkdFyCMLt7uaQJxWiEBmo6
+n2lJLy8XR9qkEfwUVdrzxYm5N8ybD1bDq8EXepZXcLH2T3+veDe5zTWC39BayRF
5jCnoou96aSz61jFDRsLJ4xJETIzB1fSSEXPCjhVh9/vhD8Eb7VZMDTT8Jh58QGJ
Q92kf3YgVlzYFQznB4cBCV6pdPeFPNbNprRJqNv7lt8VWdrFmStUBzPbcV/5fKIn
0otlM4qh+yG1RyeBS5pnUDbWUcNUZM8J5CF/QRd6JfsJ8z9ua9zy2HOeD4WEw4rw
Tbt5jnPajvAnsVTsd+DCL5wsxaZONrvTYg+bw5FUZRYzSRQMXhcjPfoDIJVa0sLI
4YOIFmm9ZxUSN7MPMzKGoqkyt14BZj3yW9dhKIwOJ65HkBg2jsEenuUmcAYWGT18
rIlqtZHsCj+TRF4gw6GVQxjE6iDTowrktARuovvcY9sY6dos76z5dwkSqAYNkTj4
G6Oj8YS26/mhWs3OixMqtRI7Mm8z21+SBgidcFjiypoKrnIbjLx+3PYX7Qct6S+d
9q009VJvxa1vAcs1FyHIzLLEmJJzz9gjr8KJIxpOxce9fbOXlmEk1fIsQ9MMBCm8
DSBtMycYMGmlbWreg7919w3w6ZhVevXpg4GUWUdf1e1Fe9sG6IHo8uuUb2nwz80k
nrAD1mMyUjyxqgDpoaQtvfuG455a8wtzW5eImFZ+rbYk0w9ELDqNneHmsPA8QIBb
8OmsMgtp1IRFLOc3KMWefdydGmnEXg0pbmLPgNcELfnw+sTUq11W8+IhEIpM2iOR
gYGmL+nDwX9LnKsKecONRqppEmb+daO4E5hjzs/x3O8+pRLWssnNyuhmvtPSdsvG
w2JUU+DyLJquWHEH5sCUeURz/h0PqGc0bkHE+Oxu3rbMs2dWwz8jTEawBu0+kv1D
WcRzDvvxu4pooyRDVlib2Z0iTz0vlAyfLxuEdSj3TGzW3CKS/erP+SoUTE6JrTaC
chm83FnYLeP+NDR7GQ2aF8C47Vv65T4jcqq2Rsupx7bgSI/kFRkOPJX4KNbcXZj9
VyPjbI32M6QFDi2PL3QXQ8RJZRVwotmcdjV6hgxeCFZq7ebHDTFp42qNOxFI7kCX
dwlWVIPdBsrtHkxzjLWtbeJRkURuc5MgTrEsNmiKsPFWR1PaEMFTj//l1QKEYufX
7lfjGRd+4logYNj/K0QRVG1gRvEb5XuGEIxMtDy3sYAH4qaoODPIvJy9WSx109NR
nnEsie5ZUTkax7lSnzgBnOFbGP4+wIa0dFu/35LFN+4n2TnV1AZAdnl60Jj0GWOl
uveKR0tVGz7iGYSmS9p5kpifnYeCVzW8zYZ7K1GuiKS4hUcMOYHzEh301Gc+DRNT
8IO8stCAd0ZqSrnMAnvKNtgSrQzKfgqsx2/H1i2m+29Rwdbe3Ir5iTWfEIpodp0a
QGwJ/dlAj9mODrhyp/pjksOBR9nLSk7QLlhh+rC/yoglHLaJtl2wjmE5JsnkY5AW
ZHXHydTiJ4aYj0EKcpDWyegU6ivoeNNemEwJYBtdpaSmWy0kGMZ5zkEDWI98xDYx
OvOmzUWxQUBw2oJW7JMDOKXaWbaqGN2f3XI3NkMzIvJ1/7u2KWF/VMDvRHsSBnj1
lRUCN6AhqyzJAjpJmxmk7NI1M72dX8H4cPUfp9ZiswZZZqxv2BcESHVUWAgKFSsL
DPLf7ixUiDnhH/Z5CZsHf6/xwyC9r0zQlWitwor2/mA5clSLn4mo1GC3gHaTo+IJ
KZllA1CEgRKRa43qyiclO7MyjPYg/ZMym9jzyWRSO1yzjoDMQFQYXKn3BRem0RQO
RXGe06d6AmCE/Q9eqLGfmBJB4RLPjBh59QTfnBhx3v6QqoSkE20Lv/dwjvxSlHSt
F/WICKDZVOIPSsUdO8b8p5PFKBqCNFqA5pkceoLcHCkOdxSXaiQqDYfBFP2QsKWa
mRc5flBAiUzofauSTA6zWqWCsF6xJVpzwdPhwcAjTb5idUzxcgATT2A7PXi4QirW
0RZ94YCMZccVUvIZ6AJzVio0ZGZD4qjy4LCy89Ln3NenKuP9IO3xQPpgMPgtkKR5
Lg3v6i8BXnEPPHeHF8ODZkB0VuEP4jbDbI61dA/wBoUExhhyNFaLuIJIKOU1ECDl
1y/jBr8iC7/uXZeK9iF2XlWH9Rk9PLcV5VK2smfQidEm0MWfMnOONy9bDkRO3N6h
8SKHJxBhfxM9EpM79dLy+DIFcWo/p7t8hO2VJ/h3jMPmS+AmeVAPI1Z9kQEMU5b7
pYe9VRPAwL7tCIPBUmKjhqp8CBpDfnFCfJHEPu8rSrenxK1wAu97NUkOlsZARDUB
xZO97sYj4wAZee1z0eJkCAdQxbPcj+LIyaiC4QrN6DGY1SeTqDRognn62/2orW3t
KmtvOg1GfojE/3fEvDdDKBj57l4NS5JvGpzPbl9s0jctaRv1njbPIsHQzBexMKmH
Ma25R+19/+qAB3ezykH+4H8mWtKSfFnjMqnzdgvSJd8N6E8U3VJAUqL1okGmk1y0
+Gqkmuu/l6X2/0TqKxf1EXMRuCNFsE3qCnkiCMfoi4ACYN1KGQB1uegC/i5R0dXs
ONGMbKaJLQvjk3jUapNuIzYubeWC2x4MXs3d73RYSbqtQd8FkMSkKGyN+c4IB7w3
SN7hgpCCFIajtf9gwUMhilASto9Rfed8gNBgK+MgKkRGc61tPllOl2lGGRCuzR6E
poGF7TKHM4N0Z7iyf19wDiv+MhZ8Bv+Fo0yCZaADfriPgBlwWQE+YWcqfwcyiy+0
DO/ETC5kvXt/FKM4tNKzL8uWu1ErRJoAZvAp8LV4tPY8vOfitmeZKXdazCXAuNq8
eCiFRunaTHhRFzL53iYk+TW2fHs6kuGEXJ6w/37hYgfB46sdd4tr1JYlpVkEt1k9
Qsyl1g3VoMr/I8UNB/Eobq9ec1DSyov9wRDR7KBqzANyRr1PKmaCtF5FxVyw9wOI
aamAKJnR1XJXX06hq1SAZOXLyvEibZk//2ae1nrS8j6BZVp7jvZP6DvAe6+YKQWs
sX9AZZnOI2pqFl4vaC8eVFeDNdYJHIFeuIH7rDW+wCygmjp6KqMzwivDNkgQK7Nv
vgT6KopWiMNC45L39oh/XsAgT6X5JYJ+S0Yxert3PNPDQFIkWOhRwRbpfpD7N3QH
YReUg+sHgOE+ReYloFdilzB7eOf5gbzi4cra2/LCXXITnQ5QpkKGwigiGl94/tRx
T772/9P0F97rhXvwP6bW6TCz5/4L6Tx6D9ljH66Y6Ht4CC9vafzM5uQOQuYByJok
6BrEutfcV952T34f8IfSh9LFeY/4eWHJ/JcjxMQYIge8YHFRRgilw+qoVdVns10A
o6d3YvTg9xfLAXwcSoWMap70MyMOFdKprmYq+hicCp/3Bn6Q1WUE1vL7KSmOqDhV
ngD4msXZXSSapcJAlRtKWf9dLvJiwu8BCsF9Ga73KhwfZZHfEg0af3DkUtxmksb4
lzCYk/gLxsGNUsk6jk097hSXsz7HfFtLS0EPqtc+gKdxyJDg9gjy72xOAhuCS1FU
1v/EIN+oW6QDY1p47x4Gi2HPl/hVL2wVu2S/1b49U/MwbUoDRYL8mxivMf15S3ry
wQvfeE1PSvsXaTXGnolfMc4WXWsuxH4NegbuMI1TXmhjADTH8ZmRF30yMZtXyFHl
RhKmZS+I0yOxbG4wC9O5lCHaGLoVA5x/4bVTTXg0mwZsLnX4+oVSG3Aavme7jx1S
g/+fVTmi0nm/VU4ci67elJ8Saiup/wEpYkPZQ7pOzfq+E/I1Kx6qeyvyM9EpJNev
A0BPfWXPqi+Brg78D75/Ld5GEzp5RAd85AvaAIEr7ooW4fm6gJQ4EHYpvMW3r92W
POhEc0nQJ1eqeNupu6TRFWh7P1mJf3VdsPGYCAvRcFq2Fhk90Yow90ICOsIj2piN
GGLPPOjszm9W9mfHIEwKl1qh5NqUG7rEtQl4JGGj3vLqZzAPI7mbiP/cQEOf0uzA
3KUg3MUgNi7MzZoTi3peJl0e7exQgpm0EIOrc0A2juYx5Dz7CZEj+UTnMUJVd7x6
RbPsGlhJ3/7/nPWoe4+qES2BXnv1LTUx4S/9k9APWtUvJN4sikLwVi+gNzOQtmZA
XEdMtE3qLiGPEGMML7WURHeFs8buTT2WUvu35CmKoRmW5C8PfYAxCEwGRFjoITsg
a7LHkiEPHmfuwJsWAVwVeAEokCLcjFwTqWrooWQ3Wrq/ZljfPtC937WLuUwf26qJ
X8wftPxGE66Y8DlslZL5JKyoSmHaN8f7OULpDg1GLACUEffBp0mpCxFdlIPDgGxN
BvOjrf89+CyvMOUuG/wrfQOl9pClrpsdCOlLZiS6KNfHi9zP5KB6AxPKQRIv5ksU
A9J9X+xecgN7nHjfmUAZnJ0Wu24Fij6nXtIvEqswOZ2ZFC6AHoh1hSA+kkAtJurY
YZP7iu55RpH4bJriAVx83SUNNBVFgK8TDJ5t/ZPdHMwPuz7n1pcS/2hy7OdFwXqI
Hn28gprYTCbUec4ZuGf1c2kmQLdxua0c58TJcxM5kGChVAnQYox/gajl6wNpAbXd
yTnSqelJneVu+LPV3b+03VDNc7k4h+UQlAscsPus6tqCwwahRGm8GpriLscHHnyR
G0CNJa43MrQwoNsnaR2wJo/y4+ybLQTPJmpjAfnysulpXpZQyMSmCym9StaB0+34
SSYAwx/AL0IUdBUBmMs6/kUbbCHOFnTvBPyc+uW3hh7RhRJCYImUknpvlvaJdoZb
nwDfdoAxTcysYjx1Bo0Jxl5qpC0gfyYohLjr6KpuTtE2RKa4Un29HEDFR7CToq9G
1Isha0MmSMgNfWe5uJIcj/7S8L8Ekacs/MUbkF9A14Kjyz44yKkymT9gIdauQQ02
r2TGVNqHTrWDScNqmqqmuXlL82mrIBi4QZQw7EYTsqurHEKuCote8ybe/QXjvES/
U2TRAADbj8UXYVtIUuA5A1ZNwexLlBDPbVtqen4CGhXLEyT9PKRq5MMLjG7jMYjM
Foe7BMqfIdECEeIwxO9jHmpZ1c3W0V0r11THxPiYCj8NI0+SHjRSeAX4hnpES5BK
8oI32mY7XfTPPWgJoaROVmcfQukxMXK0PvqDuMb0CGjw1pxdU+KroAc9qcx/5ZxG
rqyEFEXqWkcSp0jvVMBRL7nXREcQ/djue+oakz0Gde3jyxIhCLnZCf2tBaLNziOS
OBtzMrKx4jHu8aUHqKiEa8jOWbq3W7xUWNu7551/lq+ZuM0t4yIbeSrXXTQsi2aM
mW5rXdn8RZJGDPCsWOzoqnXXEgkF7NCPdWuti4n8zvW0gdB2kRS/wHCSqOL0mXGA
bd+rOSoH0ba3MqeU8ujuHjotbrXIN1bXV/E1YPJWnUcKeMc2FwTpqRkgCO9pOnsx
f049nvEjKVXoXA47Olp5I1WlqCH7t71a7HkvFikV9Hh5483cHGNNocr9iHp66Wd1
PLQqbweItQtcp8J2Nd+PRhE5v17n7FVcsF7vqbaI4Ce+hOxTOU7Ch1PECQjHbp53
gaWd8wTn/Sx8c2Q8AJKU7pKT1iS+ITVuUw1oUt9XoB86pmlsmE6vpml0H581pZbi
Sh6HDRl4bxr1dTVli434duUOVtOgAA1FmzPhcZhVxDnTee6XEV2/wck8d+RpjkIy
qCmD/L95SPP6w8FbF2vZDgXNggmi5yY0IJON9Mvay8W0JGEtB+dtTHKwFKkgHMoL
bbogsjJYRrILJXf7OTbKY40ETmTzunz97Zo2oU1sJ3dmHKt02ejOtD5dR8IVVD12
H0WtAt2wQfcETeDWB0uK1CyXFYG5i3GitDsaPAe8BIVJzB4HJ9m/3jXOCt2AhznF
+UK09Qw/fKJ7BhweJ7K4Qkf7XGRPAc+cG8jlnDCSUbXNfm7DPaKmcf+G+1t02KqX
KN+39rPlcSvKxI1cgaXk0QwMKsLGBQ9QC4iruQSJ0Hn4VHcr5rcrGePFc13L40Gu
SvqV4d9Y55pyjO3juauUKwP+6uSQn9ZBrPynEfqB5LMXtoIN6BeUw+Z0mm+wjll+
KoDIFmRx4bGHRo9EcmC0iOYTbAV6VFCm9ewLnPQvSs8C3xr8kftiynThcjMeQdl9
trpLD0hxWofrfmF5ojZEpukJxcjiQDSn77ApUPAHVD4Ted1PFym8mRTkp+IAkf7a
RSVTl7kl5vJTlNJmNaDCuF0Q7uO+e4VbVM1llD9DeNbnwZ3tt9sBIeuDDorY6/IT
j7Raqlouh0tne+MCOy9U6pGMrE6D3kYq1bfpFqCjRCo6ZAljECXKR46oSlHZmR+i
O3SK5eqZIZCqo9ZYsc9T+42n0oyByPjh15vN5XqsOOIYi9UAzuT5dbZ8GWE8t6JS
yDYPOtMtp8sdtOHzerFgkK3BYOXn4sSYjndJPLL7AVfGnPFGYYz7f1Rx5+DLAqoi
NNloFIV1UtQ/20YYrp1jwtIuWaSwcG0scM7q3X2cNZjKkFZ8oHW9ocEa1gXQvrhy
yq/IMot5uuqox9jzWL/dfc5Y2Y3aLc1k9/XkJr2DpBg6YKCp87TIOm5HqZN5Vj3h
hGgqPWGwfutmcJ3rqf/kfhy3KbpUWpRMH4z2eacgQ55ohycPi3fU+CRnwb1F99xE
MkSQ3Zw4t4/7cI9LWmx4kdt5r+JUYQav4XUWEIo8jV5aEvNnaBFqZyIkxYSBxnU9
1zMMyq2WxXZd0GNIWtU27HwaWoUhCgwzFbfeQdfoMDqiPmSHzS7J6JdGpa1ijd7s
A9vP3+Ovu40wUvBzrsJV46hCp2cMURwsgQ3W4s/Hqxoev4ql01QXRIVXsDcQp4Dc
gmUIFAx1SsIuzQHlAFcoTIBzJiI+1+ZxMJkUOaoQgmvs+TjDfddsDfej4d6QREEI
CmvWz49cEBzq1Enj5GWkCEKaehKXX7G2JT0V/Z7AqJx1WVaE/MUazb+TsxEFPDpt
Kczv6VSwEWRU1EkHHVgvNwFOsMxh57gaNQ6himLgE3ylqTo71c6mOzbDtouQcPDE
Jac4W/EGq+T+twl/xLgA3JeI/EA6+W3Z/fG/peEhtcdwBiruCq1FrTDMFJpSkrIh
T9kBU4uX6WiWxvzNbkfnM8kygCUrd5L3WAseo9oP1KbmF22w9D9GRZOAFzyLMtS8
tN/5EH0Sn4fu1yl0jgmxk3ZZIeF3XqExZsa1JI0ak02fcw4T7ZCEmcRi+xdvxXA/
2eCtZaNGWJ/CMUn2kuqCxtm3Qj+foJqw8ZJb+0KXT8lR4vYXeTkUHbfL5hKmX3xm
+gNCwLwlN0aRaw0bajcBax5PmvBUnx/JRfnMhP4ZpRbuyrhLFGsLaCsF08Wyjwqc
boZSPMbEF9u1X5um4aqdfLV9IL9g4G3JOMkjlkJEjAd58QMhAL9PQ19WjMRBd+nS
nALQX7+eBZZLKzjt/aWxehTUYPnOrPCWlZW1CjxRDDuDNBj5pKz/KD9OBqFyC/Nx
TsSzWQEPXkCTuO8AnUdSl+ktbOOxv426DXvifPh94LoUy7mz/mGgcNRtuP+nLao8
EwQ8UmBOPFC3KDkV0S5JZs82+AxWueOFgo9jFNdMf/+x23+RsgyX7D6p8Mq85N7T
yvqg7vurV4bofD/ZVGOZ/gr+0IwaPr2cUIQkg7bj5Tpcf4ruafZZGr5JyZNZZa1m
QIHFW/6DKOan2RMMMpdok7D0WS9b29XQO4zBhrr0Zi5nnjWP6XlblA9lpc6rtE4n
YkLIVWrzUdjAjLmmCrdPj6MsoeiNOotu6XcgJUS/DvyfKtWGJcTHN78pIxyzjtAw
Mwk1juH2hVigOPwnqZlNzo3zBwBdSyDi26oPmwqCN//8qmBTBKo6/9i7A4aKgHwh
g6Y+fUMUv5gamKEtSypTvWolpfYnLoM70OXxvzT4G4+1tav8K2SN9BHD4ZQ45cFM
XjONEbo9toVfmtOXJyzGLUGnSnay2IUco9twzT057oq4LcrTPA6tsQtCCJNgtIs1
Bb6euAQkhlT5lcVnsGrm9BRetGgxEZWNHR8eD2IDPeP8ym30WgQsmwVeGhJzPum+
W16H91Zq23cKukdgZ1vudpXWIcbDnA2zctt3/4joliQlBd0ZIbgafj14eMRevwLh
T+ibfrFQQZuI72soX9iUEYvF62vntNcYHNlvtdilW1qS5etPNS5UBHV1LmtNkna7
6Wo32AmTkKCAgIlxjF28hsNeI5dkFwRX/sdZYfnvpUd0X3+LXABFmWg0Wt1IvJBG
4HoQpnQEhLkFKsSP/2+Rb3xixe+I7cK9pbezYbv98+qmcx6VWmMW+TgQU4meJUtH
Ovgf75RvZHy63cJ67G0PyuA6PJ1nbiSNca0DNZMMs61nkvXgCsWsh/qXrtlzDRjE
WLjoNVUlqszzioYHqW846Frc8dJj8SaTdulAV0Q9D7tF0kP6CHLCOz64NzGGO2bR
vlZgRunisV7VFl26mcYwim4UiRe9ksaoaYwa4fC8jPAn1STxp5fH7Ey4InhO6UVV
EkgVqSqLBu+ezUiYuP4KVeM2mVPvZd8SiuVShn8HqAVNjVHTR1T7kwFMh12rg9f0
P7W9Jwv2d+50BhMNzXv+HH7zaqoBh7ieNW2UopApWjrYh9XjRMbH0OLuAfzPWH4f
8HL4Bigtgyb7Me+POLuBoGsGahTS70vosc67zsnF9NLMx08khugbYBV6q1yyIaV1
Ew2crMLZuQEfoQ1o9pTkkHmt/FaNLwjCeJBzOLxD0CkGEQqZtSuu5RC62aG8YVmy
4Qj4xBIupCyUC7wckztoVx6+lwXHdFW/9IBoMQ9R71QZ7sWfo3xBlkLu4qpW8QtJ
TcFloBBZhyGN/xBQMlMEYzExFfchBtycLwT4ibDvFwBvS4MTCWO2x/NW23dZ4yNq
MXD7dbI07+8IwpkwNGeN+bypM8wGeOChGovZtZIk21n+fWoLQKPpXmhGW73QOG18
rXMhIsJiXTpeOQ9FynJ71rHaJTgbKVLpaY6jPWkBlmb7otxicHl23cJvdng1+RTa
DTcmjOUk1ZB+onuR+A1Sh5lnx4ziHNrJ0vatIyI4digo2QvGkWaJ7CDdciC8UTUO
v4tKmAsGVXEHyQsPHqtGGMfxwW6HhynIF+deO1C56AaML1VxsxtAIvhVKvMAQQDm
u+RKTWvKWG+lY7/AKVQszpfw9j1OsB9tOReBaIHkW0MNbzsb3FeOJO15zga61Xr2
tXUgebrZSyt4nAi7NykOIsPZHw2vd6XgknmkhudU/D5ULQAwIjFmLU/uwhbGW2tN
0IqLj/YbwEWZPKE3/rmcy8AEQbWK5/EIlCHTSXhfUlvepw8B5BcIb0F/bkicu23b
OFOCCieeAJF1s+1vZu9ZiT+1Wuo3G0AYjGg7lOwCI4FBR2vTfLCX0uqt0ICaJA5N
ds2YCj1U1pLFP+LVSfODhyJE4U2wy6P4qei43/N17MniBir4UNqbjXM+zQYSC2K8
+wALgmDT43wx9EUaas0mH8s+LWJCGD+09y/RxH1LsrvwO+ui14mbfZ+3pjK0r5zr
t4ndoz4K0CZ1+SyXH9jiaV1tSZkdavaXsAxh69bCt5/7lqOQZh60vyqg4dlaQQSR
5s/XkTRhkjq1B6qfcDOyKk9Z1JfJyaaXoxq963CVLgW4CuR/8qR3t6lW6Pwe0Gvf
+arbKRiSj0Yt5KHaGDdECnRcqWg+xjxeti8HzOzAB5SyyheamM3MS902PPQ+CwqQ
Ku2t6UyFYsMpPe5GXFJCBGJGSVrMysUYpSKIu2tVKPUNhj00yNOl2596iRArbC5W
Rwp/6D5eZ2EFzV6BhieKR/MqI3edWR+FF3y/UQtZ6aw2sjFcISRBcv65VG71F0Wd
/bej1nWJekXw1rywKkornV3Ah61Jdf3JLmn9C/UKS0kEJJS54hxTkOc5i49VZUvz
5xKSK+vbru4/+oEPv0B8CiDfeOg1J3c8TFoFecbMgEm4LtxhrC8nsLo9GkPcQJdE
ip5QqGWk2GsnL8Qv3LtRqQWfNyj6Zq+UOv2iHT0WUrhHVq7TCdr4chZWIwttmdbq
boCC2fcH5chdr+rumVeM2l3ozOlJyWlfwAdhoy11Cph4Wl1w4nNafFV8sI/83dTm
x0BV1emjMu88t4tMkwyij+oT1Z/LL7UMJQKlURfVRTWN9Itxfo1kd+87GTElzP64
Gu2Ncg9lSs82RP0d3Ca/YsA8wlcd6lGecYvUbEJqMSMnX4JxIaTY4aNak61q0y3+
6cs9/23h+kIEnOInOOE+OpNyAbLsoE7KuF4AH04670mMeETpyZSfOxQpy4mCK6PL
tu8DkRtUqFFiXrWDo4MJttPsWqwwf4YZPhZ2pn17xc4B10ZajZ9IOWZcWrbKirRV
+nKR7B+kLdKP8ArQMPhixnmNzYa9WN0vCNeyLsYCdDgHljw8nyeGgimqzCqz4AVg
J3f4iKOZfQ4vW+tufrE9ZnWS0ECkc8K2bBC/F7m0D4aw4dwwjwhscrynhofO6PMW
ZZbKzoCtkladgEYsWr1LY5ZVBgMkEqX7xkOAMsYVn7IBxwTYFKUfl1lWjyjK/zUF
g6LPfHk2hZrTEv4F3cnnZ5IxHDv6naQ+ABIg1hP8x+rM26Vn5sOJ/rI2nJUvsSal
ZTkESrrL+OnibM1sqO6eAjiYHeI9213PE4LPhPE5Z7Gg+p11AGEnUKoPGOIWk25I
7GdUr75aEhNw9TkItKkTlnnne9+Qxs+7wvie+IzwBcoSsA27ig79eGEGkXQstB4K
NKuF1dOjGVM7s4mREftaGzI8E9Ka332kATX5iXmBP6harvd/22tcAsXJkuamCZaM
TYQi6GfwAqhf/gKv6bpmMncG01CV21qEKKIjFSop5fPtFaU6Y3WwvXpppGp4Xgc4
nIwShPduwbrOMPGNIbSQSYoQXNnf1/AVjUloLEZ7K/Oa0YZp2uJc9Vv2FBRI2D9Y
J574lZKjYqH+Wh9i3kIRFK3u1Uo2HnSau/8umjuqzmE5cxSsm5/hUU8a94BGr4i/
94BpSTpAqf5qHgeWGUsdnPf/kLfBpfnEc3Yp8Ggghp70hQwx7OtV0erIF5EpO/Rk
I9LmHYajGkwr4SfEpSeSG9wl1I4G/UaSU93ftiLlUErvMptArloj2mA/WkXsZ107
2olffOIwwu9fsMoUZjNOd1a6yy8ojehpLHaXzb7UAV8EqpZGB3hC2OS4aenipg4d
dwzSrecvHQpaE2DnpJPK4UtvrENIghy2G78i/M/S+A3y1ASnDLQT2DqqxzisHicV
daYpvPWh2xkfqqf177qp8KoOpEnAHTJeFTuBdZrr1BIyDcbCNjwYqYFZ2pucPxZu
69rOLeE8NHiBd0pY9JD63TC8fguyEZSwr7ytcPksebY99F3u2OEnvox7XdfJsKkt
v3AMak4XgCJwnJIR3w8AkWjdeFuarnY0H61fX/GU/zUEzECoGcfgbN8i9su/OUBt
h3O+aByZDBB1/8kN9q8uqQpFzf+KI4j6MfGAW1ud6eUiTEnJ6dX1iA5RObl2TG7Y
3wJnpnAcsPmLPXXByAS1ocFfplnnPq63zuUggWbPfVz+R8nkeLOQaS0OVbxX9QHf
jCjnERj8QQ4yIHeiHfxkQ+rHRy3whq1QrEmrECdhG83NlyO1VE+ZyPIiBgEO/DMr
FndyXexTjnfu0ce0oHboX0VxrgmVboc5bODrNZhyly3ys0wTCxUHqo7gGO0pdlaG
TBrA3qsiL9GakCjNKm9Dn9YYiZ0jyiwlZJ37MeRqUuWF2VwitoOqVnPeZHuJ/Dbw
wy/g2aO6fSBEwOTxM6G4Udhw1C474BJr6idSsaiA+iLG/pjDlz6N07CWM0VVf6pa
Br8U51HWHBAETNs/MaHus+1LfqMbGlpSmYa93gxTGEBaR5yOcNsX/VYl0gEcnaHc
87kRZn8oR0b289uphowNci0pyTgT0O8s7lqkPDFOQKDGeFgW+TUDmz55PUxHlFD6
Jmpw3fgbVD2m90D79Y62cwE/E3dhJEyiIWviGkNVXChnZGODFQCpSg/xJko0s8cX
917Vsr1R21Q5gGEd7gnpPlrlOsc2W1IP5vNSwnGyVJtEOhPLmz69Fyq6CGjEFY6/
UEVqm2M2cTda1Z57e5UK0KfMqwd5/SwZZV5ktENrJLGkHp0aabnFQxXobup92eZ3
CmOl1uSA6qIJKq+JZ8NSsKjh8ZYuRlrv0+tu3vXZc5Ugkawr1aVhGQM3tgU8O1LS
vJS1SJOizJheJKfFekHAz2OJWe93Ge7cqtgvOf+M5qeJESjMz4jMVr9Y1aaBNiAF
a4K+qgkbdlRkoDmlA0goCpgk4X3sGlKioiXo1+2J4pZgipPRKHQiNy1yDna+2mgO
YJA+lU6Fkyph8vptuxnJphXxb4dQI+IkAT3cEe64rj1DSoe3aiEwDdS61ykfWj2t
53EFdX+FrNRo1cSDvF0/kCPqfegvPTnY22NYTqAYLzshix9NGkaMdF7RL3np9lmt
SK9+8QjmEAR/BO+VNOxRanT5w00g3VMD3uu0tGLf2po9/wooyKzMP64VOzss5C+k
GQxh/QFZ/vADcOIIy7sNhcKWF0yohKRRJZxJSvW4jX449C5Wm+DMMIbCdR3nbn6x
pO3uBS+W21oFj/V3XwIWMfqKFHlN6YbHg0VPhsKAEi3Il+GY4Sa2mf8c+q74rX3t
eBLKKbROjqGEmZpH9pCtVIoqXmd/V0ZRKi9u4Tvusv/m8DSCmY+T5vm4nNP9ZXu2
PhxuFY9X0PLj5rlbwPUmeOAGauFVLQ1BDZ3N8BY4kLyUC+nafrVktUSfe475TjYs
n+e0DU8EfPyfI5dNi3gJnb1CeJFDFvZ7HvtVF41SHLowjmweGI8F4lMh9ZtK6kmv
YPF5c2yljOoWF3NjRcpVnxj7BL6uTVEYvPRWI3kLTlIz6/PgzBAL5mahkh+s5s/Z
zsipJG4BoHUFsUUkBWOcieggUnXCoCEcofwgG75hc36Z3jPFvcn2dv4lVfULjxU9
9dihadHTtnQWP7kTiiFzRSmNsnG2pKRfFcItW+9hinvME1HxAqoyyt7DVcjfskhF
eoQQBEJjLLNqlvF1z5GjaUIVCj49siDfJJ7trvzWggp0HiRrrCPI8Ehp4hQXz3ga
A/9MNHaVoRwOTrgkaYDL+brkiAbWF7+GJax3ZdYOHOYA19iV5dc7/Trn9hB9KPjb
faMJxdaiHy3ZJdORPy8hT5/4cS5MyhLLVfpsoYUIqq8OvCmuWz8njpXDJFUh+3pQ
6OL24jy/lQNsLa1V/eMaorQvaQ4JXrQqa5fgZFUXjl3d7Aom9OTtk5s8OHK9ZcAx
cTNLhkKpdFPxC89VtbROBeSMDGG5gnj11QYZRoNXbUhNMP6RDEOhnNCUFHy3zq0Q
LirIy4Tyf4XXWLWXYFvTMBrEc+kV6rFxsQoAnDJutXzEkclMF46/4uUNjeelYdwu
xYf1dQta20+/Bb+f2rl8MI6ifsemkGuWBoySLLoIxQSy6BEFoF+3FCs4dHw0YNXI
Hv3oEDbd4Ptzf7/U9qZguVr3FxjhLfjqdT6mexSbDVSeaI5zfTxnM9MScgk6nCib
/2QDLDRV6HwJdvYtzurQKI4fQNfadZeup7OHSRrpcvhMiztY/8qq++Phx65QaWBM
X7jyi4rWlAq2YCfJXxSVvExHGTNi2pWPfQC28YbSMWxCP4ERM4H1PcO9dDX0viXa
iVOYAbZUmSlAWahON2889GOyZZRFOHWD7kqP0ic/oonEimsHTlA+6w8Makmsvdf4
K5LYcsdm6bfcc0gn3FpFSUanm+5tDpTas9Ka+s8Qwphx+S3rP4bYSKUkaNmyheD+
Y4FxzvW277HQHQMglWz8bYHUTjEwiL2PX0olj1BAaErOh5fK4qpFXOy53ICCAnzm
ESjaoImVw0ZeY6gNFhQ7D4DM9VkcCsZVLpmOK/MhkZRKerY8lSN0mokCqAvyUm0d
zSGbPbyw8mFayhtv37B2uqhwW4XYq3YeO5328jJ1F6DPpeTha45rERpmUwTj32EW
/c3FvAQroXQS0Q7bdnJx5GOfIXc0Bm7khtj0CSSPn/FQ1cWDZgSgiOWW94cVLsji
pJ+3KlabHwPcRvPxDRULRPc7rQdKguubS2aJpuHEOPOYjifojMyDJSFCCy3YaO6M
4dZwYzNnu3oIf7Tce5uxmEw9785Ut6paPHz64KG2tBZpUOUbuVZ0IL/v7szkS5nD
lkeAcK/DYcO6yz6P0Wh2cNm7xPLD+VJBfKY8829NVVhQvRXz6VfqHMAN/SGVtqdd
SFXO0brBdOcBVkP80PnC+0JjQAFED7bQSK/5r4FNxVIl8930KDT6C202O/eHdCOL
iECJ8Ef0UFbroqocQRRnZDjKzMth7XIzZr7LXROwaE45lTuUqCWJtY2HvyF3aKqW
Hd/ITEhg9db4Egjc/LHJVS6BjdRU6u23JBzsVMNX12bOvucqANmLZYYatt0FHup2
lMjIxYCns2ESPvGAky0E3s+nQuOuXtCiIyNHKNJZmJwCOaY2Rf0BXaWHiuaeJHKi
zJQ0gYapDovBAPhPfmCbsscRZOroJstORL9defoIyGx7xKz2g3MJyfEtfL96RX5t
P1yNrPLae7HmQqB9q3d9e6xsKR/Dz1w8eCoMn1ue5uQNEnu5jqW9nl5b2WsBqXIq
Mvh+racCtgNiWBKeX2vKx3T2+ZSIjhvBzbMbVR7ItGsXFX3l7WpEHAZreAelP7Te
KKNWEE4WNdxtL3tFf5+oJ79TcyqW3iPp5Vx2TsQpBrwHFME0NLR0R+MVa52PT80S
x/hAfJKWitqTPX61gqmQg9Ddwz62U+bZNWeTAh5DD6Y9xQ5Yz6xrtonxIZs7ITOK
VKiRQMhyFHeKOgM1eT9jynjjpD3WNtPaRgX/vx5F0WWDpJfNbcp8PZW/VYziwPNS
MU8l5ibalqoDUzMBcR1TQl3ASkbMZyjNEMW6adoBzBfNZp93HaENJH55xP6/jLa7
D+A93r2tR+6CSpCPtPom09ZI6lilUxl/FfUTsB7k7JTlXv//cXO/OvVV2V43PP9q
Cq69FZAGAfEyEhrB1PzZnlPGvAQZZTvxINmZeNDnXgwg423btRUW+0srzfXq1hZR
sgeBG2uxHOzNbQgeTmAIMI/cYE3/0X5Y9K8bfvcp6DdhAN3ovOiw7pmDL279DYx6
gxvAq1bcym8Nnux2Yn5kpB0aOKx6N0p0aWy9pj4LXYmqPJqxIdzOhUH486S/2V3w
uNm99Dsjhkto2PRJ6s8UGHzDIc7/OgeJoAQF6UGKRz9qqfMH2QNmyXL+1/oY43xK
homxNWlEeAAY7T4zR6yGKgfPki5AImeS/V+QrOn7olkagcgJO9ycNWSG7tiNrvdU
9seIgfTdEioxR9tA1n3jp6RuD65fwv3drgvuwGE1ZUNo9h9749hHRO1iUC25yamb
J+so3cwJwJPH0LfQglrOZZQVA3U/2CfC2t5mJfP3EzHeF2ukVULr17Fv5UHowwX/
MIYQYrnsmvHhvWdCaZ2KjIQhjeObqctoaI7nW301URKgLElyxChTYvu2mglqZuA+
6XS526P1adLC+65wUS0RUKLIFcKcdeiMnpSFi0Yp4GwKh3TaTrSRFw+u4/12KmRW
RGdhZbcBE9WHzegpCgFnD6kreRvM7bP8obu4EPmLYCHIfhGsfuY3vXJSIZUz2XhZ
9c4FYPYsb4EqhInFrgVPVflHC6UNOCQC6BViHLkLIaq5arS5YkzI40ngvS7GrQoC
FLv25HL0dJ2PN3SOowkRHQ+sYjx9Y0TynkfWRHhROOhBWCorjP+Fx93UiHuqxB6g
0tBO9ggEO0ntHOAldLb0FEJOSx4ZivhAopqSZkERRqggp6p1vMb7R2VL2FIwI9Ux
lE8X3OlHg3lbYH1m3ejxbmJ+KWwlaIiDRszJudtHVhDWpOOOZtRUskoTyZ/TFCbM
XXNRIQYdML51EtvsQpVviMyYJyQra84JEa949BprdgmAN0ohTEEPKTtYLon8Xwid
vSDJlKyz+LGJ9zeqDblpul0r0VhUh9rybweg+pyUynXrEQjUfjS/GlilmmBXuNDe
k5qbzyS5IuJ+cQp96tEwq8UFX2Iz9Iwb5sK6Rovfz4tDfi+5asyv4RlJ/USxE4Oo
qdTB8bE58A4RvnJgDJXnNG9EptYbQxLTi90XyIIDvTJvj+U2Y8K54Ox5zz4BnYU4
7rKC8Gs4/WdhqzVmhL8FWlUnKSoPUIj2b5r6oW2figUoxhaRM2X3UtnhqmF2dp8L
zbQgqei4ok4jQ3f9Tfg+r3iB34FOHceTNSpBsjYubqJsHeQtoTR1mZgJ201Kp6+Y
gzwvj+7qwYPKHUbux4dTdAn9SAp5VDs8jLKzn/0gVWZzCm9nf5EdOlRcZh+p8E+6
wzcoWq/xmOkTvZ//w2GMTX4V05LqMdWVsp5E950sx3ZFtlMfMTcF+DTkZixlqszn
JKvDKd9mmz9j0vGLX05OorYN5fTRUWbzG+CJWUvEl3v/OAOuCxqs/VM6o506m6Da
FbP/7lUgBmuEgY1x45iFegHR5uxUYVLqvShZL6VWGedSFxnqNeDb1dTdtmXcP/bL
wu+yKd7fLE8ev/DBaLPRBuaMhI8QJU90oHbx1CEhsRlL0026UjZ+mPjdvI179WUp
zWxLoA5wrqu5vIfQnx3MQ6zFcCMKFBlkhjJjMqQXfoA0ctuQyQCHNsTvqY2XCl++
aMXu6ef7IboFTEME9D+/9YQp3gvBCrAAjAdZlV10/zQZ1ZrHXOwHVHZvohqTLXqX
FWooZcn+JWzSaSqI/8OvQ2cSw6LTDkDJDXhTe568M+JQXzNqLaeF9ZCSQ4DA7PkK
PLT7Gs84G4cEn4CNu8jBnekoIP2ykdEtwqqCME8+RNxRJbRRDjilYhvyyy4j9Qx4
ordTS09OfVP9fWZmlks6MYLlkUnZN0a1QKHlzOtkp7oVIfcB8oHEp+45/iDfN2sf
uvv5DTpfpPDRyyTmMvo1uXbXRssdN6GHrkGL7S7n68FQFdK1vR+pFbe6T7U0r/67
1p64B3UEeS0hL6cx649ijT/NLM7ja1jRVHsk0nc/ZsajE1MZdBY9QM4/Xjvjs+yw
K1x3HqsZ/pkK8soz+78j5qv7jDHZ/POlVKgCEXNBRMIjeUkT+Wb7ARSTwfq1BAoj
I3yBiSu2doay+ZFejKRz1waYF5zFEkse4aopF1mAjz2bQFuUHa7O3Ffe9BTj4f9g
bT25eQiw1JUjXyxnYomSCLnGtgo6ihiwzNKHnTETyT0W0mhA7unpF3Li6RyF8I1Q
gVdCkvL88vOSKkFPciE+n/H86yjJxGBa5izPCf1fdvnG3huXLxzzzNyQRj0DAPVk
8z7s5pdhh34uC1X+l2ycrhhA6vlDnD/+kDOSQ7d+YEMDTR5S2herDOKUmAas3L3Q
Xjq/GUcyGUPtUDsZSt2wdwzGVNgyv/vWbS0JspcJN9+YcWhNSgz4zb+6Sr0DtNDO
MlfWIkgKzHXNrMSkrS/7uPbxu8QRThv2asNK4LCFx/vV0XmUtZne+JAeSdo8qnIP
QVVL5mGDRsCD+ayBoSqSevdJD7wBfekTKRO0+V2xDgE8Ip3Gkl16PXvSFr5lM+3H
yBaxF8uMdhJBmfjE/RjrR/brIJE7/FFXIJOVK9U+3O2KVMfR0eMh//XC12TXg4RZ
5m3kuG8svDSJ3lPhrW938ZrcKSCPuLXNflk9f0f3oi30gp0OY/7js36aBLBmsyUA
MCF6sq4lpPmp91C503JfHhMNfsfer69rKJ8uWrxriSIZXolBBIv8zXxGT6ML4nJK
FjemdchN2sk8cRnDLFvrSU1zCJkPkOhrn1m5SOFyIBrvU0nX82ebw9IKO899AaZa
8iEnsJHiiGAbPYiMdA+BPP2EBKFxF4TnhMjOfkgzKtyMmWaSMgQPuybHvlr6drC8
lA8h8Me1SY+pFWZe6+w8UwCrm6bjHjr4nqh/s3xMq2vwGNUmvav8JN9Fo9yaUW7k
2cFbSt+4Ozo2wgC9TQ22vtBJPvy+uDlj5Vy9Z24yWnL/lu0hMuCrSadNyFSlT+Y0
ILZAVloF3csUKz+E5u13h+Qza4DNJoJ6vwtnPwk1LlytW07dd5vRRca6zNz6c7So
wyw16sgGf3BPsIZfzXKKuyHfLOedXyKGJ/rW+lUJZvuHgDT2Y48d5xq7X+oeYJeP
yiOyouYinvvketB0bGScJnoOqtL7EprC02HltlQu+ssY/+DrZO0p17YBelStZ5Hp
cYlfyenWmW/MvX0dbDkMtZVRaf2Hxyowd1eWyY5FA4mVYAec4BldZRCbvwaOA6vu
n8EGzGishf/lUJ3YaNPKuAs0WeFZ2dGQjtqzTC5lBKIDGYaw7wWs6oNbIz/kiAc9
xOgLxuliwzgwGuQKe6MkpnpgIYW2ibR/HvQiPhGDhm9sZcwtmIewtQ9t454kb3mu
qjVRBEh/KgW8JzcDzGuRWPTQYy9nxRN8PsGtxYu3PrJ8S4k0eistrNGcpl+0MBs1
MIk/MAQCCZz6h4GmTnEFRfJaDHJeVZXt9LcxDDTVf0I072FC4T4iDmR/e4h4CCXU
YG8bwjSVKqfmAdEp40v9H9SJlfR3yTFKeq7UTxdMx/hDuRitqnmH6/r0THVx31Nt
y635CXc0At/EBxIGk9mf2rpTZLwaid7xGd8UM27oTjmcbktciVtLGRVW9bxrAUMW
yzyvozx610F/YAkVtxow7KOF5xRZhLdxFIm6oAuXS1eCVhdso+t7US8v+XrVUeqr
S1inYWJ+0LD0IOa7+mYimnzt7XdJ/56W+qbo62FAokSyb26Jk0BjwJfaVOHSU6vx
Pr4JBamVPsblYZyWo8H3FCye2dVBxWC85UxAXYmwdps+C2TyotEp71OhdBijv2EZ
xJgUxW80o1kPvzmDSGU3Ay61OLM2JNayFrW2eNaYXy4AmzdGpANZlz0GxQPPvVD4
IKGFta6hpWw2K4eBsbfvTK4WQ1laZwYpBPv6eHEFNQT7b9y9JgJQryho1GHsicx1
A85/FO3edEQh0DuQFltJqU1fzHRQKio5u5zt5NkZjhi/AGFQJWW3Re6fqQ3LgtTc
de6c1Jc7rbD6NPVCGBjg4D5TbV9GHzQvwpCUn+JhTUiTExPHP5to3Q8hy9gZi1Sj
YipBil7N7O3qbp5z4cuQNPUf5b8glwSdEuCkFlxR1R40gfE0iNGAbvvp80ZqDgFP
0h/0YZfTcgzdln3U0mH5S2G7q5Nmw5Rc781ZIb/BrU3M1vWbWkHZ+FBlmV+3nvqv
wo8WNtS50IBATFSVu2P9+rLA3U8RdRo6m/HWSyiiKzsadzDicMdGF32V9TlzD+wu
y9B5MKoIM+OOU3weFN4Ld4dwrMcPclHD0QU8OL6OzoYMOLWcq60CDuFrR66UQ8r7
4hK5I8cmN9AKvaSXfhhYR4F6aj97YWz/VM0nQJUEj7gaImffkxaIUhVMVnUxZN/E
C+Q/Q5WUr6szt1qH2XXozDTol3EMzOYWolnQJoWGyDM/enzrj3lyfgBvEF3mEzBL
XB7GIF7gfrdnx2q4zPUKbdbnemq6W3rcj6hFnCxeNQE0QzYtE+CdxODGHVFAE85R
0t1ASrw95Ye1brkPo9coT77HsgVdAK5RvgtJB7kbkbNX6y3B9GMF+fmsrh9ClrDv
0++1kHPpMPTiFSE8e71SKNz32VlcGQLNV+GMKPp8CSmUFy8YmsMgt6bPH+CVHvuK
hOABUTzf24pedNHg2UAeU4SZrLRY7rURjdrJdTAMVEL9993p+PCl75cUwUH52FCv
iao1qo8kYU44F6vh5ybUvr/Twmx+9lemzstxLDEB6xkzy2+MtYpsgbNBjvreCU8W
HziHYhlEAXemWA74dPnfIKNc1R71CH7eWCE2gapgT3/dDUEzDNotzq6BcOWNPtxN
Hyaivfrq+omIE0DQGGRXyAYNKmRRcQ5xaxff5O5EykD0RrBpRVZYr+m3oHiCywoc
y6uj0Q1hkSxeg/NoXgLnWsR8Xh49iB1sQMLSdfUUREh0aRJC92KInH88K1IVfKDz
BjWrUXfWW0THLkWTkzLOgLKGAztIk34SwC8e7kkJ9tDO4erL00Od5iWkVHY0YZdX
XJge+VNxl/w7baJs+fqeqsNfxVqXozoFTEX5dBmpANbhAi8cNa0UQwFmwJdrnhza
7sSAaPGkuTTJF+3ROjgXjpgOSAsFh/gY2zCDJ6At+bS4MkG4klBZLG0FbOyR0PHm
EhNX+y+Je3WcFauGvMRPe0DwvL/+z1hcBouK20TPiFEx0bkhr1TJCguKCTcG94by
MtII2wUZ1zJIMOX517r8sS00BVmECHGQTNWOS+rg+jm4aAuCve9WRHE6azLYiS7j
kq8KRP57OkeZT21r3zUPzGXkFdTHTzUHLWqX0GkO4gE179uN87e6IZ4/0O9yr//d
riy+eEys0BpupL2HPRi5a9fITpUIP/rI2r8mvaJhO2HSGBWa9QTd5szd4U5FHEAg
r7HRDg7iwj87pgXYXC/pxigfZoKKWkI2XFs3/aGw7xFJszFgP5tx82NFiUzzZ/aT
TXqBtvSpDytutDAQ/p8lX4BPR/DBoEVeJ5UnbB42W02fIpJDj23Qg9bUHl8IpQew
vZWC2Z1pdwY1qYsrMCgIOgZipTpuOtMjXZ7BoavsvjVkuky0gUJeFYsJiXfqJlht
C0/412gh/c/iW32UJxvcOCuSbYQyrPQ7sTsvBqePATysgpRQ6DCZzBK0b7CGFmiu
/NwHb1yNi/WCDzwxabn9IlAHrIVFUmeN9Vk8+M164LFcBZZqFyUwCJhsuVf2UzGo
WFtlJuE2Pc/RYEygeX5tH3QziJMJ6OQ/nhmjVAZY3/yXPgeQklN8aJ7unwY72eZ+
+Qm2K9mHNK/okNkXKas0/U1TqjAC4WTMsQuNIxsiLPrfeCHSpiWqDDIaZujjxM0y
kfle2XMnAFdrveLp07YLpDyXB3JDe08EvPZyoG1KN+XFJVY5+ZbCeSb7MxPrzAFD
MMwMoyXthI+bW6NXOi6IyVmkHyuwjdIAcJ91WozdM8pe0G7RH/ezM132+/yn7ACE
JJ4rOhDIw6aKfTUjBK/dd8poNah7dKUbbeCE62LFuTgOYvl++Hvu1chYnrnZYxxn
jbVpnk7P6QM5E+EzEbjtWlGPQMcxBLsjVB+Of5jjpOWTyFVNtYu4Br9Luc/URp8g
dXCaEJLC1fvf1ojB7ITjPxDOnQz+xi1mYOEtzj5e9fXmBpR2hf7+28EqXlJLtmBE
XuKkZ7ZnpavYFggzb81CZwN78nqKW62iYlFi+eckqP5fxZ9U+nwzD4vd9typf2gM
8UJurW8n6/OmW/oyPOXtDEXUmwm26CNgg5AMKDi6cI9uJJ6GKdEPrBs0/WuV4vip
evqi3uSAQIfok34XJDD0lyNm5TcIABAiXZ1WpR78eLPAER3bZGygzj9TkfsJyZx6
Mf9S5U5Nbum2q4Eqg4aRfE7JQJvRPGhoSf1EwBnTp1UmTd4FA2rxsCJBTCD6feu4
bYG7XxKGks+wkTVEqm38q4M6P1LlPbEp+jiMzwUqEpnLBPXZaSvf3FgjHNyqvQz4
VSgUIDFfBp5Xxu3EWmG4WryNyx4NKk7lWC2FMgdvDEL4lQzT04/Qr8Jizw35AJKQ
gMTwUKJXhKZE+X4UC6KwFisEmMc32+DdoVZ/AVVl1d90mtISRJoETeoFnSZC20Jp
4m3u5DRUtnu0rlaI2YKYwmDmi0IpUGiWPhZXkQvk0CbPmps4abJ9FnTkLaH+9BQT
Ub4aQWkg6TmV3nldAc4Jra6GEKnA7K1j34jgqau9787tOXq4l0kJpIP+UfzEIIWK
ivrdOM6blWV0Xfu+GHCub024YpgTDVSJUQPPAoAuFX+DwBXEc6gFOP2dJjLvwUYd
S1fCN43Z1FRN6lZGVOZZhkor13a2nk/g5Oa7Cb5iDmHXoQ1bbkHycBiePo/5A6r7
SxlgSNztvB+C2zpUS2uzZBSpdQp60DdDBIYLx23nwavlgsoR+LRSdG2L/fNLPTEb
jn4ZutMFsZKRUrP5Lp1DtEb0p2kJ8gz5wQcZeD0Shgg9LFw+/ZDOIbLRGM8xOH5M
bK2DXbBmy/sRGpiJZ2Lw6ACSmdq6qt4+7/pTRnfCe82CAel5tPjo+7qVgSYGgTwD
S4H/NXc58nFqGebGCp1DE/ZMq8ciuR0nIWhO/7WPmFhyMQuGuocWs1x/+y9V65WD
fcTg9UJUSB9yYHOkF9mwArLJKOx6G0ijpq/hmyDcog2eGT/fWTt0Pq47I4mZl3jd
QYdEvGmUWPc7ni31f5Z4HZRSFbDbr6l32pOhkhrs4eFi0FNHWLIqZJr51fCSJMIJ
Qm7T/yYV+K842jVrdybYArGCWa539JJ99BxNx/2z1dZmLNiNct7fX7YewkxjY0qF
9BOsBwdPrGfto8Aet2aZuVBZqwY51ZOGPUyi1GnGXTYE4kIdQqgNza1XnAp8HGwE
agkPQ5H5RdUuz9OTu+I8B5Bf+F9If0HqtN8lJKzALxaTJV9xQLIOUbyjpzJ/sSIQ
mnK0CScGIDakXTIxupFvxLhIj20xqsASL0oNM+eQErvZQdeBylNiqiM+7nXgBynE
w4DiqiORAstZ6eIqq+uEgP37ByszXXWnXsHfpouk3j15c2xiZlxjqUYJgShhq+pQ
35WcJQWetXoelOVnwtlKdiagKUxetm9YTxs9+le1wyrPI7Rdv48CjcyQjlzOElI4
22GJ26KjDI8TsJweZAPu2Q17UqqudBGGe1ULIkUs6brXIbpkvVYgBm1phToI0jYj
E38Zr52LlVqDYP098oUJlcTKLmdw1EVhVeyGng+BPspdkqZnhplBNjsfARbX0aGZ
khm+y10XAdRSEt9VoW6gKTpZGdgZblBq2WtKOAK+nincoRCOBj8dv5cH71s7iZxJ
fo6+nxMI3CJgFqrrqYhuAe+bR9ylZsv7qPhO2m9p4MLAwVFNdJrlHumHMz9DiI3T
2FyI/VIyjoHs3epS6ANjuyLFVBur+RC4MRnMZJA7gC3i5dndXVzyThDqvpafxCmq
oxD1gjm2ZrebGsGRuVDNJHgHbxLrOdPOLhjLJMUprxBNlOypLw98g2dy96x3r6qe
tdPeIAsMLCD/bTYiYLenzbhpKeFN/zwunvK6gSb3xxu/i+2nmGMrgiE5pHuaG8HJ
fzCCXia3rGGKJMZgmh+wp5yFK6MyXiuMew7JbybdjIasc4CYPuWBoZ5q2rbRvDn9
pfASv/U5AtwpRYmWDO7oLS+dGN5SaqwRRqOhoK5/McB2YBGfLEqNPgZF/aLebLPc
0il7VReiHCgaxuY5nV63Ufh+iPmbwwvkpbckQlEz1KfSbY3zkKajAoRT0f1An8t4
ZKmywctE0NN9mv1u4BFgfU9hyot7etJdQWLXKy+vaKssPaQ2MDIMvbQ8lZ3i54ny
wpi3T6ULVxuJ09ZAGcvr2Z0xCbnisDfixhWdmY4unTjJ5D4hN9xFfKKacXHJOPzY
dWq3JgmbjKj717RN7Vg9rZVVUfCkESbowNgJAZOmq1SKIE7cU8ShhVXxqoEL2/zo
B5EL3evvyj7y3UT6ePE6u/Zk0glRIXiM+glLXOQpHNfHSVinL+ljKfmrfMIVM12W
LUdhz1+rkaL3WRlm5w8if4uCaXazlGgXGseT2Z1RlzrJ4o3dyhfOZNVrh7sWPCkM
VdxtM4IzaQReRM4i/Ni5W9IINkU82XVwF3SOxBkb+Q1EJXCA0gIT18PCkV3qVCC2
pFSJinQKb7WVej9GLGMBoSfuTjFl68KvcWiQEYCpNL7+QE8PZYNwK5+S5ISjNM8a
fNJ+LYI4jl3qCQeLH9s+/qr3SpZDKF/Nl2tr2+bxDb0D00pP7c4cUCjSZ06G9Wi5
KzcgsUirTY3nmX1LBNYAuMK8u/R1Y7/6f0aynSaaKXa3CrSpuoCV6sgknC//Kdwo
9sOpJutfr7kcTljHdjsfgwWvmrHnp3Cz9xpXHOTR1i8nu2fJlRNVIiFedDT1iGNf
rHoiWxe/nEKbQS7IwqHYj7hc0uuxsBOyjQJiBE+BFlDan5UD3VwPggctWOeTUIuT
XDDmdiO04yeK2cCSGzjZO7SomGOFeVhYLardsmwFcOIqWWlXFbojJ/eXUj/fcIww
qTOUWdjvotsaEQ5H+IVfrX0isSCd+e5T9SAISouSPcOF/TyED6EaWfM2En61HVkx
IpYS/e6hO0NWHLDaye8G8+D3FX7VbC8Qs7qYXkYuWhFynDep0leHS33zFMrtxiOa
OVYbgbzWr0uRCMx40mW+2vz9y9DFyq4F2394MM7Q9geNPKc/85v7IoB7NjfMa8Dn
sW4nwlOFTk0iL1DdYf+ISb2lyUARTszp8t7gq1Uyi7gTCXvbH2+zK8cJtehDwTu6
fCBnr2rwL5u434n44TFJ6fFFUMx3TibUufR6D+y2JnIx5mm8W6nf70lsYGYYwQLj
OnNzrvkcqX2x9OQc0SBKbO/d4tiS+/QNnJSlKQgZUNgjh1gFJDVO5oRXlrFEzF1G
GajpQXOnjHTreE4plKpDsSJcF/XVAsQIWDNi7SWylZT88hqHn/SyObH1vmM52n4F
UG0PLnxnoGGDzMHH2V3ZseFu5Yr3VI4114A+KKl5ewE+2SRxlLpDLIMqoQzXgig0
5UNsQD/HHrEHa/cfHhYo0CXz4oakH65FPumWaWL1UCtJCOXrtUbbTHm3OOFodaKo
bp3ZmEwFTrATcpwxpHsLJT80o6qGat0UVG26Soa0UlhIN23xBlxVRa7sENngKAn4
+uPaFvwjYQXyefrO2MnSS0dT5xs/UTzJPEgvBUqZMOnDpovS9LD1mF0WX5dBJ/oV
8+QWU8pk0yOEiICcZy4p14xfz7tD+1mRfXPbe463JiZgGlRtJpIbMRGQ7bEBxNzQ
1MXuLYI3XgkNnkNYt6cr3zsXCDWfo4e+8mrrwdbnOrti2ibiV79TN4uPIbrtHVrG
zJ69pjFICFrvRkioE/5rUTbIO05WThn5md6r30MApzmJuKl2WB7dRWVmAqjok4Vb
jMgQ9aWDDR5omEUw8e3iOdmSf74S0iwJlK8eiqTzFkM7GswzVBJ90AhuybFFs5/N
hRkhTj1wJzwGzWUof8ofre9Uh/ABMm4zkJa5vFKdwT38D/9XqWgOwKOqm+0j28rM
Pd18Ecp86dn5iDAWiyKUEeth9tvkcxb60DD+cADl69n+6HkPV8/sZ6KuytXUszTe
RMQWb4QXJapjRwSTi+gAlKlAFRrq7wtUgVe5mGi2PE96W+OvkZTzWeMmQRKQcJHD
ty1qhmaFlmiGVSh209aP1aMMhwMQYL7rRvF2c8A2yKqGL58aWhrUDsNtqC3lg6sX
K63JYjAcppRerW20y6tAqWu8uI+nUbBb15lq4g5FHKbA6JsJgLsN+C8vomPZi3xc
qeTQJakF800NRTJ7U4cRozgb4hiZFAZfvTJOSVow6xOrkO9fzYd3SRBGhz7tUiJ1
wV/JYfCDI+3MdInM45l/KMVn94n19Oq6xowCPc4nASoY0MOmt0P5n1Xed8XOy7sr
tIH1dEDmN2klkfzy8apAQJXTQlkX+KDm4T7lU/nN9Nr4cp5yR0h4sRqjhioEw0M4
/UEEhGs9uFmH2FUw5r0JgrGprKMs4bWI4XnS89kjnhvw8I9h161xDoF7nnYciHpp
olF37gHHcMfkJksJMDg0IS6Xriv90G1RBOqLo6pb0tDfqwwOnZuxX9qtimTn7Svm
mIhbw0Iqk5jPouOUcb9o+DTxmReagjvt6t6JltAoYSdcoYaqUwG79x4Y8LhdibQt
H9e3ZpHRWtw+WVcwkPAtJDsayh0xbEtbO6ks4UGeezwbdFjjD8FeJ/Tmj12hbrSH
V0iOZgQ8oos94azl2Jv/tCqDMaeTDsqdKO+NyOUlmjMsdIhH7rNV33HL1Eyh7KDY
uBJvL6L7wIu5kcuM4NXQwUuVaL01T1+Y8HaFv49fuox4ViEHWo7od8nmo7924Gxn
XG4Wjzm4vDm6wPWOUFo4iIgOytBbtoEP5jBpqCBjBPnq+cHluXSGIZMu7LuEiK3V
OHIM/dBSROjyDlIR0/Jia8tdNUMXXxESCFF+Fxon6K/nJ1bG10aP8VIfmQdSXMgb
YvCA/ILak/+9aWl0PrT6HTSJnO/5ssg9C8MYSduuidi6e+3qzZOTvWatNSOpmUAD
XzM5TPCz0JwHo5cV0hL2O+cyHleeihoAAaclHKrSkYCfdkU7GiaV2px36Pxt+AUJ
PPHqiwfS1Cfx2F4f6O+27LtfdD+cuGC/QN8MPFC4LnfUwDxBMuI8UOLwN2soKaFf
cUaUH7UBe7THQp3I5fRUXkoJbSG2BYFzGKXvFC+PQi1JE8aHaDRg+Ms+eTR0ninW
hYetYtzDFSbZDqHwmgIrz0moPCa0FLb+Hlqjx8ThIhMHQu6Re96yQz4H1V+wDVYH
laCtbsZLXJ9lljvGf4Ke/VViKoeYvDGpQJp9aK3WwKmgcCfQQiOlj7i5V0+WgmV9
HZXc3SKSPZGd3eryJVrYCiTfkcedocpimMCT0k63l7RNMY++JFiTcD3eTPpomxQf
49P0XFp4+FcxDnPANgm6HFefaLmSn3kdTImxS87bt7bBRAbx2u+WXEwUR9MSklDp
Se7nhAIOC5st/DiHisCj40JSuwh2wKd3w1C9Jz5Jpxq04DQGDrVEkrC3FXXwrQ/l
977iSHPLoI9cdlCd9DzvpnuIr5D2Ocv+M5q46HiYNkrEuSM1G8vPJgVAgt7MFH1m
DuVhAlxtfms6KiJzM9jUHSdYx+eiMoCXXFIMsyQsSnmp6fKccoufroCB5sGDlqaI
ShvLmFWQy0podyU+W4B7l8XVJLHsIjewiw8B0QSv+ueNoHTe8z9LqK2JkdOvOxpm
0lJh7T9Nl5iDwZReVn7TVpYRlnKxJHD6A0beBlxQqTS/gKFaXrPIMiFS+sl1Yzhf
C8i1NKhD+DXyv4DeJ8/tuE8M0xrchmKgGelyiG6y+EAwet/wT+VT5EYUpK4CM68N
WLzLy6HQIGDqWgz9N51fxFcdXrKtWhB5gYu2myKRhu6WVIh9k8CADFfwdoeEppQL
Xuo2GeAzNDR6G7bN2poWa7zN1CfqpmBxtna2NRoRFc0XaCo+cRUebDTm5jleIBn8
TlTNl3tTmXFg8iWEHd23KQ02EJENHPifsjelHnuJ/LM3sxWfrxf7zA+BoM8QR7Mh
yBWH4Wg3dfgCXw1lIlppljgdZonhPc9qQOE2an/9xG6egOIOVTCjOM583L+wqkXC
vIt0JEyKOo9eyYj4giO5kOMpMUpjI3fmyc2U1Ir0yHnQPoWDOVi/n06o6AzEpVeQ
Dy/0dBkwEouI6aTq2EdFok0KKN1ncB9IlIrzqamoHOg/Ao4a0NXCQy9QD8+GGVun
roWvLWc0YLNGMkQhJUNDm+zVNUC/UGLg7ytn5jDazyN04l9vOOY3OB1T64iZ8z40
DeIDolOtoD2lJnsrgkuDt+eQ2785uPmxNnho4WSyX9RiSF7pVijwG+7FUUIiC87V
UBSqLSep2jrMJgvBs4PijEesU+1KQGVKDocjvz30NXmsXp9YaD/5aKFXtyNwZ+ZW
HYYsGZUakdwLYiHBtMng8ZytbFCnl5qgOWrnEKekM6XXKwnhx2HJHDaQWt3t+l/A
mivJOQqaEHQH0wt/pBvZ+LtkPiAqlsR7AvYJY9q/3a78KSOkDbopc6f74Rcan7ko
S83KCUergSz9Adv+8kaX3ATkNzuH+7XUnwIQtaKivtLSHdkefn5Wcj/jA8QhMKBq
2ThSgdClPcj0VA4D+eDYXMBu+VADYmG+NE+sBBG/k7+YikmLEjZzFI/qXObuIJX8
zwTJvrtMw8ySXPGCgerm1IU27FL2PVJdEuArWpBsTkxLn1LauQFJfrjnGshdiGCG
KwTJFvasqOTWU5Q9B1yBKAF+gkYIAhmFFjlbUp/SPxbsdkBOHCzQBzH+nL1umXcP
CG2PgVXtLxgxIpCzyEikUX3pdn4QqOJHos4ZGDdAc9613yJBVz7yAsXf/9KApi0v
amTEFBCX+O8c2izbBRtsu2BGSh4RN0qf2sytZW7Oo1C9lUKNn5d3LOdD+s20dC1L
eC+6WU4qm8MLJ14bk8H3lOCfWZWfkKIxSttQ4yRQxunxB8p5XqnstZup6aLjg2sM
ZKT+G2p8NRTGDHESWEWUMhLbwVpxA9Kc+X3RVKLC8oDvtOCQN6QMpg0pF7WZO5UZ
cc9DJVOFd7njGiTf0N7qENBQbbvRJq6rdUHmh6XYAk56O+2A7QXu4UTbyBFtAWjY
AcJvyo1tzcRYSRUmhcjYsj4OM/yW4dXYck+LM8KyKFElh/1S1V7nloBHr/eHo0DJ
W9+8DHj0349HNMX8ACwji77h/pmU2hhcEsQS5Sa9eAVNWE6vWg0LupgrfLhKr8BT
LmTxcifPOIgpiNje5iWaOz954K3EWNxjcukoVaZoYjYpaiywYhRZ0MuoGDPT+sre
kG7kalvjvdk5XJBKAepeWTWOz0OqU+XhmknhUkwz9My9Ii5sE9iXfwQnvqjxStgU
+3uRSJWn0JzXp5t4hfC+IC0ZTM+WVeQ9qKbh2w/qinOjorR+F19lZP41LlD8Ufst
Y9ZaQYQGpnoySQgjCM1v9Eg2AqGqNlHvr0+tHcboRBJdL9hWBFZwoYQ+bbNpinxt
dM5L5flDvpjCzwNjWJTvrBj/XArycJuHUh1FVaYsXGRp711dOaIUi0m79vgTY6fz
LK1OyfFMaQs/Y2gLGD/XsOgj2xQX3QwpazCiMkWqWQ65xMTW+EIOvCbIayvsYusB
xPMFl0dxs9SEZMsYE2MZOldRbnKcwHYnn+NleTSSs4jF91jB60tiqzuscAK1unNV
92hBaLjdC8P6baHkewGvqVxKse30VYro6WsH35c8UyBKxlHLnDAbCzc69/LjJ6y0
VOKf3/shEU+JEjicpfbWUlt0phR5hJBkhPGvHTX8TXb1kvPunqqlUBes4y0v2tSz
iI52fD2whgMN0lcFC5sXmQGBNXJ8Rjth5URzD7a0Z/WmVv0lP8n3Fp09Jd5BlOFo
UxVheJehSDWojV5T6wtMwCfyFoV3wv4Nojt3hajE0SronqEPD8SDoWe1pyVtCRm2
Ui46tXzzIuivkV8CPJu+Fmz1cWm9mQa0YqG2BYSopVSW++zoESX5PfcgdGJxcYAT
66hOhwTp9iz47fw507W3Jeyndzn9yp09WVuAgjv153jrd+Sxsy3Mirxc/G3QP+sI
DHUFmYX1zjgNuPHLjowvwvUQFwWEjLW7/BloRn4M1pg5/z/xcnkiU8R/aNSfbP4J
syLWU7CeW0C6/E3Vi2xt7ZoEjngCJ1DW1GAisPb0mlv7eOfdAKrB4ymE6aNY+zXy
Cl7G7NbYgU9k75+4FCV0uQHw0rEmqzbZOU4oSsPfLUlGYzdwk5l4U2kn+29uZtDr
bQDE1GIQvnNyaYslX0i0BnL0gGI8YwmvMU/tqjVpWS285wBRNonaanFkKxbkX6An
vJUG8MIHn6/u8sfCYLwwinl/HADcUiJqIC9B//dNxv8LCVl5Fr0zVtOsJ8ZKkyUN
OvOEo6S+hcbfEB+bGArn/RltGprwxYwfZMTs7Gg0OVwQac9zbLPWZI7lPmtLtWue
Oc4vPlYZXS7v2eAQJz7ADjp5vLobWgdXMALYAbIsDVFBXksFfeXV4kRkZIm/QFlh
IyeG3PYU+Fonzk+gT4S4hzBz+cGigjAK06h0kFpO/I2m/+Hs7qbrIhJAr9wRQhyf
wdWz1X0TskI4qyO4WUl+iMUoDUPvnYQpvFVfnJ1R4v5kzg3daLtXQcWjrBZjYFiU
hY7ZdgrmQjMKuRxDJj1gb5rgg2GpVS+jl7HUouAldJmSZA81BQj5xkJepHuaJCW2
GRHQVolstOWzBpHLDkXvBpHL47bZQnTo09zvFEVDcF1nPRkyrwHTQQRHns5f898m
y0VNPM6zKC9u0glqxEa9JYCVuXv1/SOWK+azPYaH7LpjJf3rz2oTrNWQeoV9yADI
U07E4w/vgywU4vuRWDX70woIw0JFD9JKsaotdxZUeaxUcqquDdumTF25yTB2cmx0
+B5+MDeajZFpvZNpwG9T2QYKHlhlXMy2TuekPgjHsA/7uP5IR9T/s03TIy8zyKaT
8s6SJk0VcquZGIBf/fsIgY91GmHZehaY+yQpKzAtrXWuX+FMsVo6wif569g+XWaq
3pYos0Zv5bQLdRpgSLU28QbYLozy/rS0GOVjO3oof4BStHBlTqWgaI7npwbM2W+p
khutYuY6AwLds0XUtmIDFKYSuRKnzWgDTh4muesUvAVSEuRQmOFVM5+CYpv0gNRd
ItGrknpcnUR6zbepTLm0mg9qTGdXoBlIbUVTbVQNwfGud3pZ1v0U0JB3VTf7gJLS
zRih6AAV5LR+4kIy5MN7QP987mTK/TEztBu0oU7MB1kaMmVmDgQJ8jJxgJPaMEAB
sOiUaQpVCQtqb5z3j3iry+5ww6NDEwIk26JHLL5xfxSicetWrrB8PR2bVad088PF
DWRMzTvlAQb7E5YD9JDp5U5LeAAQhzs0V0LePvUaJd/53YUeoX2jRgXeib3WbRfa
i/HcMPUayxK5d5Zm2UIWiXm/9UhPZrGXTfwvhYzWHDRqIlvcO3bPaZ8m6wOV8V04
qV//xqNQ3BFqCmjOIKymQLWnoblEj6TSKRawRtSG0b+B9jEOxgECwQnKq33nEAwz
tvtVEEcL1ApfZnwFSOZXvWZdlw2O3WWOzHANE16iU+8j7+gLIdVcRu0jYrdvTSdx
JSET7f0fqmxAhRUqp+G+eiXarnHS/meMii10D1Do3PEIMrMu2rlkK8RbPx4Rk1Dq
h13VVd91pvHt44ixUVJ/jgEbMBVjCDCwpCN2HUFBvunXiDbPuMpWmMrMfAui/gyY
GsDBnizfAvY1EKeYjdKbDjvOCyLV3AxHdPlx+DYJw3L94ghOEkuMt6xAvSaVlv7W
X6SP+Y9ESBuK5s22213lsiUTKZ3wYHbrepX+iNxIczpPOJ6/DMh31QOZAwSIxiqB
s4r9jK22JchtryzoAFEWVOa/Lx1ZtM4iBWNteRLlH0hQNNOxK/wWgXCuf11YMkeS
3p24f9C758q1oJLABxPlxUNqEYHGDyCW/wFFSlElrECZZb1zsZRFQ/uOd98+JVmE
aGnIjgFEp50FLHCwSfHPiVlrastBVXBQEOU5YTtdjf0Oce+ncO4KbSGOqKHqRFqR
QkRuV0k3yX9CIab0AtEyLvEbZFiPk02HtiJ1DWfrRRA7U36Dy6q2umG9k6P41F+1
1CO8zCu4d0/o45LutHKozLy+rqNlJPXVxf2+IJEF9t1VujmTAndNysuADQBhP4Ed
JRWyjK9f9Q+oQ6lIk5O3nwrqqPLlWtPoITbqv0lBnFDu0ShHG1Tb2cmcpByZG1HR
P0w5M9kj3zT3sWYeXHifDjljTC/8PiuvG0Swz2P/KzHNKiyUQmj1lMgHE8qH7dSV
iOWi/tw3orrnfnKwSQQHSbOsIa1vQGoc2KH+gmf3xt79+Qoq/Gw2/I5cMetIqmgz
+yk6DMnsAkHx/wW/ylfUP1liIfxCraIpKH8nYZ5Cj5lvySVrVo/ihhmpS8ZZlj7K
43hzvHwv749MJbRYepr8LlMLXfGwYP9jLKahCamB1LUUrrm3JyKEXOcUfh0MJHvm
j1CvdlBTeqfRfDIpiAGmdyUOnZDvtevf8p5Db4qCMqWc3BSjWt5cxqa7a6Aan2ef
I5wcDMS8LJsV8IbsB+mb/7QqNPfADO7G0jnrvOUvf6Oq4q3XKvcCz2Ro+JsQdzhZ
W6BARY0HaLe9LvI4FccJXbe3nMzWqfXfSwt1cXs3+G37Xn0gaq9F6IY4ctkJE4kE
W3MkCmfASD3inWjpccmQygoxk+UzVHjhZX6/vvAX2uluXia0ZgivX157ODhmvocL
SC47SGOpNCNs7A4ibOQKtqNwKOXZ6GRA/CD2pV4LkTmN+RyEgoyzVMR9e3Z8OwFi
8rV2lMwWf7VUTbSXJHLRfCeKTkuUoXKIHfShvQFQgR/CBs8HF1gKP/ZsuBBqfGst
ZBHHuYJ1w5zHir4D1It4oHiAekIqOSZjQ52XL88aP43YuyRr0WeaKrGdjYBXOR9Y
dvsPtjywbPEndqqjVKUt+3AySuy7w/NGpLDIB3QWczpbwxgrSi1LEGDf2C6hdSF2
vQwvovSe71AqImYTmXzsrdn6uQ766XaiH+wl7lhC6G0uXxirisFgZgF+OM9ng7HF
OFWuKhntuDvJ/ClyphZ67A3podpOqYoKuWWaHejklqn21Ijy8ftvGuh9+Fp9ssGQ
XyhpzB35Dbh56Dkkx9kB4XYDf1sbxMZwvp62iCidGPopUuBlyT6TFntVSfvZY5e8
l5x797ODH7+aC5PllSRFmPqDGBVNw5dXhB022TEg+oq3j9nql1Wz9QTlAgVyFdS1
yiK98SGPihOJIwaQVk9Kui5av83ySc1da+WZoo7Qw8ZOr2ci3THk+EuyKKUcSjY2
pZxxjllV+cV/ar7LYIS0sqkjvF8CzUEJ3qWZRRJGTvx+ju3r1qwsPjzOEjcNRJoc
uBpNmI3uRUxtSf+N/jqSqaWkNPsMLHCEBYM0vTRQSFrJP6eVtEmpy+i07h0RfezT
vixwUqkOE4GN65yFujRiiGiyUKkEHWWIaVhA0NX4DUFnOemTUAmuiXBy2LN9e/CQ
arUfPwikW0LFql7FARo7tstPBqhhuqGQbUmgoBcJcGbXnayeKInFV5HACVFBDhH/
2a9TGYQB2bgkLQMZFxAWcaW5jcNIS4daXd1CBR9Y4fuzbNUlqsSRZsXdKeXxTRdM
P/yi8Ij4rxmJ6czhZayZZbtEcttOVW8oe2JOuPPkYAeI9mVnGEp6rjj42JwrB7qc
AMG8gGPxkltWG2OolPkz6iLG28ZXlJB3POmZdEsknnsjoMNyCPCpumS0ZJZP7FqJ
Ql2x0p8zq7EdNNC5AavHvqp7pDSqwzFHlK8ndWePXNXjw5C6rC3WDucmabBqcIjE
ZqwrXLFriQy9QJ0eJNEL1h+sifN1b8zziqVvvACTbKZxzzhreB/C23r+xHRDGXgQ
6FmtU/Kxfud1mkbKaBkzsjrYXEz7bAc5PG4KwVrF/0yWTuptoUb9f6NJ2nB09d3P
xGnrzwsUz9VfRJ4gZik/MkwRZhMCyBQsYTWphsr/lWwAUCeLfZjOW6molX9Z8AA8
4qnfjvaWtjb6EGVxHi/WdzhpqZ94cQHT3rIhrQJIzPa+VRLbNtavBjPX6C9jKLAd
jdR9FcCo0JSKJNq5yQEf8D6vxwhz+UQlPp+PADcWtrUbFaRzYAfFmBoGojkN68Eg
08sHXVaf35IEue7g8TuJnixf0W7TIC1EhYKNzCFcAlTxwldHoWW6bXWX/A/iqdgr
TqPZ9rm4V+IR+faSLR0QmsPxFHGID3hk3tAhMQCXC+dodrcjjDoG1AtSS48g4O2E
KjHIB4+x6yKPFAsdzwiIEGzJ1rFTDI0A8VPd/ew0qSQ/EnCmChpGJUjPGlwARnlx
bWoNwxpiLBrUmmg4IQsa4a7MZyTco1GoCkc54YNLzYPtJEQYPDJZ52/9MJGHwcGV
Ot0wL9Z40nq2lVtu0hXxUfhI9PmAUnWd4SJkvqDSwHVA+u32HNf+cR0UBaryC7Bb
c2Pwd1dPnyczyZRYjY9xCvLXvUYm4pxCZoBbCqH0+mB3iNmPpx+SQE25DXWF/J2Y
h8HABzU3kBUVwBFbZ+IODXkhSRSps2rDKhtuelklbMArvQOgLXmD4rHHSt/dzesR
+BKN0nBqa9DFycJoGG6TTzdSPjOQaw8k6hADdUBtbmR0ITlwAGLDaF8y2OVNBhWv
W6G5tuaQelOKCQMmZEqbY4PJJ8c/XZnXy5x8X3LescxTNxArLkG3kE5ufpUvyzpF
6kkwz09dk7dg+w8nvLHprsSaTvSNsoPHu5FHIUY3/6QIy8J2dnhsMqFxYU/PmVUN
B1PNaQHoXL/k3CLrTQ7+cfUxbmStr6iVSnfyHIF2LE3nBApnrK8FCFVKgs8YlrRN
J5+y8wU2Awe1ggS8mDAQ0W5mAoNulJT60mYfpO23aN663GE1RDA+UGWlihC+JUAw
BqJAR5K9IDXL6oNR10pwkLB9QvMctBSPBfrpAP2diQvfqXGnkbTNZDY+Ium7oNVr
IFJMz/9x4kyIjU0Jm6A41PGTNFwYi307296/Eh/OKYeEakSbaLztmELbpFT75U2z
qiPOGivmfs8R9MFsN3X8325gnCRTIm0NqeJlCAlFQ05Kx66KV1qMp1C08LuM12bH
qBoAqE0sYaARkgxdG1n5BKPwdkod7ajmqFdKdqk9BVU6YTYd0YWwxZP5TuNoTCGW
BHW1fpOcs/ZTglm952EsEXc85a1S7lzcJCEY/hzIQB/Vbjx3ZK8iNaDOAWK+bKHC
p3IVLPnYIBGD/DMnwRZK13BiT3Rcmz8g22q2GrcLTW8XvCJxL8c8mdjzUGto9GD9
pqLx2aNsbXzZicvHiQzUFQPEOlnHT0ngKq99jKGMeP04ev5xJiyo+LV0wIqh2wLz
6LLHnu8WgRlwSXUvgaNuiqNSiSVmZabCmzXmEXCsvOS9Ca/UJlxw8sBnlr+bvBfz
TQOnRkQcA8tR7H/GeZ96biP4gW6wY7HNkFduCpU2XwMCa6Em1GyHVRn8jGdxhknw
3p20Ra+izZZCfrbZaI/XdX+RKWQ5B2db93WWBcbYooPOEE9bgpAQ82diYbI/Wzji
HeyXHloT92woaesfWuMqPPmDEPuJddMFTO/sooeu4xMysY1IPlFgKIQvKfZn4Sxz
bwP7FfO+NU0UoOL/PN2dulzgq1ASyJj6c0E9lHKZNrPOXJEvBnvTQCOH3LMzuQCq
FqrcBuYqtwDD2ep8JWgc6BGMHUiVoQX5k1G7QfOsQn6XXgbfjXKaEGAIHGhKZ5+I
kxfaPloo1uIkNc4kLFLoHTnqWB31Kc7CX9u1pErkJTUpDc3dmR/yYrein+VoaoOF
GhuS+7ZnUG0az2FtmYz86WAFnhw0LND5xgmhWdq/XNzfOM9jHUB/IJbGFXlsy1pH
OTL+he5BIZScstvPn03sxM8nira/0Z9ku8cw+VOHTeZw+CsYV3hpVmXq+SljFSMH
HkJLeTIKnCOYPtPUejcAA3jUhkLdQrn3qMn3omTsGqTyBaWnA5AUrZfpdAVbpHpC
roKN9H5NwQcvAyPkKeb9qapE5NMAkMv62JxsB+yoEuBXRDzXNu8K7dHO2pFpH8j2
+zQlTFgtj5e7hNah958b+AtuojmfvUOqrEJzbQ+EUWSM/EfWYCNbMYxsndEcXXSY
hKBez0bnSbm8LioSCCvGZ5XuKVyw524sKti11NEf561k7H0fBrEyIhc3LRNhY3WI
STNVcZcs9uYz7uo1ZBqWcX61Ozy8VWb9J74XGltCOhdC7TSfjOJ+pGO831uZOyk8
t3lnmkAoaxVKHwOUv2ccKR++t3GiLJTJL7sXIYoZ6anC3kVyWpHh9oKoKi+zU+/4
9oDGIYhnzpuHYyKx2SMI+YTNWut+9PUXbSnEq0JZqI9GzmDPeYuzJIGQueN450g+
o4dahIBQX6Yz/2SCl0vJ9AIFD7onz21Kd6qu8QaLO8II243uGQSRVl+ECsG9qXFj
1NqD1HqrVLmFmWMh7ufJjA2ELAmhbubli1SKMAND++eMAXFBLRUgNoG+I3dgSO3k
P2lOWSsnSTK0vM20RClcYodpEHgco8MzfuKO8Shrn7sovw/w1c5e4apEOPQoEAQ5
ZFcGr7jPpIEE2gCo7d673YUrnoV1sfdBqn+k5hU0tEYExqDAlxipyX8ZRrFltNyw
uFfcdg+42Sz5Xb8BolOwT0kBY5N5Dl7yX+E33gMrnybSPXzzg7eBjEJka34LscEv
QlDhC9zXZYEpfKUvE/kLxGQO4SBLMnulVB4Boh/MILp6jLnRLN+Y0Iq69N1B8Y02
guHOCIBUWVwy3dyZvSM2491ZMS+TDsYA8GnFgUB1DB9sycQf1WCs7Sm4oq3Wkape
gt//l0HD+TYATf53Y+Jzf3eYvfmBhNC/UZOZWdy6Eu0guebH6jMtJMmknMd566cl
uKgOS7IKRrOgqy1TEtJ5dmzq0annyO2ol+AkRk4PFtceG3yfO4OFFlTPpk8I1Tkx
2c0r/+vuVk2FslzubHSIi5IaqGLJ68vXBb4qxZ9MdEqhiAZygPIj/2DG+ENRPAmH
5GozWZwmqzDiGYSLBWZ9qg8EShNAsYVFlEnwV7mjC8AcMXcbCRunqnXi3wPGjO3U
XkIiCL2z/gbqnw8v9Y2uIbdDNMRYCMSMvsnzaz3qvcoNMkWK5XzRdOYmsBLKXdqO
VVlYxVFAuccNjRYiVfGCwk41g8qoMz4x1wS0Prg7HGnK6f2ajKWD6BlypJOmg7IP
j1swCDA17VGoNUL4X78/BqQas2YWleThgsgvoZbeaFtm+9KqjqfsFobRQqG/b7rX
UWRr8E3Y8tiXX2SGzjWxy5+94PuWGoacs5ZwlosL47bZgYCNSLZBR+KPiEYPe0aF
ZACG/GJp/PCiZNpHMOiSJgw7E+bBepHtN1kMsHrNOr97XQ6v22060ZNhdBoPL/+N
vSS3cYN4RCfFpkzZUJk1nZ3XfPpfcTQzwE2w+3azmnbZXjnwzQJ22T+YF8RyXfgz
HL+Jtg79uNYADCwWUvk6MZCKwMV9UD3j9npsNDoJaMv/em0y3HTMSlALAF6/Gjgb
e8XAr3AuhsWLbS1f63ABcpAeKC3B5Kbh6gjcFUfou1FZO2iV5Jkl0C3vW/eitvS9
EO2NbY+1QMHwPae/uXOCnHi2NW2txLE0DIv+6UxcMDNrHGNeDY6nyE7hIMZF7z4n
L9O64fOZWm/7tbTzb71UPvr4zhEHSjvm+lw3ZSmqQ5051rpgB34Aa5t2HXaewu64
E70qf946wcGCzKSbKshicW174JsLJ0/spdc5Cx/MkwM3lfdKhFW9fmLqtMqvA8jV
/B2I8DSrZ/5v3Rks4Vct6+VM+CmZvl9+DUxDk9GQ1I/TmuwqJ/Q0Hd/dUUynw3O1
UgOBS8ylUSc57E7OcPifYMcPNWAW7lDNM37y+rrFOUHigchU4TfVt9spiMaPW1J5
e7zf3MyOKyc6zV6/YVx1OH1tpSEbDOlYjg1gJXXUylPGmSpROTYwIUpLlwalXScF
xpfQyVlgZ9O5pqBHeb8XQ5l3O+8CXrWcvrrTRVyRRTSS+Xf7tfBsZu9tn2fC0dUM
ScUKLtlAC5GvJnz5Kew90QAA0p66qOO/XLkQT/ZYZS4JaEl3vhItcXjgn4NlynEa
ISNEb98oUD4i//Kvefx9B8DdcijwUb6MjV/pBrpw4wj5CCMD58h6/ZuEKQa+MAip
vycu5B2lyRKC54LsnqzJNAiI30V7lqrAbsygcYNfqlRVvoVUKd7+gylIaJMjYj+Z
1IdQrw7CKAbRSOiLVQh+JGB5KX3OBJhfu9Lf46G2tOJoKVpnd3UbURKvbAG13UV2
6veVpHdBbhLlFWZDzR6FgL9UMRCigpKrprqRlGrIsg1sV1TbM7Yn4cLOsnzUJmDD
zDM9Jv+FW80dp3ovrCBQnlhrRviI1SZ5WYf2M9eh3jCr4MPtS3oduhc1IsTLPZgr
4C1JMrbsX7rJHB+sbc13umIfn4txfc1+3wVUddF+O89zeYc/J0rF0ZOv5uuCOT/R
+cvmi+MqMjnOVVwmsP+nfuuAQ339/AaFfGPNsx5TogVQ2I+mEe1spKV20f/Vqw82
Pr3PYXXCN3ABi42oB3RfZpXtUQVQ2nYmDsXJdGck91cHbkQeWlhN+9LmTZliEdPC
DEvFoq5dBtwu+C8iZbbjWR3YktU42UvoDbvjG7TgoyPIm+DDL+fZwlRo5d8wrTpv
KsZ5+HtQRanlnNgfJfj2SCwPaC7yabRKHBNuoBe3x0Tg5BwhiV8zID/euDLDKLG2
9dgo0Ns1dRCQytzdXPisN3vrfiI9X8pOmLPEk1kXH2PcI/6ds+dLr9LKGiO+SSyA
nf+GAVUdOpnReVvsQMiYh3dGPdYKMrPpAESGOAzN1x2rpPu5WRMZkgJUei4fFI+8
okPQsxqPxTDEzeFU0/ci/KX+DjeQhPWo+BcXfiJ4YDHMW0I0eJ64o1Qj/kpbTanB
cLdKxyr7J7txyeKx80fEaiEWF0TFsb1JjFijiBYW1s8Ca4aG1Z/aSc9pAxxKhgk2
dgkpn6o9jWQq/eGo/c/bSBgqu2p4jbIrR32/kRB+8vFKj27t/RKQYNtSf2Bdth8S
JAuPhGiuLcqo5fiJ5YqkouBroPTCHWeJUNFw/OmFU0zgn1a63Ook2ZOzYRguY+2u
UC4HpyXsNiK/LIkZQAds3MGQHFTt0ReRgTSaVwyW42oYNJ+UedEadu+728AR7+5i
z4XBisl2zuig94RIbPDDspa/E4uco3oc4gqTVvqt8Hqzf4xlfzmuJN1bVt/L0o3B
+fuhnbALLM3l1ulO93QsQ0GDCMi++IlZI/wkSS1TWAi6PCTe18wg+PuiGjh6KVGV
mLTDKsOUu97gdUd4Zw31KKBpfXnsJv4ICk9q7md0jNSSqDnUR6BvOlTAZJqhKeic
72YHQ0ItuDMc1JRBvBM6xF7DRq01Uz52P0nX4ijok2uFI34OggawBK/D2j0Rpgyi
uFCWtu7Q3L4u6MqEJR4eRBT0/6XB2DNfjTtsDcVFQEu6MSon84avEM6ZIx6PPk92
7epw2VSLuSTgFaIH2H38Dn7R0ZqdLD9tUKRKtt1R0lcnKzUpMU3ncmGRANDMaWoz
qzv54iyFzOUVBL1EgvtxQUb6glpMgjY2QGXP+DyU+nHusGMqkLfFA0Jxj4dlGJxH
TZZjmgleQtU+fxAhiNK36duvAYfpjElb39gCMFZ9M3K4cw4/mYc8zmSCulkB2Al4
z/MS631V+VRe/7C0aaJiqcEl9ZtccIWh6fhNMp0RjpIEmO8O9zHFN9WuhmfpLbS4
yXz/bSgqF16uGhx5AjNm60g0qUL47KZ66RuMAApGXjBzzpKHbVt7FVJ/nsVszgd1
3SFws43sWPUMmnb+4MWECTxTZ+2Ge+ecFvGLfdcCpcLkMUWpho95RZw9gb+dGdIE
oEXKd9whoSL8vdKiuW2M6hUSCRJ0dWZD++jdlXbvlqP5kGR88BkejorppU05smvy
YbO0M4/8G4eg9A4FyYszN325X0ObBS0h5qZH7lMTKRjjtl1rImIMwUH0Pt7BVicp
iDfcbqQ0Wi2a6JScSd/vCXam8U/UjZ1LJFPLi4fbGoLkgCP6ULjjbjKOZ8yy36Ki
GjvO5DME6waHZGF80kMYNJPAIxSexMmsVhQRk3y40UitLp7gYotu9nGG8u19sdWB
6usFXnpB6ZFj4wezaMfQGK9xF1Up0dLrsCf0BiEy3DFI7yI2n8NVjuy2JBrBDqKH
zkIuobDTj1lERFOpfy6j6KT5pNpraVHku6SZlGK/OPzdvdur+i4z9TJ6fOFFjHGP
G+B8v3nH0o1CPKaF5I7rNJLKyEBPcC0iftp/dunrnczdSjFsqqBMEworrH29Cufe
4smZt1nOuExrp1nNrPbDahVn5anVyBSwXPoj8sRvFvn2UoJZrXJnRrATDVzw8B2k
gnaw1CEBWlDRqf3BYEC6a/RUmExb56t4pfSQSgysVN0MtZM8I4RjWrLlqvbeH7jR
fvpotyVFikatpB/7WEa1ePjsdiQ07a/nVA1Ushkk46mNx4Xq5zN+JaXbFGqL2qTa
sfT5iDUJ5dP1nsQJYzQ4iCkYRJQVs3EQDZUoBIP0C/De6o2SxfyUHm3QZPtDLq2t
2sLbMJQ1heLZoo7fxZK7qt1cBpw6DBe/O7TojHWyfC/r2fNpjMM5LqE3wPRCcdbU
TVhLRtmZsoJsgrRFh2UvXHTy50/bSvqQbzfFLRmodQRSxGsz1obo0lcg6sQGs4hN
dP/NTZp7byYMnEqC/o87eGr8peym5E5GsO4BVDDwwZuI/fIjIK6dVaoZynHt+uL9
wpBc7mJd1rM7cLcJye14X2CRO+tptRpqcYWmk7gvq/jNo6p3HlNyaP98XV7zfLhP
tAribtTY7oC0yBllRecNFGup1T5UUsQmoON78gDI/TbLr6avG8lr9DKblc+am4LN
Mu44/TTX6pWvnF6L0EN7MRXnX9f2C3V8HMjdPbANWrzkZldZ2beq84H+7HPx86Uy
U8HpaE1OcCdOj8N2L312jC//ryi+3JI9BcOOy+6DR75E+gD4zRurg3Lufrw+UuYK
OpE4RmtLQEUxA/tUzJDE5MJ4h6iKNHCJ5wEx9UB/pKT9Jz7zB0Vkjxdrlh9vOKjT
4iYjmMh12Iu0v+hKoRJYD49UkBFckWHBoAjYef2wJAFm9yohqoMdPg1U39PiS8EB
HpoaeLDbW9w/qv6K/OTJbderoQyRThLMhUOALq44BmbEf8M3WBJL6qfQ7C2/E+xs
XST7Xewtnf+cdzg8cxGyLJ5cgk1bFRPw7NiqRwrWQ0PB7Yi+uWw2Rjc4n5fqdV0s
udA9o508f2zlTtha4tlOmil74jKPvLJ4K8dlqFk+XdBrAoucy5MLT2KymFpQwMA7
3LKlxjXh9U4jMuvEsSURZ3SFEShRaD6YBpd2MCQpdf08fZJL2IYzGx4qsYx6HaGF
ukjo9b2BPZDZ3eayUACu5ZdG1E/07Su9HH0RM7yoDTeZwK9Vbw7V4EC4ZQVa9zkH
qhPIgC03ydo3/pXLZRVGUC9Vj0OOJocnASIO7K5W54mEh5HdgKfqrlnjN2oI83lb
EgdpWk9Epov6IfjXN4zca+z9O3WVjlwBOdUqW3QYqbLjxAIfwUTUpp0xoGOJIT8w
VdCTW9j6jf28UYUQaITREAfg3xLXVsm+pfGC6u4I8PRXPq0gD66bjrBzFa0yQbU8
oVO4u0zHW7e7CP7JjZ0oszYYv8HmVoydlwbhTgpWllRe4DclCW0p0UYG6X4V4YTj
zmX3pJlPNfBjEvgIp0nsTIm130p5oDyFOH6j1V6PjkdyFi1eT7/0wSVGtRMhDsZ/
NUYFr6nMzzGiBjSLA47IuGzFXgPlyyZuw/HKFFJQh259KEXFrgZR8UExTT2UgrhD
G6Ayll9htCkDDH86H68BKJHZT7lI5cQf1vhiN4M/Wm7L1V0Gvryu8tXG43jBaR8k
YpFiqAZ0Lt/m4FFVICl1Ct119e6rxSEbVOrNumuo01k6XbxU739MMWTkHpNibT5R
Z8pI/yQDas/U+1vOSpnxFVCbsvLqhf20zx32xjyul8B2RA0+Gab8eRqZuXXzuwZ9
R5KdyC+J3ooOqsgVsbgWRL5mikGSytkUiOGCiNpXb81WexfdOqrc8+P3uQqTrM3b
C3JP/Ui37uY+vorprXS1NM3q2ANXGYEdg8YqGL2SCfa+VoEhL2YbnysuGqQ+IHXH
f4j0R1/IrJfdDOxpkDVNlA4CZDjBeyOhw06GwqIiqnsuVRsABSyM5VWBcoF+mSie
qcVrcxig03gdKvuJToBId4cZkzNLwGhROLK2iNCrp4pfB6mObGXJ2kPOnawCiEva
m5HxhROZNEp59YDzVf3+SAVVIBrD64Y/76djrxW+Al2Mj6yI89mHIzLfQBBJKyDl
OXDHpq2vSrgCTMAl3+siyFnbDzVgHVD+60QEwZA/SqSXLmDKXimtWNJHRbtZOdLr
ZQZFFdVnLXPPQ6JdmoifUZ+xedhTt9Ydc071gQkvKVQM9BsW9UO2nmfq1Ggd2mH4
9g3VuDbbw+HtIwwzaWbwpt+wLBDjJNKz3RuJbqZJBOg0EPrLCn/y78vJuCDG5WEt
jcsu1Sg8iixqF+sVHCRtf1E+oOwQHdl4GC2B+eJzRvaadKWZira/EEFf5hb61TB2
WqGvoq1Pt6EOW01kbg6iDNfHxgsBNlx25QAEInAE1OaaCoJCvrKc2+HEmYY3gKzt
6D0lTUX/8TmieP9M0P2jBmjMcd+ROPprucJFgeNychJqIruAlydrzXTKihMxI1GC
Z8OTggvXtPZd1Sflpl+MIU3LqzFlj2bvVJkZKtePZrjOmO/IzKes3jMnblu0roMH
Pk+N5Hb+JBCgoVNzted0sp/KzvEmiMOlpbrDa/HiM4tRuhOmPYc3g2KzdAdnW5+1
oajlobjOSOgnvcTuCS2WfRgKZoI5JUANjGZ8HzYXxIL94OY04Z4LZ57fvmvLNkoJ
mZw/uEc7u/GzdMbkCb9wlfeS0gNN++K5raMGx4iBfa8pN5pWHbKalg14DW70FUfI
W6hnocX1te4zPER79zxLX7v702UEbrWTUDY9n9BZp3Jxgm3+/SyV24sxkO1vuMhN
7AR8IV4MNm46qxVdpibSVDTFt2mUsN1wmHydtWRMEd3kZbx0x2NkSymhiANzLflm
N/AA2+FhndpwtXEwD2mJ9hMAKP/j4lwahzsgR8mXcxzJStAUmHYXvMelBABKHcgB
eYRd1sbrfLbcF3DSzs5VxDiNBkiQTXONXn4YAo56j0e/fo7UvxHm7eU8O1RnI8Nd
dHAAzm0K+a4GQ/gaSkkecE/r67BiIUf45D4ONT/ooAO5+L26wzqEapZEl0RcK6zA
n3fYzeQtz5VuCEa5sJuWmvdYIzs94uFKB7ocCGL5jropgQdIADYhkh+N3+pNr4vm
6+oimtHl6ULv6/H7MOgrmuCX/Uenvm/qZjXvt4kWZRE/j0TYIBAJ6Kv/ziplVFlS
cY5KXBnvKZ2rGEpBj4wO96UfqY0MSBcSj36xd0TjkSM78NdafSqR9wLHIbPxu8H1
W3keuvyyQIeQKp4CWlsU8ga8MXwj+JafgrfCd9qC30atv2CaNKFYDKGVOkR0EafN
pxbM2YGN74xxQZxF+UKqlGSt4g0bLGFdL78pZcqbstd4dbcazsgkaJtM/oZPDfQM
rXkyV2RexXvv7FxHKnYqqUn6L+Jdlj7pfuCeZw5lnQdoJqycGjD52SYuB7GjiKXo
74YAfXTW3pc3Dyu880gMJ16Q3p7WwxnGEydZeHsWaoVz1dio8sZ+eJNoM9JNdkKv
Sdk7Bn4adW7jI/9TP7Or67+TSbZ3dZhoOKuQ2r4L2AENPcpFO++ld1+5VKqDWSlp
vPEdbuqdN0p8X388gSMLkte48DhnzOn+bkIglsU8wpRjyp6BYkWEOh3fkTSuRrtj
AsaKyDl7ZzYd4AvF2q3K1DLHManR2f/wcL9b1Ss5F6y0EvwiKtMO5CaDAl4ZyrWx
BUFJPxJohSEU0trUm9AjAbMI4YFh/JE46TeZnNIytF9486GBeSXenRW4Nj7MnkON
/D6255K8+N67AApCx7W5yxmAwL3z2Aws60g0BY5D4XZg69b9xQN4B0RzA+iKYXsk
Z6mllonmNjEtuVwOQ31YY5dM5DxLOXIa0+7hpOTxVwgAVqJRnuaNBvxjYj7l/9Zr
xVLMGHHeYO0L0+uEU7gpVgN1CMOrCPbVZLxl+yDh1t0GfylPMO1lFk8zW9/qFyif
H47U0AY4eSD7dmPZMl8IvBzsthfAtjOSYYKWOFqidl0CH9H4ARX1ufTL4tFLtTx9
lFrMhKMvzskT1rAhGA1rD9T6nNV5Z0Ei0V0qZQxskttcXPQgsj+O+gu94tFnbI3J
Tds1bsXl1zIbRjdmustpERIA4FaGRTXjlKWUaTchrruV6ihdw++FiWLfD2Dzoqea
X0/gayvl3p/LTca4wf7YkNT/7SXy3FC9maOVG886nHiBHlA/+6F7UtXFfn9CWCg8
Ly4CVu1Qq28heYbZYDFXPuv4FL7jloqhuqfAjC54O2UEoWRjw5UtO6vOh7rWyqae
5NWMRn1jsy6vUdE4BuTUdC4rf7upioWVXEtErXcI1CqFocLqcU5HsHeXVHq0Mpx0
L4Cd3SlBh0NGydNW8imqgzSpupDxucafTEcrb1tj5Ahf9DotX8iKWkMbJk+TLhZ0
Vxih+3CmSzxBVQMMrDqtsNpAQ/aoDOAUH1nBW4ohu4OtmOf5ETfsh62/ynaro4fl
uTPQ+TpfBvYdCM/x5ULjlIOoJBLsWalAjJsJL+LrTtIGXLxkeB1Bp1YE0gYpeYaJ
NmHq884bUDYD4jUXOdaTUnOq+5z2dZA+yZ6ptylec2OnqTcgWLYM9ZII3zaNmxpu
nx3pRlPq8vYEc+nrOAm8XxrTRSMtg7DY3aNvasB921JLkw+ByXUPN4K/9s3u30UE
mLFCINf1C6tNkC0H9za/DltczcuT3ILHmgjQsbO9dj4=
`protect end_protected