`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzY2+EFIYXUoRGNXzJ9ubqwafGWU+mAErY77eC+3yQSII
wFF89zD/L+wytCUnsLUqSQ/lYI4Daosg7V9Bc32BdMe3WJhzHbSURIyj5Kq/pK9R
jDzJXwRMCHeCCYWI55erYT1qhh8QGG9SZ9LNoNEOg4BP4DWUO/+0JJK7iFilB31q
ZYPZkFlpd+1IqXGlOAi2RN4VSVjqqpv7sVPEdjpOx5M8/PALK46n13yGA2fzwXzk
27D/AzzyktSzv1kyAspTv3UZcJrvAjnb05MXZYuScTIFlmiki7An/oX+/XA/f44J
oMwftFMLVUKo9ejA7/vomczFMM7L4d8vqqXQUBrBeqEKn6lYHDOH5UB6M3hmG1ki
LexcumbHinbDsilPSjdShJmDl6rRHt2EtYvdSmadZ4Zhqb0ABiPWiREPGOp4AtG1
ExKZ+Effb241VRV8hxrr+LIDBqc2lcYghy6rgzQTxMp5HpfpE5voyoHWbNjfbzCx
JSCvMTm9uJl1fOO1L1hTMVPznOtgaHXiCefdbI0QfupVlkdPrzOi1R8O4qdA97x3
uNqGTmLmZl09BBD2Egv4uzuNhoyMbD6hqNBZ1P189Ft6+E6Dxd2t18T6YiV+8vv0
+3URiuVwJAa4GBWbvyxooI+UDDkg8LbE95tde4ESYxNOn52DIEP60qf1At+l1vb8
f0H52tiDgJuoR/JgjkYyX0g+kKQuopeTUaY9ujum7lenZ+udAoXZctnbVIw0zT5Z
h1TPio3WkKF2XIDaJwCwQxbQqOQ0wVLjJq7uQltvhrXEblxIiei+PtMgwOn3cAOa
ge7ZACpV0db+IoP9pk+CcJyIAjcd2bMNM0dieb3kiJpeH3xMGtRz1jIL3/HG0Ora
MaY9KtlA9SVElsvsibiO8U8KKOEqtKiqDtkq/4ek3gKLpPZVZZFkt7AvGs57J3yv
gYL+55mUyPN8l3orpckoBGE2lcLqcaIgKpk0U8MVmGQq5s7Q8Dn67jWAKMBi5Aa2
PsDIKBJu4ClRYhGLmHfY1IYCG+OXfhVjuGiv+dSFKQLrS/wwajv10bBrPKEvnJdA
Z8eI4u9Gj+7fX3cO9qzz3578vLtMurKO/2wleVa9IVZMn+0QPRBgbIwBXXS83Cqy
e4C/BW3bykKQ5DTxv9UuqVts7XHCRh41E5KHeqflFEXWrtXYNFKoT+h/qbAnOzQB
igirNfCBj/K4AJ6SzL0Khbq0ted/YXxpKR+HwdIuTMqIZ5llsm1790lEiu2b+nRA
u7qiXGMADisGvwtfWJeZ9USICLGpJHvK8w5o/geeSqP/wuV3HFvU0vswvCLcjrJP
bJOr53oLIhAiumgI9so5RHz0QT52bcsAmgcYoBPJzimnNBJPvk0KoySVtVkf2nbt
nm6dr7KiAT4+ZB7235I0HgYz+7Fl0NFZWgOeBcNyIYjbe+qn3hTOkjf6hTdPr/W+
eMoMnHSe0XG9nlLo3gV/cbOjvEF9r9+FUJJbw8Ke2d+QbaunUCwwKRIvuivy1WAg
BbiFOJETrIktk0Bm6/28HOrteKXdCfV/YZMJ5Bab7zF+YAnVfhdIahpXfHpHihQI
yQ2ZYaiTpLwuvY+pZeE+mrx6EeTankOK3jwOq35Hz+u2OfPka9JTBg5EqA6jNIvk
oTp8EvVo942GEGiwC2v5FKoJ6cw7k3An9ArFR1dBJA/fgrOOG1r+tWR/N5jRLmEw
mk2ioVb6ov+O4kXNpeKsCZ0BwR2frONSX2g+nuS2Tf5DCKjYgWjlOnp9OMXnTL+f
Vqe67N+MROv6HaC3tEZJBhB/lQqmTyvxcJ7p2bOFpi7r4tJlXpiEgcpScMdcD+Pd
sm0vabFOB6JNxp3i3blmo9xPhShdYiEvwQc3sc8iCRHWtJDifiHzMw+rjIczvGfU
wDKYjZ5U2gxlIxyaudXZpmEBcLgQ1lRvjrgSdCOasuu5K58eMABozW7G8j1g3FB3
P8j8jjHXESX1LsyHFb5e3is7+wKy4SR6nj8NZfWaIS5U+B1IGilR8TL0d7/4Pifw
T/p2F6KjBdCOosvvVjsbxYWMu/mgozlMbsh2FImfvwl6HKPdj9C2vCopZMvrghQC
37VSHgnHfMFAVDQZN7xtB9W5mcOZ4it7oz6TNJa/DOpR5QsiWTHe3y+vdnl1fbKf
t6mOYV71CnqKRpbkd+XDPCT8V5H38HBox/w1NLOl86xZmPC0S4qXVPK82tVUhG/0
HM19w/Ccy8o8uHE09r3Nsy3oTnROKGALjI6MT294m6FsbYOrDr97GyzwM4YDyNfo
1QwuIYxN77gw+or5a51TXB878JjMEpDf13utIAtbMv7UMbM1drQ3KLDtNCOTn7HI
ipSN5yrXtCZbY4J36LAxv35XYKIOmpPOl6KwQre+D6Zbb61bnwu+qmJSnBtL7pqb
18c6Xpddp0aePvUH6v0RaZTGjjFNbeMgsAvfwVCrUtjyo4amgbcPsVT09CCzBElS
VZae02cFjtcPCkQcfhIEZBgWc48SbwlIS3UAkDJBJNiVBHbWOECiwo4coNsVosew
JS9hG/4bUQu90UIroRsWnSIe4N3ndKDKqbMO8K5t7OEdfkroGRqFcqUuh1AjzVxs
gFrcndI2cXcKjKmAq+SRXonHEZ+VCoOtlaE0WN8Sc/4E89Ykfp3o9qMJ/0Au4CjO
JN6rvc9XGQh+XmxswE2FS2iqWVOUcSXcf3tp3/J74bm16j5Tanqkc75+JBzFbi0J
UC6iDWO91arpkicvCfFmyiAF7G+Zx4OezbFSQ8T7dtuMQls+aLV4wiWPUB8PSfgq
n62okaZbkhJqKgee/STzmFX6y7eXL6QDO8BKHkAoJDIeL4FtCFhRFnFw+PF4pOTa
prUQuM6nB22lGr2Oro8pWlupk5IlmN/MTkpMUZKUfvp7gTCK16osWXyOxqT19oTG
SeKP/y9xk6KCxNZEudLuRNYB+Gg8xv/007CWM/Xgt1TRTvHW8A0PNhvux6rcSw6r
Ux0ZZAgmRZLgl8dxVZx5vAcCkoRCIJ+xfIc0Ns423juQxfZBcLEVUU2aCUZ3s0kH
2m8zgcCzLc+C0T8OJWFVey9y3Snm2aRSaQMACStZu7LQKxXd5X5BFXod4JYxb4Co
f1vysOO20VIzr8HSf6KJLh5iAkW5yCBwSg4WjRWpYiBq94qj+4lRLFL6hIKXwjK6
SXp4MYbX/l0TvGj/pcQ0THJT/3TKkMRgTwShrqVsdc6p41LABNpCFJdgj9oepsaO
Nue6Tnf0+NAXxrbE60tvi4WPnxzjnDoGL1GOyn4LFzS5lVz515BgzFmiXhQX/tYT
b3wvCcqTr5AWBBlKlrG6a8c4xtTKSrni2PZsPboRcCfZHYTM2OYOd/MhGU8iXLY5
tqg374mUM/XGJoGn5HsMTlvnIJdiiEj4f86eeYawhMkY0RCUMFjfxEnYTBNcNyOq
q202RnP0XNqCsnvzHX5N3v9aQlufyhTfmwxF/Ngy/V1aIe+//RDfkkqnZ2l+dMYl
SqJhhDEYf2BmgU8Zuk0MEO7F84mrcL7cT6RuRJrKVgBkIUpimdIM4CRFj/aWInai
NpAhKnIxgA5m1pw8HSMpxzrljXl+FS44SVYli9jrLqrt23klIboQlzGy1iUdVnC0
vO/yBwwMTzX4QKEyEq76aFwAu9+jPmUUSvtwR/JKTTbHY/hGQFRSsoe5CpMdIRe5
+tdCzofsRlO9oiNcIo1SaDHjB0DO/9C4bHOrtYzZIr5G7wIPSwF2+zAEP0pAYIU+
6pKLs9byN5GZhAZg5FuXbeI0hDjHN95wzZ4ehmeAcyIGPzPdyTBbhhi0f7eewGvj
ycMccqJ88FFp5zanBNluIRCkB5ZnP8Ri0JVwf+3hoPJyseIlxp5e3vPBckAUVX6q
C4LrNyudk46z/z7ygs7TI05PztHOruMtzELZIMqD80V9co6/jo+zhTdmlmo6XdDM
MLOyiN1XEWRKfHICgaFxE88bawUxfs8YLpB5YnRw8MNzJ2ZRdT8pK4WxtoWc7Uu5
TjtviTS818eRuGfBFQYcAnwIE2RzdZHuN2V9LNJyQ9WNysaYJmv8WTxuFP2h37kL
mDvL4g8Auj1Xtixc9ePIxj9iiS3QVaJGNTaQDis8HRZlBgQgg/1d1xu5hi+PHkBb
A+OmPF90W3kc0QOmr7eyjmLj4SjS0hllUZS7hqLYPt28YYQfbCruQRVIwqpC+ACo
/askAFkzkAeBdWbW8MZxQlSburCERkzx8uelABiKhxs4c5eohzPeONzLIYkj7Q5q
grMfoTDdAWVslJ8uicClG2hmjZPaUeysLU1873X/7JNG2etL2KOkxZ5OP5VPDBbT
NOw8JXKlVWqs8rp2TLcyysKwhUNIoeclJNF/EwfxLr/VIK1q0cdkWqx/3CFr2W1X
C/sPTtOUd89n7RCRbBkOqngzhEv5ae3I/RFaurRnWYF9Y7LGMwP4fhjWte/B6UvN
+fJpFrALd/bPH/tuH0q9ih+vYWCWhbRW/0t5pxfgxt+0FcWddDC7ZJCMU2xcvgj+
YHMy+XRzIXpSgfQ6ko2ZU3xO4O7KNfuWAtOVzKhVwdc74bDBFMJa7JsU4EWZcsAd
QjCDKVYZyr1XP67BZtMDfr7dBFrLnRpVz8kYtq7IkPoEZZqhvnOTRfXX+iUe9/b/
CuM9C+ydpmvTUqPt9GfgMiFfz49vuo8cRLIUgsO3qHQAhnnTWCPnNS5oA2OaI8Hm
oxT5YcnKFtmTKgd3H8bGtCf+dYb1BRP4d6HfbG7m0tvBIzuoVFpNBC7DnqtTp+88
8JYqlqw2+9lYBuTCccmAcSliJEHlMr1l8Ou/2m7nf+LpXsLUfg1Fe5gL5O4jEOEQ
Cse3UfAPd+sy/j2RhopIWco036XU14ixe7dSDBtKqfuEx9OVCTZYzcWbxYlDDlzm
iWis1eWn1Kv9sA/yYJLuz9MNh7fB+MKXVVhR+yZMCw2NFMvbNrj3Y7tnzZLIS17V
yHKOzAnzRR6rM4DXLm5uaVa+owOdv9oXj0q+NRMlqBuHgsq+nNS3ZRFYLqYeoDho
ZsePPVE1NJ2YtrUk1m7OcH/AJo/akgK+19m3UuhaKV3EGlrzxo2v4Xa9K3Ki05bN
Zz4K5CGnHH9zmmgFnv1JO/4QXvvD7yqXL2tJt/0Rs1tCzEm8xSRu16jWT4MhwMAH
/0nkMRHeHXmr/TODhcW0kUreD7nJ1yTEjOrFGBzwK77t5PGTrrxbkmFORAPVRKMs
7ZYwxyyKR9z5gu8fgn35lWlHpDmUId01fcuZjWiStyjW38ZwNtyqUJoZ3z7aND72
HLNta92yELdgjWzP3vmY9IVs6kK0fcs0uklnFElIdnd3EOhUizQ30vRktxzl7Ui9
fDYYiRdPn/YUXInZ6ubqxuJ654xQHLL+7Wyp5dhCcDmaimJrjsAXaTvTnrvROKEJ
0RalBYB5LVucG6M0m5+TPpvAxv0Wn4+/9MZ/gkoV3VA3oS7Fo1ureCBvtIr9WIRq
+XOtZz/OOXifw2VSoz6KVvIAbd7OqRlXii0Cd5+grOtJQZ71LV9YL/rO7uSBK8+J
GJ+syKYs9TlktA4D1qeHVJ7z5r3Oyde+W92kMjPnG6Ywc7Jte+0x0DksC/XxuGSP
Llxn57nfmNyJZlmsjDGfqP9AwdJxQ5Q88P33A7lyYNKtRP1MvM7A1vKlTyK8iuoO
q2LmFBWF/0V82eAvkKCwrwQMW8AYGSbGQd081SHoOQbvVXQHMQZ7Z9obQexvwQ7o
fSLOuwQg58gMikLxeHy2guEoZVVvnZ+FXCPtbWXQUHgv8WgSXXgYgRmIzsjBC7fF
gEMlo03CAnjgrM5SgZlG1Emg8svhv3IUQ5MaaBEePNg+QrEP0K8DIRG0JhbGKDCd
G9Ctl9rTe1zslT+TXG380wjJ1wFtWl8zuNoT472ShrdqoLiB59R8dj/4eWWUu9lp
szw9xw+FJtTjPYeqfO/eEOMrt1tiMgMo/iYdAXLMHf9B+BGGOUhfNLJTXGzFoa35
/EW/lXjSFIGpki0GnqOcFivuLaLGO97cHnIEqF589ycXxyUzSu4zzbEOI0oRYMcW
V/w0r5BhT9dB/M0ubW1tV87ZEqJijlk+Cx5M8qmpzLG6VIgNcyNbjhR3hYiW7qBO
Hd70NUY+YjqRbS3pgZ2GlFFpuaTL3VqGEZDrcnAr7y4EVcmLjpiL5RrxVNGYE+0+
OgN4iw2ZPtz/c/vU+TH8jBpqndtS9y/F8XnyIyNCamB3YycLu0X0pcqv0w5XlLlM
RjrthGJGIgW1T4B6qBQfvnTOVbp8xNZ7kUrHHELtQlhTwsyoYvYZvLHh0CgReFc2
MwRQijzmW4A6kI1Khbwhi+o9aAWOf61z3wrzTlr6XMoMgLwrNbBzhQ1r1i/t5IlW
5bgxMhcudJO1hR5O6WGQ05OjFDzohZcnM8dzwgOl6/fT56e7tOQ/JviaPn0oSsgR
P5kEzE8G0C7VGckfAjluxNjjZcymJfFsOI31O1UAvfVGlKD+kRgQ859drd7qFHaO
z0VvaWYgicy/7cT3IN0zwSxyDDVblAJgeateItm2jJV5u+TeaezRV5ysCN0FSmGJ
5fLPzPe6Ta1u2USV/7jQxseZ/MDH4+a1taA1EfDlTwweh10eTFqPBX+LlRSt93QL
ETAAZqCvYD96zyOT+Z5cfrA6HQaLutt+AgZ2Nh16rxxtMB0HJ4CxUPhpRqiaCylY
7fNgPi0i1S5gWMZRFdPk0WdhUVddS3OgdeaVdVjnJWzSfG/u08gggzyqeCxd1lT9
OWvMO923/RSam2YeJSv6kN+jrw5nlnyrukq4OYKyFqnLlH5tl50IcWbAEcMUNYtr
6StwW3IQnHX/6lE7iXtQz/5dqIKQBATnE2EPWivZdtM0kDIG/dtmpSBqgxi1kok9
b+S6NA6c909/ve14U9H4cNkJJZ4CBu1cor5fhpZCErP7+0e+M8XmRLpGO0vvTXEF
HASawmfnQah3kzCBX6ehKBcWkw4L1Z+5HF/V+ICOMduCI8FhCJRn2E4g9SR3WuX8
MQh8BFGIHUVryGM0Pmj8DDuWz0hKKhinRHq/0E1RIBlm5cQEOlx6D1vXT0ff9RD6
Jm3ZiUJiQgV1InKOFag0myr7fgKwQPaPW1TERYWL8OKai+RgRw22olAd4ffnRnrf
i20V4dg9g70lzNWFNWi4bhkEVdTlm/WzPmGXPMUphny+dblsYH9vWlLYgVBI1fny
ygAajmovSYoGNCug5g+iUpry1AJJSlCvKUVt9YWKDXZr0NCJoxm1tgI3i9CqjedM
TnrAdttWQ9oEj4w3RTtOmv+1cqJFEt9wrKIo8UTRTBpWamuw+3pcqPfjrbt5e5Gn
mrVSF4jAA77+tEnYC4yVCCTpi8Ne9zQ/khVH6czZea3JY2pu59jwDdRZnC7ty1Co
gst2JFWYtwOYEbozorRHEnGM0kF4RZ/ImkTRv0No2Yq3l1PElj+YUQ6BG00tcOKq
2XPwg5wi0FIlogZ8U/YNlNZM3jXlBCI+PyCOrg3d/EUf6hyYcEL5zhVUprySVsbk
XTqy0PqfYzdwdIR0pdpnPqWatAENkG2w4r8DTNtojCsYemrVhT9x1+JmWnfV1GZY
2xc7GB4Tp8QgWDCB1SsRgcqO5DjKxjZ++3SKlEqTKgQ9NW6HllHfAm3qkrCx/DjE
i5ewVbUo9YrcPt72SDfdXnJi4TcH27DTULqxg1/GZxUIhhZB/HwcjhrOWZ8iDFEt
U3oBHi7iWFV2dDY7776sAEgfIW7s2ie0z/ZS7qHQvhFAUsSjoeZjsIGR7mg/hOD7
ZJGNUmd5Ly+gwbgZ0Pp8EQSdpOPasfbJdovoiBlDEq8mQkJU4FTkZN9PopNpLvas
+MZoAHCZtmdB3BUYRv4sGgeiKy19llSXBsJnDCqFhy6USLBvjj3SjSt1bgYM9Tl0
iiHH96asHDbWhWrGlAFoTSo83xOnbhY3sS+7iVE1KGQdwmJvE0+8lCCUrQMsPf1L
7PA82fNrIpzPIW3e2W8/7azbN0XAxTZZueF6ujCyKq4amloJXz9IaEf+oaUm5pPP
vOvy5JOTcRvErXsVwlndPz2YeFxbfghx2KKIpiVnScBN+w/vE5NhFYbLRmRIEyQ1
pZLJKkni0uU+lEy27BuVJtjAFEgILAdza6fXgO85ByR6OEl1dqj9uTJVtMcCV7Q4
gSimORn2cWXUG1bU7ZZVxJqscMx5FpDrw4XcuRZmhOVr5XE+4VfDMQcPXXTVKd4z
tM2DxqpXf72xOyjRXXDWg358YchyGl9/zTlJ9al+6/MaiW6jr0gOoQt2X6XmMbvj
bm61sUmzfVTmi8+g8YBcoFNlYlmOrfBddxPp6eaB03/lXNSlxl/aSXYErEtX/WuW
5cFHZ9UPnt8kQnFuBqzf4cqzbdjWQ/dpuxQp0HPyWeg4fnrHbcNdB4oTcNUQBOFm
Rh0gSL2nOZTxl22trr0SPz5k89sgMxU8jT2WVBsQgQbE1S6dK5sswD3JFyhDjWWj
6wbcrCo/ibVVlL9kEAJfV/Rri3+lBmcmsXg15M/skiKP184+LveCJAMHPZDw9KRC
AZ7Y3P8CPHcoqbgL+zpseqMjW8wv0Kms3nrL5aPlwBvEGYhAfvPjR7GKOsNJ5whC
wUTAC9yisDV4e5Yb+KdwdyizG5P6b0C1eCA2tmTPlPsA4fo3T19loZ6RYRbtMDDy
cwdTiCmNvVflTRFWPxfvZOze6B2suGqjy4h0LVJi6K+CEOR2WX8YI/MCzBq+icy6
s8L01coyrm55Sy5OPXKfkmyhb1GZoMU9z6+fjBJI1b+rrztVT43RZQV5RIAIAyUU
o0FZwa8MFMzfgBKxIESt1NAN9BPczbUBGFWdsvSDgvTlPvNriZrWcchRHNo81B9I
M/kwo68HpHmF2jurqskj1tpR2z3de0ovqt2YUJQS4udL0Ebx4ZDdY39AaaEe3EMP
51luyNrsoMJ2zHS2Mdzwy9IejBju6tF9Y0qdqy1tL/Lc3kLUFGL4bLBtgwHL5mqX
8cOBwq9EstnwSbv+JUhfiY8rP7+mKBefH9G92bZyYTlMJDn+DiW7yw1jqhDgKLSH
6TjQfe0plsQw06M5h44i4s6hXeYRZ0UuCudKfWttjcflRYqz3mpWh3z2P2FrEOyF
ZyYC2oefXJLzSH4WROFiSMLREKeDZNFT9uCJqtAtYglJrUv2EIyEUoa+yNXMFYjg
ujZOYMVbGB7NQYVUTjW6PaXRea2JNDSd3TYPBBpYe4Mv24mN/sM02Y1qzhVOR6mb
nMmVjmLt7ZPSf6RWi1+QNvjuAavsjvjtv4FdJx/qYEQSryk+K9aLj//Uz2DBt6JQ
GTo7+HwwsJUFO4DsPjPiNUrAfr9SpsdzD0gUlPaMNGXb9NIBKwd48NdJ5b2iP9kh
4OjsqLIHSChVcCooMmsFovY8wDq+6kEiPVeWVhVZk/LfOo4veRsEELdhTUdkEUHi
bm04NujuhodVtCruXOnTbghfmWdPHR/eHsCS385qXVq/ASDmzbMP0Mcxf5FE5eTg
4/vNy21L+O1NMlTUUzlUnmWmwG81Vq1pY3kcdGnEtguZm9W6uPhDwkVrYkS/DoPj
IX2ie60YmHU54C44LLfbUmAvLKZnPw5Y+mzfrByWNKjV9gJ2gNxMNaX0+K9p4+P6
iY6PKXTRVMS2cswC4KSxmaZaHFPE2jko7YByK0xfSmfzKzlhT1WUkhY1edSds4Qm
9WbcmlBPuJZD2x6GxhdBlXi2XKmDT488od+c4mMaf2GtrC6P+tkuftZ+rcLszY8y
A0rQWnFDFF8C1n7181803jrQ1zBrGtFnxN5lr+fJ1NSKmfPGDtTwb1jsk+rKXS11
eFfCITvqxGQf2u0DE6qyJNrcsYNdcWqnGpbunN1ERX4U8j0zS2n3ey50uV+csyAf
ddkqIqft7oYIGY2vUQ8fcgrPo99uVF7ugJS0wv7QpSShb9+Hcodyx8uXbxEvtI+V
2D5PQTZghbS/cPnTk5IDY+i+xdtfGaoRkl7NTOVhrN5NCVm5Jb7E3obm41FRCA2F
1pM7EWRtYtf2hmTKRMCJuTxhGdGXnfTtP0nJRSW7DGX9VzqMd5b4HqQ7JR4UHUTk
huaKA7ixA5xf1WfDV3SodjPRFl/KVbrhvauyGdnlVAbLRAi7252GWTZ3Q6WfYwmV
84mleiO09KKdiAoYpxw8KBurWXTnoOz668Z/LvtyvzTIkYoCu/bn7Nqxa7Ioz8qS
OFywNcWumduWyQlapjnQt6Im44H8+EsBXZ5lJ7YC7G++ONRdO6pwT5UEsvRtqhRh
7j8DHtTgBhdnhZ/V4JWNA0wuhwQ6GkJ2+Ym8PfGKTDaBzPByN0+uvZGzuHaHDNjG
ZzAW6RqL/SCuCgzkn3Vm8GwoWixds+8UkEpmHTNY5k+QJdNKj/7qe3fAXS48DE19
Cziv1HeMTd+jf56W+WnyPmCuWRrxVkSc5NqqPdZTMPx7B+bpOhfToeg6UZiYmieK
YZQfOv6ikQcXrbETr78Dj1honrsA+X+ldI7GvSiaP0vHysjZDDDtUim3a4wsy6p9
JAGRTiCSC0FVAfB+ecJ1/FLWl9SYKSn+cU5YDHFCS8DNhHpMt1SCDwNwMl58TCe9
cEOP62nJbg7ZIVhGscYO0OQXhDWtCQWj//Ih57nKs6iL2SUze6ju5qzLnvUfbijq
KEW8q98NOY/O3NtSL35s5P3+BSEuQ848iWGiEXGrRE0X38rmIt9xkZHcrRFsx6e3
Cx/oCKHN7vBTl6krDQUMdfsrsDQ1rMhwuxWUqMi0hW+kLkpR7oOT1RZKPIMvPgWp
hVFAWJWIdhaVjKJW7l7InLZcPMzCL1OJTUgseCALqUEJ2PcLqT9VMuEZrfk4i3dK
LmIAL3RhUGgATjy6yx3mMQN+3dsW6trQRAIJWPebTiN/XiGb9ilGo9VxDBI8WYO9
/zf9/9SNFcW/fFkl7Va9ys1sHfX0tVW7DpiPkn29J7ondvx/qYNNh7mF+wIZZTJz
fTQrl4rr9SJaAtT6KIXXHKsyFldI0EW7HHtSSkS/09+/EhDwj5lIhpwyypwSasi2
5NkOizMWhZmX+SIdekBLS7q6Sf06qjvzyzVZxBxC4YGkNuIxdaFulPxNeBiFlnTA
T1zd+QY5keQRzd9ikv39zdC8bOLuNkQmDhCnNTIfGj39wWFxcKn7IgXpLLKglK8S
ydlMFzLl4uoEIKXUeuKw6fZ2yQBXImnvOb5pMwwEWugUNjKglRZXY2Rqz7X5ueQQ
5U2PpVl3q0PVOnhMhhCK7Lc9pkeiptlNwGvi49p4EYHJxD0R/9/D5ccAH24zp3K7
VCersP1Uh4dy8c/i8/EXfVLqjU2e5/MpP821bgUNvMwFvOk2HVgmAbw79rwYb30J
/JPs6vqtuiMFEYCUvbq3YQq2RNJHpysXDvcv7l0pmLk06JGqpunwcqJTePWdhwjN
t1FER/Hqzpo+yoajx6FPe1xPDomkQdimZgG6LwKrqa2d5C2OyRhcpBZGgHY6v9/1
spFluSb8halB+c5xNNg+GB2+Pc3cXVjgkWkosUF6x7wD7cFqJwwH4Fd2xY+MbDuA
dYDPfx66fZBSythHc0SU85EiLy40CA45bst9nbWcdMP4zP162eMuSWkF9C26NVGF
9e8w3016SaSEXRCygHOaFIlYAjimQGhk3yG4esxRIPiXgwz3bF/wX683zqIA+BT7
PjmtkYlZGAYBRJIniBsAapxkP+5f6/CcD2RcHaBRnDzK5caba7VnDEF5Qyt6jUKx
536sdkVgha/Hc6yQ4UGZjl7gzlXIO8SfVU+cbTSIOr98za7JzBrDyAJa6aTy60vq
6PjYr/bsEw/95MOFm3TpQ1g5BNtYDCb02MNp7VjJM7zFI/p4hJkM3H/5OX/Y2Lbx
xADawPtWArI3p1XSPSxlAzc85zmsABIBehsefYA1hG3HH9kze1VlR1/rKxl2j1Y4
wixvk/pyrsP31wIZw7H3wnEEYcTQtc9FfVkKFlD7U7fXLKy5MJMMRJjdP2+TVce4
KkSA/0TayXXyxEvrWx2DUw7T/KBPVZPrsqPBFrnUiJijpzz2n9Eer11/1o6g6ozv
Bz+2isck0Psfzwei51vtcQXe+LgZNu0skNu9SXoF648oylpHlaJUuj02hqwvjmNt
ar9QTNtNsOhzHs2pEi8Z5GKZbVyCKcI7x8jMUPfWP+O6x9cvpiqvHGF2wQOoYTiJ
WiDPgxhN58Nq5weaBlabtdYi8Xn1nhxgenTuaXwN9i/L0p61SBpXtuT69o3EU5XO
WNEMTm6NDCw+3/VN6CTJc4VnS5gRRvwWTp7CJwG3XWj2qt7xcP5EmovS5lHy7mYF
esbzno1zv5zygk2jdCMSULwBcn+zZKNKkKw/gqzQ+CJStYVuFht3Iahilu8rAOpV
duumP/OkOHDffGgOHjXj2q0YmuK+kGru7jmMD8R8ZsxEBk9KYDeTkp7zIWGECjWx
PxEib3XUg8sIBbnkGTQDGBfFPT3NTSiN/o722aOsgThmuGtrLkVdasiDdJxmCGk7
64ZLddn8VtgTcHPU0MiPsJALChG3eGelHAIdl6vbJwViAyy5t/lUMaXFkV36HWwD
Ezdwhs2Hks3/XE8Dz06Jfz8AayR1DN4woFX5i7lJ6tQSaqtBhKaGSX7z4vkRRI8T
Ixv/ucezjEx9vkpYg11NgIvjIhZCk8txqeNd6p0mmLmvLFBC2hl6SvOcicbVMTZD
HR+zhbMC2fZ7yM4L+AeNgZz6aPfO2YxhYNea4uVwtb9boppB9oR83SkE5ueqWGOp
KTKiUqn+s8gI8tgjCIWxKaQrpeorc91/44IlUNcLfZbGx5o/Uov/IXrWZbEK+eEu
SYE56vqPNLeOeH8nLXj1vI8oaaS9MQgpXZLydmHvIxzYAcFExXdtGbkHBayaPsGO
IPd/bX6Y9q7E8nx2GCVrLhhDGONx9jTpP1cM2r9xy8WLyJLmzWa9NjbYNrvGr6h7
dK6cJVpZC+O9HrsriWEhmywpZjSdQD1VnebF6RGluDq1r/HzJTw7z39FKcOY65ur
8MdXCL6rUkniQHZswH+ly78GIWvDqKc9bxoc2B3xTBhOTrrAnKL8ynuzQCgYJoWc
971CFdz0cJ2S5uhqpg89hhnb0M50c2wNhPLf6pqL3WmaskB8bsxXq2703YwHR7/9
iVyJUE/C1RBTkdDL095vAkGritnhnhyUH3FIy0eVVIQG+kfmyZAONXXRIVgsLe6B
Eo2XNRiWl4A9pZx4Uroo3MSDIyPnzHMq2QEB9mXYj35tF93aXlSJYNBKw7a1ybgA
6KIVaSH1pC4b5HAVRN0c4GYivMXJI8oWS0382frX2y3IihMzrZfQVz9+CL+txwL1
z+QzjnG5jaXONFvB93o2BQ/r4DjS2N4Fqvzz2xo1yDuLQwLe6T4SW9k806dggjDb
g/tQmv5gPor/Tg5fR9dW3bjqbT+Rsft18WAvGDnBSIWL0zWRy+jpUZTDg+ZpSms4
fEcdli0/ypeNN7ukqK3NtQiPZ0zDD1KiJlr/8JgBJjeYg69USSaIKEAkE8ZHM+t+
tOOsl1gf42MpKnRcxvFtQG+h6CHIMSbc4OIYcX8wvQob5EEIfK0kk9nrVyT+rbrC
CaCFWdv+wPxizhL5hCz5jvZBtIJdp0rghgA0x4w2gCLRF+R3q/TZMRFeZfeNx5yo
/lHljhz+EigzOAi6PBmClWv8XCjXfFRijiMTsX1vznLmW3CR8l2SiNny5DyLuApy
vDRf42QdpsurPjsU/irug7o8jAoDD5D+h8Lx0J3PdobV9E+DSZrZaTRiznMKFuHJ
h6M07keU/pWi/aQmGKYLpNgjz/NL0TiiIoGBoIoWJOWsFW1LrA498GPzcOA+6USk
6Ag+VLI7OgjzX8AXkhBFwKmwqUX0PG0yJU0t8UoeG2Abe/uf5ifpYJmlTFoAvVar
PtAvB1f+eB6g+bqYN5Tz5VTMw9x/gTqtQHYmcYNgZKh/Bb5E2tMalQ9xDdTw/In2
sPhTu37wOhKHTsnTuC9zpSFMEI7O1fFLqMMHoAW3esxzRiPLClfHrx0HAC4uaqyk
EXSmUwFUWeY+HF9QJUyI2mS/5jJXOzpWgh5Aqrrzoy4tG1MvJgT+2vb5Fl+JdrRh
DOSAxc7nR6H/4vB29Y3ohokjAOi6hSZR3vvGA8YLgrP3C1sbh6BF6YWp2TCgNNIa
ZrmXjUETlYcBujQpw0GR9QwpMRgB0u5KHIMERG822drT7cFhwWzOJR8ib8qn7GFu
uli0AHiu8VWQibB2qmE0dOX99HPAjpgP0Uind9ZOxMKkiPFsUaJQrY7LuqkHFRh0
w2xiY9pt7hcsCeFrswHQToCj0Z/+FiNamjG5dmyJu2gLQM7jG6FzRwB27NG6dAog
znzT8/cMlwcRbQNFQ9IFULS173IfUu+CqJlNbnMF2DCmxMFxhvQSpeuI9BTOhTfc
5hxiIssBjOXU6ZJzFl4p1pyqClk2bNGMSxbpBBz5yz79BcavaD61bEjbZr09Q6vY
wkbPCmZI8DQ92OtzglbgG+nuibOAeMlA65x6vDGB0BouscDiTxZGfboMRB9Syp7U
27ZYRoXORKpumh9RLW9LfnjfrwQTssXHppycBJOmmA9deezUeXGcsyJCpTkfDqN2
gcPMRBkOfEBOwSKB0Jv0Jd4TYdNJGwnwsbOSw5siqbM7U7VuO8ZlrvrhoMXaSykp
I8MlIgFtL/qk/8swVpB1rzQaL3dzb+NZnz48X2G8c+7K9y04SZaLDhCRGUYwjNoX
v9tosAPGZngpcmfew7BI40cfuBusHlpyZ2OiJ6vDcJcNREEfjzXZBLSfhTxT2vDG
NKHkBrATQXW/f+DSgdDsPGNMXul6AzbaFXu3+Tp74aeCaJkASzlCsA0ppis/myN7
a9Y6U2MqTY4nosF8N2kD4NGYtZqcCSyMDhpuaHL6hVTacvr+zLbMQ8YPZ+duwClK
F9NEOu6cGNBGTQV4PoRBUJmd/wnL36xUn1Gyw9/rFKNyOo0BmSF9GmZd6hh0H3nn
3MVCpxw8SlOERz1EKhYgw0mZMA6t4ruxS7SrsfRVOmahX/P9bYqMSggxUNNMHFx3
jx87pUD2CYyTsVuHNm7iXsYw2ARmgkzory+G4DNQx4Lf/+EQJLdS66506Anb7H6c
Po2EL1cJttbWWC5PvhMp9d2GXYOCRFjH+NIBvzDaytMAX1DygE3d9EsXjona0huj
3KbukUt8/LrvGHEbsl1E4me1tWvRd1QGs0uhCy2gvwY6uHR6Jx0/qP69v66EtF1W
adRv8wpFmv+PTlaKOAD8kCKYWJf+riGdBZu5MpEbUsaJxl7YDYcpDKWv5tt1v8+P
U+b/20Ky0Izu4c5KjSGgh9H0SM1xse2EAZggUk8dGiUoz/m1ry/MsGXMoGqaBRLO
G/SMMWL65ryAp2D9qS8lf/cZw5OvBpsRr+8SUiEzro9bwBwKuK0ag2c/nBcEO0zT
d2MytNh2IK4US6oe4MNkCmabsNzfJlylGcDTvpaK1+vjYGuHJCMpSztvYneN7cug
w55G2PCkDYSQnikxE1g3gfwez4K88/f/QSjHKEhosSMYVLPgHXSK0oyq4sWysW35
41o0Y0j1E+2apUUUyLhR98T0rhEetZ/X+fBhoOzFGYEyN90mCehxgUs4JfUp+f46
riMnEUa+Dw6idlb1EyDseroubydKy5Jhm7rx8A64yt4L54CwyzlwkRw5biqPQTRE
HHoAK6Zg1kkfXsIqfrlM419kN1+3g10buvoi4ZIu4X97cEf998Su4P29+w00F+tU
vTm962j7hz63kbYiB6Va5WR/8Ay9MHEzFmlk9GFMgk6pyVwv6yKJ9h/Vvh34nivk
6fxTyESWpRRtgDySBflAtaNXMJ3poGNoZMDPL6p+AJZlFFgHWTGLos/HeVr09CAL
9ZKWl/qH8pc/IxrXg9SwAicKnIM0fybB58pYpFOL97BmC5GBGIEPzHA73hLeWcfP
cntJHrCqMo27V0RyKebPLTNmEjjI/IE9R+m3xezmahs3C1N/lwAc7ipH9LVdflWT
zi6mGxDT7xqJ34Vw8qNtSaSdyGhXWyZ+09S/n5LcGn7f/rz1smWt/K9iXkCJOaSK
Pp8W84NfwL+W6Tj1tUxfebgH4q+qD/FbWxY9d5tiVQYqDQaNaSkJcJ5RCGyk2ZiK
s+9SiD0CitHWZFgSowFoENHJdvlIpXc9DP+OXiicJPp+ICJbSFZZR1SOB1OWihXs
NnF1mNri/SIBZ6wu+ednQTrUaLf+1Fe6Rf+5dysx8b5iHl/MFmMkrQlwG/KWn0mZ
3aVOtCyGlR0NjBm1EzHgNphw0lhUrBLNpKaDFvdHr0afkfLUbwAa/03RAeksSc6v
P0mN2Yscm4Gs4NcqnbHrrSo+pn79N3Ahf67wOvNmNggoTYN8UA1xCuBnbEmcDkCc
FhIzd8rV+Nu4CARtsnEtcoVGBZ8TpQhM+vTxn5FBR+soDcXkgm8pcfvuNByJG3hh
mKuByz3wGPDZAYBJUjs9b2qJk0CdMZe+QDGNdRS/XXk5IOWQTHJ4JTWoBUQuX/qv
n2agEwUPuCXEIkyPJEYb0/rGK6D4B5vUzDRuRIDCpWwYb/yCNOubOf1vrOqsgszH
3ZvZ7Jjdrh444NYC5XAEHC8JHe/bxxPO3dQCvQRllVM6DhBMDUvr05lfjR4Tydad
LtvsVdi/QDdV4UwhDE3gASxi/3AeVlndb7gGZEm+cHRovhknUjZv5ciQFNNQR0h0
dzNT5rEh3/bk42xrHnNfW94j7cev2RvbtJV/bfBPVCzRWXZkP99H7O+6PhFNgaLC
L0yQ3Zh0LynpOqNaYZ4v2Kg97grPpWqBQUAuXb/g8y+vvkKD9GugFwCVfJAj8fy6
ePgF+TdK7p4CDqeHjc41W3ICxhz2lpd8ujqoIVGH06cYpn26AVl/fg9hvjLCPVAP
z8UzqtTa/KN9aXX6zzEktdAdhSIXmgpEavryTpcCzP5ikmbdAHVmOQu1CWY2dEhV
Qx60+Dv6u0FHCHjGoKv1l4+uJ27sAWrFxH4qJubAPXnnjaLPGOGUSk6wEwfjIb9W
8uBFuTV1iFlCFda0eyabkzbMfV+bKwCthkusnSbAQT1GGymi9/3sV/J1tIXT93WH
C5gkqdabW9bSDxI9/8XSJxVN2vnR/2b82vEFXLHszVKKbvW8GVyBSVdZmmiCLNql
eLEUt0Uh+h0uyDfnVhE7DRoq+6oNDF4CbeMa/v/gQiNXiY2BREK2vUImOdUQE5+O
Zr/dSbuOYkYC1xhoqd77WJ0bf84aTtza6pLZ3swb0YDo8M5jFxJQINtKXgVTLtKE
K9EJVSK4sqPcDseth6MXRo6NzEGCOoEo7vPWeSt7ZF0nk+k+322DuHTw9uXZ8/O2
U1MW8m87px3KImfBPE0nY74Pc00hjWMHIVyjKlN1AfQrei1c7prI6NNQgM7DHs82
44E8KzMPOItW13HHKnWhVRn/9+fwiIM6ndlVQIuLn0pUSCqIZQzybwjEndwLTd9l
GyY32KhwsvF/UkNuBi3eTow0iWGSCJmGfu0E3q8MqhOtPm9nCRyisu8OjK8180qL
BV0AikLD3dARLm3TMfM+2kGk10wfjPXdOmIT/+haGG3aVavhfPcL4tQaVhF3xzc6
Pf5palxQeoXKXUSrBgFwnTnD1YhIrYcWaophEoo9LFokVzI2slRq+gKFZLta4+aT
6+x/1y7ypxl7InVLfsYUChn4NciNNaOWsJu9QbPgMQ2WKuY+zPxAFJaZj+hByg/V
DgLfk2tV6F6R8fk6KJyYYduLedSgIwbJNT9Gh69ZPREMQNAnFLwbfrqdNCZPMBVS
wlatF15ImUKeBPE68WWERt2d6O2yiSg3Jlo0fsdaplT594wq8PrLwUgdQ177cp27
E0nUiGa9gsMXnIPX2ySWhswqDXvH9syl1nYEPTdVcgpvcvl+3pdmG9O9TVjKK+7D
279C4vEqpF4TEVB+/7+yuofW87a4YP5QlKLk6jCh2vxqpr3RXcar91Puo0qaUJbh
Ky6i6Z/4I8mLiKggBBBEozP9fIofGLhveTppQXuL6FRFesXIF4n5Q4iE7x0ItSTV
HKkhwOIWmP+rPKJnw76UTru1huEy54m2BVJ1O39UqaLKUdy1v5TkmuzOyklPda/z
f3f9FS9fodT8C4/TG8pnh461ZALK1b9iraK9MCgQ2xPq1l7k1+cuuULT10z7Waj9
Z8liKZyAI/TP7CHybHw5141XNUT+x3GqQmEt6gXVDGtoOUgzimX37XLHu8pC8KG+
BQ4UEdtJ8HQwdB4vjWIJcHMcFncmWr5tOW9qApmCIAzk2BbZxE4M/FrKHpKA7afI
MOLoUuLsGRM34mUcFxdfBOHw3Tbe+ERkF/jXOMQTHyrF3zgOopFtOhKl2svVHOtY
tSkJA/5+/f/NYHKaZr+ZB0+DnXRtoQMwtC+20i6+nFadSTXewVTp3e1aOvi8vumz
+55qF2mA/wv4Po4KFprw+VVGIjATn+E+/P8c0KS9NsVicrXf21kRK2xt53ijsR0L
3Zg0U083G5b9BM1K3Ey98uEP/xrpCSJscyFWJkLLnRB4eq6QD/r6c9ZEQeMOJ7mT
fK18lMDDzXdF1MrY6jC7QMoB0oZ5hi9h0bTDeJbBAF7qPqXQIWVatkD8X9sLiD7D
Qui06LMm7HyRLi8hZOh3VUw6Av1bNH7iGKZUcGLUPJJgPzocagiMpGs5LJ34MrMj
gXMW7PV006byYi4FohdEfFQLm6gzhrDJYXKKYee07HsMtcZjSzMOQRY0RYr9T9GP
vZTXlyyWoDy1jjpGf3W3ZE8vKUbohBV4h5bkFjPVxmJnfiPydXWGkbZxlL0So22E
7LKe17ICnp8pZwFpIx+2NYFhmSEo3/Z4PVrbTzSdSYqqP2RhI6uObJr/u6ge5XCy
AQSpVRiIpeMDK5ZbDisCPdZODTOArcCIFVpf54NBQ6B8NdexVwp10AgJpKD9DYv9
U/EHDPQzonWkHOtCgy5UgoVVJI8SA+iXVChLunXKlA9PfmgyPILGxMlNPQFGIGAb
Xud00sCrTJapJwggo5OmQTax7ZpkeyEK5J+Tj1JcGXIwEgl+YS/cyUyDxbIuDu56
VuSCMStWnneHNcqRzcxdon8LjpTyIe20EHXl8kr0449C+XQuWJ3G/GAZBDh27Pp7
HR5ptOgEMn8pP4oAvM63IrsIeZO/rquk/npDvJhIDofasbZ0MtI+NOL7j/wmnhnz
LDJeZ40zY++SYJU+gvVA7Fl2/MoDWfyyv/pKrVtqBg2qcWX+6hZD1JNyy5pczpKI
/7dJDbamxKZj3kjPW9cWrsJ+pQSckGBl/dUPhdhrKHFgZLaW902jJTq6ulfSzXbs
4JdQ+DEZNayQpfgtlqRpwuBT5kUAnzR7ZVcOhYtKPIMZVl8o5wbJnEojI6kJF1s8
Dg+gra7VFabSIQvcGt3hRTN/LBzQcg4JBXZY0VNvAgdpH4mcqsG0A5uSVZbWeMZ+
RqTEBaD+GLWdeC4CC0+yRiyHxggdeclhaJiGPyeH1R7d3320o3ALe/MiiDl7UNht
LRWGL/b5vuf7oEVjLeFtBd6plVgulzWuVVPCYiQMxIhqqcAE5+N49qo9dPKRSvQZ
NFpplnBRRBLVH2HqoSDeEDALsg/0GWUwG9SnMFdZ8omqG13TXO41dvFy+wnhDi6T
S+0p/axZmZPBwUhsL560oE2FPN7zmxa9NgwusCmaSSqjUcVQZjiL/IcnF8/zgFw/
I8EqhB0SSfCzrN+Odfr23cbki0n82Jp/7MoUls7Suc9QZv9c3D2EAGZqMaFip5Gj
XUyuD+Z0SCIigFwMNPshjwHTaKjPNguqHuQlEKWXB2t09+Sr43qpXjnqrAZ/T6HA
ZytQUhcLhZrHgzsvQ0ThZS0H/vi6bqzUyxofrxxdYPm3g9HHIwk0tE1z9XdGcx1R
BcKe0rf0Mm33TSvY1HibBbYd93YSJkHmpyKFYnVzBHhdbyCZr7ia3FCmopQ5VnUA
mx980IauCnXHSUsJtq09ixapTMNpcdspkcZYwUDqwdyRKDFkv2YiUH/AzP2SM5yR
UGZIoiW+hcYSceAMYTsE/D543ywoO568yoxXaAP3mAwRBA+iFxaa4UOm+5kMjz7D
3zGBx/DNcKgRcPb2qGkhSte4M6/NsDQ+8JreRxYDVWE+HL9ROR55ykS6DkdQwzxe
89+YUqEH+DKYtNhJjT3B5kG0Pc7yHtNBJkIPYlvX9oMlaqyyPDsPCnDhbHVkYu04
66LPJlUM1mQUNaPxPJpUGh2HY3cizBOGuWF92zV1nyX4bSWfXmCfEqqF3XE3/8Vv
LSlB9mM0pSYCdRW3ut3m8af7fpMsrZHnqdJHeh38Uk8axmy1BtMw3eIoY2UYGDit
fIDTrL8S731drmJbL+6itbs+t+tSNEI4w8Z7CPiYR4pziKifFUd0fws2g5ybMJM0
YdUcaXEKBxnwRVrK4dpOWAvVPKf9lOR+4qLekO3a40+ZcsQd6F6Uqyfy532eYmOp
VQ3UsvKi7+txczWTcPwKGR9L/Zj2q0tGG3y7l05uGS7DLB0fRJN0h3Pc9EUz4xaO
nJl7sMb2w0mT1x8n1qB2nV/ft4TQaV06sWPI0cVWm8wWvIrz3pWQAo2riBpH03RA
fKYw53+hGMV9HZVs6EQhtIkMdfG1jOVG5z6MTMoNTyHOMMqWnDoWrrK5zYMbdnR5
miJEerZhnhbauUYFGOhRlyTtuo4cdHNd38mBUd+d8hbu0Qc3X0sT4oAFAm23qMYA
6MjVuReSmmULnYtN/1s9gR3isNNzgYixNaFzEN/kgHh7bYERbuwjGNR91y+kQ8y2
0hxE1kvF3LRgJWiEXP8KOAVrKHHvFknY1KeWA/BTrtXGmoha1nNwfipx2SbTe3b6
FF6vm1ZVj/pewLfAJcJ89iCYEd1CdiO147VOggHrS0qUfZvBOi5SkWw7Ndqdhf0Q
ak766oYc4q93XLK7/BvqSvor8p1mGTQVELcdKCVdm/Yw3kE3nEO8ju2VAl0lrBiD
baQam3oitnJ2JdXBNDNMbxmtcuqtZGEMJdycfEc1eYFXIfak6Wx3KT7dTawgaTVt
HiirpZ8ZriO0qHEx0CAkRqXCUHh4EznBrn2cl7rRxd3OkeSvp55otloIYAeGULON
y+B7l3diPiOAGBgYSYPlREYo22YjY2cDzvLkXO+9g+wiI7mn2D1us5eP74XE+qzU
3WXhHjZDFCWfTuS4XbaolrUksAGSDAjriRc5FXml6AOrytf/WfBwMCO5PUnmfIfN
W4Uf0ekvubn158kUzWm70ossnXqEnJUdodhyF+iA1E7/YoBB6cplf6qiP6TVOs22
gVHiuTnhpQbCTXSuTfga35WjuZ2WqwXCs5rDBIImEZPXXrxUYiQiSbKS4aQc6V8j
Sd2Ire6sI+NzW5nCMPDd5Lb+Dv+tfO/IimTO4IdMbdkr7W9JHIVxLUFcZllXc+te
0zKq3QuVV6t8bLRAjPks+qEAZUd5PKyJIwT8rAohm2sag6o544+d0fUBjCn2DvQK
DDOMA+Aqwxl8BQX31YfIjxDCPtovIumgz9mDjPpRid76VSqfAcjN4b3dB9Mi1neT
+hMj8ulunQmv/OX0OowbXiAjItx14LbOc0IId+TC70jmF/ICvULsVxxstw5VI2Bb
6M/Q9re5kcbutn6QL3F0eY1ugDqaScxJaQVkOQRzA/37fP5m0UTPmAJPrU3QgyiX
YL2fHR9QB0AMkUtbmj9Y+475ojI5YPCUWhDsHpWfzU4IWAr+19J7756c8WhJnc+d
kpo+zSfZuS28frKAW1PAZp9QY++h+wNc+jyrx02n3G9iza0Qzj5diHJTGNJW4529
tcKwBo3DjoY7Y+77m+FCymOOqZvbZwSCfA1ePDoTlVDxlpOFpmO1+B3KFNNlKLxc
YTn8EcmTNzD8+a9KT14wmMZkAQjwsR81hClISqXsTLKa6pjo4G138MLaDdWWhKZ/
d7V8SJewAgZ/442rnKJI2CjOz5uDpf73vhMlVMCpO1M37vcMjuL8WU58WTY/upAD
GBVqFb4mjg0oc5bI64+Xq9eug3B6TiOZohJUKCbI/Na1JxXhBgp7bWIcUesl3Vau
+rK93GrAIot0xjgVpkLhfzhh8vBmfpPIN/Pbl+si+lE45un50i+xIOzxmzgS6ASC
MRo2X9oJj0KsJNSBa8NCjVDxtBKkQg0zBxWAZ37KQT8V6SoCDzSnWJZaGFVbNnZH
+MI0QfOAUPPqhz4O9GreIKvNtS/FguuEsD5wakHe3yj95YSjdFRcTSyOsdpvFCx0
TCUf/DNGf4zEPctX3bdPVsXPfeNJt+QH/Z3klHKII6luHNyhsw5N7ZM69cDXJAUg
3nEIEQVLvN5hq+MHdeuQ2nhRynAWT0zGEyrPwa+Ps3VEnw9MTPqvbJA32untJuoK
fGOkj6GR/vbnAC31wojKSyqUwCgeBUhOcy67ieMDl3cn3YLh2ETN088x8ric/6kp
JKRV05G7CPXZKvAGHB769/3utQnEkEnKY7BeER8HmBYaLmrM6USRB/h+BpD0bDYA
cDGhOyaM8NLNEcLMKZpdMP2IF0K4nQfUTzuGUBchvpZANx88QdEWpsLF0mOyi6nq
o5HsJdPlJs92Lz4NIrkRzLUBm4nBcPy5EnEKZsej6os2eBkHWKDhSH//eunhqRjU
Zq+uyZGzluVDMfeynLTI0aIyhAMjqS9xvGDBzwhuqarIEq6UO3KUpIsALf1JLimn
hRUq900HDlB2pFm0jD5e6THIM/TgulVzcQPy4A+JBGBokfvnWjH2b1H61Wps/0IA
kLrecHKUR9X/8IGzCUKrZcJiXFbbe5KTPNS7c9EVwp61wbTMV2nAtq6Ln0J3sQ3m
PiFLOHqbLJ4vvKsZsCHUg+0sxrsb1hW14wPiZimSwIu6KAhRsz4wlfXswFWlA8KW
DAa5GyaOzB/xTGhwYiOYgHbBCyCtp7QqtWe3bcVXkNjIpk6UdrDOHNjeRa+sjXHR
YDEMJ2VgD/Xsc0Hr4uZGW+hctCL8OnbNZJKMwSLI5Bb/ifxtkIZMsns55jiVQItE
GD5FJJX1YUoyQ8vjbJFz4yJtUeazXnw6uXvTHit6vHGaDqFr2BcDvClsaigEK1qR
U9hWRj5cc6mTznvcP4NCJch9QnKnAPZRkE5hhxVodoN3fID4Pk1yWzX+amRoDm8t
SsatNn6cCtnnLPZ7kVtYPSnelDg+k/th9ogh+Wdbw4xCNtH2YiLy1tD4r2wR8RY6
q+pKbZDGmX2diYYZ6j+hHmkRB6v29IqPY07KlojP9BgLP9EwjqObzSyR0IWK5Eib
0r8ngV2TF9YPCZbGQUkGGpfZHnIOCNXg9Q4LebiaTzg1O2C5WOLvViyiDpOuiUZI
v6BUCNkPRoEQAwo9pZRe0DQMwCUs8W0fKW6PRd4BWg4aa1r9D4qq1nVabLztX05U
nUFcJY6Rncql4PQGte2IWs9gK2mUOLT784f7inZxNQtbYqioY5uC69iJMJMip8qq
Dj3oMqhUwOiZbB/FYPK7n5Uf9/Ip870RcegMyPBkmZDVK+MKGZSi9NJpy4g+Qhvm
4FapyEtA1D1wxV3oYpGpMN9K5ZNSMhSFpAkhDZEXC+Sm71qxFntsXDCGBRdilzqT
7cAUmhiupeNeY2gOxy9XeHkNMCHb1qDOPj9zJhQgdYJ65nX1A62xCPaA5hEH07Qx
nl8s7gfJ+4bEz9ufTJGw4nz6saGUWr9aLKxXD0SWqePm4TBlsUEEkCtRl5CPO6G5
QDfrFSzMT50pGiNyu6nEYQeVjK/BsJ912woLg7lJrRAUQEnaHqxA9h7QTe4Hgo3j
8/Z+Y6248rhDfX9nHuYGIXxoX0wlZEbcQjOf/EjWB78YFR1cCHK/MLK+ASnY2yDR
zJy1f1FcMxTaGMnc6ylKGhl4Dtcj1Umm6wupZlW5ZqVb0cxogVN8bgN0H8d0Dw4h
lpbjiqTxs1a7wQRBchMz3BdIiNhizDJDxdSHmwL+sh77pH9/NqUbRsDF5UX0LET3
06XMU1RXZDJoo70JOWuvnahJP0+5/cATrxmZ2LYoEEdSQ+YkQwAfAFN55BlzjvH+
P654uPgoaeR1yY5udd0S+UG4b/xVZa/9rBibtwrdVXeGxK7fLUrTuiZo1smEnynw
J8vue5hAUtpBrPfvGRWNv+8hRaF9tHAhAfz03fLWTz9tQeEV2MGIq07LGEEMGRzb
m/cYh/7wgOcsXYhebXGXW4SEti3e2xdM6yWdUjgu1CNwUzGowwyWyyudgBgDn2/0
rLnz4oMU1vfDOqczdapFFqMO1DlOWJUmyraqzY6pOQ8bTd/fxk3nxsyMsbPFelQ7
3WaHLp8bGoVYvMZJyS5JoFHFrB33GWOKEr753JKEC5SS8iJN23JMAONhmtboBRQ2
jJ9I1Q2f5C5h3xtiGQlf6R6/R6h9mVTfnE4ktu1IAoDF7Isln8ScDX+zhPlmBbPX
Wh77VNz3n5PyTd5uHLz42/k2uw/MJuS2ljgpZkP6CuRam+ugwcrdkKJ7VNPMtbfz
o5DmjbfkaZdNYwpjZLFCWU07+ob1KLuP7PIXzTrqVJ5ibgycQciTmLJNgw0wsf+O
S9ZFztx8IF+ambCdl0oxlteTlJB7FJmTUULMyWY/HLByzSy0UrRjVZeGMDuzA1L/
kK1vtgZop6cPBiJ2pK9eeOimvRBvrNJi5p3DuFuMJgPQTOi3JmB8Vif/f/fwKpeo
UMICbd1WHaT+PDZq4e135WPmpgodXZTacSAhDQ93FMKEf231lroTJ4EXzZroIV12
v4QIU5Xl6QODSJPRTQS1zyi1s7YuNvDtm0lpUUJVOAWhV7Hux2EywlZNOp+GQe/m
eVI59DqcaYuz6YYXbrBdz54WN1D27FShh2YnzPH8FKS1MSEWtBq8ZhY2ZSQp+eAB
959lgCNUr702VxDooNVBrSzbmz0uQujnZOpPQX0LzX8lUowTlmeEraLqFUcqoJ3j
DkfTPLz3FBOrXl8qrZCSj8BCm6ndy2YzEbNHNKtWqkM+grKP0x9LtpOdV4ncfD4U
Ra7nWyIiMrwbzGdJYawmb6nbBbC8d4WlNWXo1LFv6olaif2/FA2ZIMaV1Md4wSIW
uMNXhylxMGbKb5TDyBOcsZmx/7pCWoCABwHtygmHbYDk/aiRv9uzjn2SUAz0i8ii
hFUA3DML2kCCmfy7X/ST1ZRT1fqm5hSH+1rf9d2aEDy+lFs/sWBB+URJaYrrnpAw
T2NFfjmYfkl+KXM3NK61C/j/uiBRjhpaqZUQ8wmlunK2J6c3aellSK0O7tMoP+0E
ZdDS+dCu/4Hc4gwr6aU2L3xVJ5iyR+tC5SjD/qRqaI8XuqF9vvEPS0AYSYgmcqOb
iu3L7jsq1hMYMeTlvc8+EfD/hfni8vXyi3k30gm9dpA4i0LLoL36//j7jZWNslq0
XogNDWtA3oJyREcQn3DGMEMP4oKe0kmcFoO7K5QUC1UNmScwvj4DZJRRqFl+9lnx
oy+u+zWntuAQ2jwDsu7SAXipDpdw8Ax07yHnqQUwi2TzaYbmsV517yv+5V2xvoUh
ikWrUCmIqEcFhEq2tmccikxdoueO9OQYvE64pbHXeeq6DZMnYz7m9aKKF+MPlccI
A7SILM8V2SZXTbPvzGwrVNZ+RvWsDaxJcO6eZe5NvlL2eAm/dZ0e6od0rG9Nv6mn
9eZqwo0LvBd+TkhtFMwvlMMoC1ThN6C2SSQT4FUYlcxoBTL2utG4fZRCQLP1SdFG
masBUJqxekwPxREdL3orh3+pnNZnpA10EZq7i7KlKjuZEPuaut8FUyw0RkDJ6ZpG
4BoR0aQJyQcZ7oBJo37U6oHjxqBvzzoAN3nn1dDx5ac2ca3mljp94s6NTRs32hWo
FFjjfaSKUk/Q/YMeQWmGLa3i5+aQfxbcMeHTDy6Z829QSP2SSPsSYeolYjz8/2wN
kBjcK3vGksloUfnLd/XBj9p5LLEdN0K3Dl26yW2kuZq869soxi02ZwTdLpFLm04i
`protect end_protected