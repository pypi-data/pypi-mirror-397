`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
ys0fr3rzP3RAlV5qetsYN1o2G1RlLzFAxlspN2cavb+csfs07F5WnRTNm5poKQe9
MpCQLEoRHHGUEFz8H8J6rgpL5aLkFA4KkR8mK8TuOtRwgxVrsV5GmvOkt9v6QAdo
/hcyUaIyP9BZNT2pFhOljDu6+4HqOkaFeeBCIumi36GGmxaas3RKYDEVJmp+LC/5
5ZiLEq7QbDjeyLCVPs37HxEglC64C8gmVxBoVCUfC+T7jS6c1DTtdvpuKBu5cWh4
0iYCDl4GADrgW51lf5wv0zJ/rKDaTDLGptyv0nA/J4Xlya0X/W9xoPmwBzWyBK55
HAa9RwICyP5D/G81CrXD80ESwMiUmntf79+/R9Pb/SggWR1Blic7rKYgc9Wmtg87
R3xEU7unF408KId/3fl+Jfz8ml3o/noNdQ0liQmTDl/qqln0uC7MFRjhqI+dUk5t
xGZVOIymm7katxNRYX2JvGO0KjRtkS4LiqZZebNBta2lT2fZ19mdC/IkpyzyP6S7
tFBvOXzh1HoOAMASdLxjnmNrh9xqXMfdvw3qQpD+kkmKSqSeZf3jYbcPI6RdZIFW
G4i+6RreMaorrNG2zr5qn3EOLnxw0DsVqjObPC6WNxcC9tutoWnIxeLm5Am9Mltk
TZTvZL41qkqfzd7FNJjQbMAjERyPrRTcIJfbMv+8kIVt+sPDaCW5xQ86EfqbFwmE
JjlNeK7M7ykXWgamCgO59wsfmvAdL8ZedrIRW16/XnUXC9s0tcUHEBQ+RgxOmE9I
KM9f+Q1Y7iYW+X9pKQfsT9saIJ3SicfwObpHnlbQ45ti++xLQC0YwfjJAby/LW6P
f4wk1GAab3a8vWZNt+p+fiYjyxgsPO/MzGtJi0a1y5ksXwsvzN98ccL+lsUpjSGs
KIfhk0ZoG3Nr/gVbkE+25vAW59b1G1UOPqnwSVWAVJDIyCUNVZgxJWsgYcvujJZz
4e8AzDDZhr+v0L2VjqNW1Xgouwpoy9cLgTxm2QvJQvLhuMg8qn+meds3Tkl26psa
oR6BojUQLgGQ/TN2QVbxbfcQUnXydryWkAG/2bajwPj7It66pa7BDvSABYbD8LDC
XFB5/E1uSc5GBD+QmxDWnXUa2Ye1A1dtFun7Iz3F77RS6eBCjgFuhesAN3U+XT7p
7Uqwmez7+GMZeuVeCEmCNH3Eplhwv3gam+x6O0/tTP1ir7f1jgxVicgzuk7N2NBJ
Mvbe0QYwQEz7IzU6eFVIvzmSUNtg7EdIgGKDPkEd8pNQZjC0UuodPNacy4W4HcTn
oz2y9GtBSBOvL+jvilfiaVr5e8y/lWlk2PMH0ZXIoZh045RqR0qszC5VzxqLgnPd
Ph/rusRq2YwcfLWiyO0Qnw6IqievQgXPOxrwHJ4e/1C/bM3iHGl1a+WuAsH3R3fZ
qvSuaR27ftgW9cJx/Vh476Q5tOaUPwopBci6QjoxRLbKcR8OEP6a6Ubc1XgkELNi
0dxUMZO2D0ljFZhwSCNVgYHf6R23sT5CZhMCMQvJJfHj1svNHipSRNdFijH0xu8p
V9PoaAG6/Kw+JoB7UNkLP8Y2Rx/Q5fBBw9kBBEquoghreqs1jlY3mum/to7quBVj
hYqoYPX8M5ycoXSjc0k7g7HrHlS0of3FXfOnSssdEKa//2dByIwbxV1s4C06/jHQ
EfFkaYCSJO5GFS3pTcMQ8DXj0YkWJGX52u9sZoHkqbX2LADA14U71SgdkJxGYP7X
oQ/qpxyyW5fNPCfIs6+2sIMPnWlKag7dLFQYAVCdRRgnFmezqTK6Ih4+WbKOk6Xf
LM+Ex4LKFLzxHGDDD7DYTZtoybBYVyRHmiLrf3LlMi3kHbpkLqxguHE3TfHKpFhx
ZGpAgBG5vdD56ll2COuFFYbRe7rJX9Nv4MBL8z1WuIT8kgH/ilOQfsM7rWqlmrO7
4DzZ787Ct2bxapOgJsWxQ3VYJp7VkwItbW1UjKBgWKz1r8VNsBTR/B3pv9700n+o
FYAvMj8mqw9T/+3K9Lwhdnm1q72cKArF4/ypMjTSE0KBQ12qc8HHAvN59I7UNubD
o/beQB8wpXI+KcKrEG1hFkJlRnafbEz83Vyc0SqYe5XkgNfX8O6WfwwLTcWEh5ov
u54mVGGevep+xzlXnknqZBKjMhKrl2Uck5umjyd/nAYTjEDP4ROPJNPRGokcNemk
i9dG2e/NB4EJ329g/BHLW/8H+iX3YsPJiiDIQc0/DvCmQeIe7QnSuAsPlCc04icR
6lr4nPmK3UgbCTsiw+gOd7yAOtsTZGhha6A4Qq3yMsjEybpp71D3geEXICmHRAt9
kY0Pba7invQr2OfOQOxadS47QOT5S/5gEENNl8v4Z9HUOUxHsvzbYpYsdJ9x2dKh
8iHReopjt5zXJivat3vGfVDpGy3fXPDUzigWBfWwcX0N34PVtg9dFvb3VSPH9eQv
YQakgW0GjnoYhoKcYRkYhgQp2UOpBdbaGtvXJpBTnwQeesYXsubVax5jZdTtQDAE
nuAu+ZNFyHTYOzRDpIxEIBtxPhpL3nxX9ZCNIENYe1nR30uz/F9HZ9pz3fYQSOjP
k1nETACrFKI8rGSgtkmNXQq8DEk0xrI4hkBgXTXPfoo8A7/4lFagTwl3VMh47TOx
SsLhj/1sdOvTkNwXg/Wzpys6MNwmAVTLjgGFubx6l98fgSv4O70oM4GvLofrSoGE
F5zxpGCNq9UOkwfk+p4TqWq9JLPmRTXG49AcTNUoOGo2o06SeejYdTkKW+MeHhyV
4n3TLtvEQtL/2jxXf2ef4r3GEOTRXmu9qvyHrFhy0IKX9773K/KRQYFnEjffOcB4
Hg/lnHud5mxz6FLkirO635NpsJEVvL1S9OUy4WLBKGWttux//2BkPSvYcpFblRgX
J4NMA1rmBLd5Yu9uELQxW7e7lv8o019REFkUBNXnwz5+ZyLpQhfaIFpYgJZBpOZy
kq9ZSjY7vZDp3piv/oq6WW42J7s4GvKLBmr+dvnNv0Xj9yfjEHEjzyutW6OA+AMm
Ntb1o71qXCS3s7Iv30lYOU80yVqfnvVU5EexF4ebTc8p68tiqtjfjiTgaaqR4aW1
UHiDMn7wGVQHupcn8bppKbiVkpZ4eAnpbtVZ76Lap3v3mJGBM2FBtH1z/TOrCRa1
M2dF8FGma9bNd6UXhNwrQ8kQaEFXCRYDmhx+ehJeNMfkMppMFd4FVGXuV7dex8vJ
WhhQksjmHs7XPdlcqM7YkM29IksRcOkuAv/g1zVwobIxonbQO/jQXJG9V9ShJTTw
wjluN2iKnVRGRj37WPSNBVrZW9Bjyjs2DlTmk0QYd3KsFnwf53mu8sndMfUt1FEm
MsCoIidaQfyNUnvxcv3rxZWArWSJHQ4FV28Ftjq7Xo0YobN2hrY+TvHlxl46L+Nb
ukIs/e9NViPhM8z8yUtuUY0/gH0zmEkwdddKonJ8o1cSXKzz92S/9QywpjvpzXC8
PBV6JbewtIxtEoRLTMfY4XuyMqQX2y7CBlmXbIq2TAIAUgh4mMcGsTpILANG3eQb
DbgivwUowlciCAPtX5o/Tr94pFRQbNNcNfPJkxRWiz5hm0dNRd4ZuRRQJVrUMSBl
ZeeLphdfNZyDo+pTB7/W9EoafEZeTyq0dB/LCD01DE1iuEGQcThajHz1hwn2RZV8
cq9jq6lrWrHP4ktoYKJswNnrs9mL+7QmrpsxrTtLKHF1K07MR3LIoWNV4Cahphoh
VwOlv49VY+WQRYSabVDQkX+IPTiGC2qx+kM+vYx5V7PwNt0tO86C+x3OPV1t0mT0
+/BH2oCMa7IpeVbeVJRep88woSXL7DGnzHCmS5EK4XlArbaSa/MUO5rkibYNv0N3
BHuYmg4vGl21bxSSewlERMq4//l86TNNoSWK3uiUD9t3aC4A5D0CvnY/RL8blhpL
pWqeWudBfVvaIJYeUk2zx5ENSiwKa4Sn9rJ7ccyJVqV4xtazsvxTlY3qPyc6ML2D
1B2SIK9wUdmCusSCskQJBEhSr2SMBFO1Qn3OHQNryUxZIpGizyD+xP7Ng57dtKFA
CDoYl0kbKg/Q8ImnGuFvYISHTN7s/wkhaDGesI/U0nY9rIEAlwUIR4ovmfYFY2Wb
fyETK5fUR3pILDkVujpBV/l9WZeBuJW1fVXRJv6WGQZN3Tnq6oxFYxyWs9r7nu6Y
fHMLWVq5DhmbTtNNtm4/2SkbS747/uUVDAo1j1SMS0n+vdL4AaqwhIL6tm88o4hF
bkuoplhQcUWMaL9oFGXWkt1gzyCb0XNna4i0kRmQrjyMc48DcY2UriIg/lVDxFDm
gm8+4zYvPfks7eKACZEFQRvoG2rmSEx4Xf3PNNwjAPQCWwS3o0tx45TpaMbDKHS1
SP7IFqAHCGeVs9Voug8ylACy3vXr06/CJRBRhQ34FSr5T/rGjZmrWz/bYvIa611A
unMJQP7N8z8OeaQLeBhrcPy8cZdeZEj7TivgunKO+2AsOCPyL0O8AwWR4LZgW/S5
TrysZjdfgH1DUNUjwMFEImZw/EW6p2zE3azCyBOnhRqmK8hLCsfMhtAdfnMJmLBk
saki9bxkhbMasGJnU3Vn8uNOSfEy3Gn3Hz80FHlaq6ifOJZhMmQ7czHkK/vfVZXr
j9Q23Bsa/ucbjalePzCeMROENK8DmHEgg8S3i6z1NriuQOKUiorU9OtOUfwk7gHX
d83rte4jDdw+wrk8Ce4Tu/6PrtaRQ21pq7BnuuwHibsrdlhWIhheDAN30tIOqLxS
R4pAoWdiepDlrYNIeTfTEfbB+KNDwiw2hWOCAjmuPrxj+YZEgI9Y27ncpEEkmQ4e
/TtIS2Z5d2J6kAIxM/hDhmMHGKarGOaYssO2mZUSBecuF+hyVLYsYPSkst/Bd5uk
NJ/JGL/gWlVwx2/g/AD6udZF6yYw+5PTCnnLAMytEu+TrS7cuLBc5zYIdHqLdh53
`protect end_protected