`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzcAd88RKffVsQ5om+J3eBoEksCuENCh9aLKvjtZH9k0U
sLVElb+Oaq6nObTmGNPTowLrssUjW4ETcb9iE8JDgvAIojhCX9DfTetNOfOs9XfG
w0BoHI/MDyIVFkUHfLdZdv7soqMEAxcNVpbfF3vpMdteBm87ijdswJ7ftMiPESbi
S//xV32ndHdqv7JykKocIHPi2+5ZUN+dZp4gGqZ3GKvT80icmrCEVJffR+sLeWuu
0P040aBxXDqP6g0x+uXlu+00rzrmNWcoRW9jh8MW3NONvqeLSULGrufyUGM3gMp1
PaKCk8o8jegL5Rj8wfn8XAJAfDCOcoH3m6q8QHZjduWaNjNWxEHj6qTOUpE7aGy+
vPJ0FtzzMMLMeVSZGfO79PYakyd6vt66x5xdF2PdOKPvxrPo/6Y/mP3KH6iej3zY
XN4p4slB/wHRkWZhVGk6QVB7IrtzXKqKCMvUFXwSQjsy64bKuJcFp6rUCTDnkvwn
qIcHYZyZiL9PLl5ZBwtM3M5n/GsO35DCdMFdqcO4fsSLtXm4xiIVzgFV4KXQ6/pL
L0z5z+NQnyC63cmCzToFmqk90A6uOgN7fYhMC7nOAvkQWjA+2oGiz+0/uxCcOHcP
ftuFjw/EQx0cP9eJF9cCFASH7yU80qEZutW53+DpujifTiZIwBIgn2JNeOIk5FlQ
KePhjcb2qQuV44yffY2QWn0xhwxKtUcjw3w/Sd6tFRY/FwNEAiag5qAlB5MzcUSO
+gNod8FKYrTrL9gjbnmDVd8qUDIqM/OLCO6f+LqID4YjpuEz9ANCnJKIZSwj2igK
J7bUgwTx992BqZzxZMnaH3INXMMlULau94WmCXlhD5kxTl3S2epJeXTgdyNfeRUv
8il+7A6XWw5ROBzFx9ab1OntMM6gqojJIMZQjfV8vPqa7Ak0VsBY6bLRFz/635/+
6WWNDuevHqUDxJUOcUuxNgcJ0i/NoCyhTKf4708beTc4qHyFR9A7DDScmS7uRU+T
/2txEyAogUw5h0kLV1UqERXQ0HjMmcoIxqafSHbpoJ+aiDLNhBSb/OlDZmSjsxEl
XzeyElcjCIMwjjJ8O9mYa9l1jz0BWc16NWvGhP+C7OwXtXpBN/mHwJ1dokLdldUr
mikVx2elbGrvsfPTUSjaIpBtKGfUDeyzbSPKsilF4yvYqL1aaYf99IIbu/UUgSfN
aBu0AEGb9jDTGaXyjQJR+97XsBQxFD8ABTDZB1E0QBkwN8CDKbPUbRedHCfYQ/72
0tlnVQCXR+WgK/aGNrXaEoQCoP+6FDw0FSxIWHFvkQkM4F9+/9qBm1csNQObMSG+
xJY78F4P+WNkETICiCjPVcS1LEs5jZ6MX7GrFnNzizXNoSP6XSIbLzliamRJZUAw
IhvcLA/sRNus1490oj7nlvDitGfzyCFg8IJd3qg4sYxZmnvYpILNLcgEKkZ9KJuA
hCj034mG8Q8Nhhw1XNuKQXX9Rj9nbo8IC3w3XT21PdUdxu9zbYS1w5+GK8PCj4mj
HQh4iBfMPowJ8RzfPP2BnfJRchj+FOEfqwR5FOye+qQ3XqSzLTxD9D3GpAn9ryWE
GgqXRz2qkI9iWIk/ZbtiiJy5q6ZdSKU5waLqU0ovqD3697XWJtUI3FkstaOnP8WK
cNvsEpw+GW/c5dxcMaK2HemhJFq/JgGb/+lPWFP58aClXRRJ/RvPfYQjxxDPYmbl
wt/4p/Pr6+zbph0CET/uzhK9HrgkVBTgKdRPIBcgqvNmcLAx68dlywh/tYix5B3S
VeZitlYnCRvuYL1leNJYg1Hxu6bqqxPu6VbfMpPhSEawMvX6s9XvsEmLPYw+i9po
r/GJ1/4oC6jy2slwsyNG3eNML9TbrVDl97PNgnHPRIqpJoniOY04OlXJaHWOBl2a
EjHlsfeoGt4I2npq+4VpfzK4j52qfv20jb0Kc5xrOS44BHH4/9P8ZPdzUMg31isU
qNdi4u19CXUhRsNH6PY3SK5PKBEmEFoRanK9TiGUtULEM/htvPkpkPRBDnYu69gl
oVOobUU8mA8D0GHbYuCHaih2yzGH6LqoQwM9XZejFMzTFbaLV4jgraOT5zNyREc2
t/Fo60j5ShYuQnePIsBO4HQk+XyI1p7CQSzL93d3QFAaLYsQ11JMmKipi0KdcFgy
Nm8N3icN1aJ1kK2iFRrvLNFaLhWR8+6z5h53PFnlC0EVOJjK4cal320/4A6ATdkQ
VBxCaY99y/JhG5fESMxW8NkxhDIQCo/K6NIG0cZorC7ysbaJCizvP6ejPKcF0OPH
YOVHEqFHz17TMYUidTgQthzq1K0gfqiqBGzV5xEh/lhQeVrz/9YzJYbh8xxK6KZo
vu+JsiQwCsz714/LS/Onx5ft3myYY5IYnHHUTTApoHaHKDQ08GwDa/kbRVXocdzT
Bqd8ABjCojLJLSczTm0S+k4hFwpHz/LE2qng4B7C//Ro1bQD8ZAqZM6bozGe8Gnm
T4zg6CjLvIMOKu/+faoZ1vt9/aoeZaMsnuhAcQWozX7EW33iggpyRtpzME1nY+gp
XJG4tmk2f/+4ezumEwviL56We7jxBvIo+S/H5aLM+6bVgfF7stFJBNGnslTLH+7V
rP5enhtogwGyaIuoo4MgN7y5fI5CnN+rdgHt1Vm5VkHTeSRdj75RMruth8nI9hUD
pvvyTToy2RIEdG9QsnWR+qh6NN41pJzHBo5nM1RiXWmxY4jXhsBiafwowj8JyDYK
qeKrMJ+4uXIIsvnCjai7gwrqtgQtw62MQvLkp1XxD1zZ0s/tNJXgPtv5msfClteQ
Cp/qim/Q5X0POjbMhsyHWs1JbWw1hwnLLFep0QnWJeTGR2s/tLoSgOImcH9edAQq
+2L2FUNj8pKgXWzhJx9c49LAWyJCu8s893XUIQH9HWsHDaYYNcUXADMUwEBvuDrf
FTQHQtJAzQHa+HrbscIXQVhE5omXeafbm8CKC4YfJLXLuxCZZMzop/RZUecliWYI
8bUWYKP4Nu+mn2CxI5Z4QRCYyxXNBhQRCr7iqD854FRReFn844ZvtdqyM2tbeYkT
cTgZ4U/y5SksZ/r9OmburAPwLhFBHl3WdEtQewwkPSuJ/MIdIP3REULj+28sJwlE
4ALwNBN5HNOPgCVUivSGB0FjmwMRDjUYoGMc9voBvuFAkOzOBMLrcQJx0Mg0CaOS
683ETvHrk1f5J7AiWZp/EBanFW1De7Ig0u5nZ0UwF2sah4FdJkBd+PUvH7o9iO3q
RalzhzdF8+PrTFVYoR6okkJ+4HXxTkNAgkB+Rl9tpfkxVW4wckNacX098o+WC956
KwgOsmCphWWTlP7pRcox9nB8eOkkKstEwRWANYsfu3BkXAb4vHjDA1ccQDGDiQmx
ejvv4uVUPOT577Xnvi98tfz0ORIDGMGuUYXLv+N+en74kqt19W86SvQEEQDb6FZE
PQWltIbGoRQpR7BPtioV+SyUkSYsrIjmYgCl2Y4B2C7MsEscJ0R3q6DhJG3q11Up
MKn8PsSJJYzMT9MFI0I+HoUws1q612YMP2xzf1YRVyhQ1ds5bUpYMuvfdNiie5Yb
rf5N2DES7JL+xoPI4GLb96AlU8X8k1MaYVPZMgpUh1ErKpYVUqDs9F1RmKIYu/A4
jlPn7p9J1Lmzkw27ef3/RiqMRal04oPgfhoVm/mUVPspxbhBbOdsil/lDxUNF1JQ
xM2mlkM/k6oHut42tanqc1MYx86w4aeiEvNY549+7rg0Xy30YG80RUl9hQk5w2rj
8GbbIk9jeFFHuoUcAXTgl73gPy6pCaiT+luRIiqSwj8gGKZeUXrojlXvCtB6AMCi
p0DZMavT2cQPNjBx8ZIWnRNtZOejmTU7BgcjMszILHhLTrIqyeYIfUxY6MHbm009
Op4ZmQXc+0K3Gz+BD4P05XPmgCGkXC2ngfWd77tW/fhE/r4/7Fijl6t7KTPUo8ac
YW4pGXkRQyj5pP2RmcpUPmwlXW4sYe7AtW9Qg8VFeDqTIDlS5Mli6pPokXds/57P
d30hNhosWkZ2owvIFaKS6hmL8X6HE4p8/DIwbkKYfc5ZCnDFaueBK5SqBMIZwKld
vOdNCyteN/HjUb/A8D7UXZsVwMr9Vv9oVjYgqo/0VF2j97/AIPcy811UPaPuC2+Y
K/zq1k+YdQVGiGYqj+EAwEeUyZg0bgaX8Lk4+sdjEBWgMTs2LkZ3vmll4nyLs1Vc
ZJr/khBgwgG7nA/BZ/9oM369b1cHf3+kRJVdk7tJoBvhj0iXYTX1WQEVFTLPIsuZ
nM6UhForlsAY+ziAMM+AcBKOz0YlXdyoBFfk5GhzDNDhIW7JZgfnv+u3F7yKTzK7
QGyisFrszqMV7rfktmiwv1bu/fBAlKfYb138jGQGl44fAtubnRD4lqR7aP2kBrL5
QAHcOf00BLFScKlxXn190DjHs0l2k52M0FK1evcIllSQi7Kbkxs/0MZk5BDUxWS6
AfYKUj1rT0oEoLBgjsvGj+1ewD6JUHRv/FtJxRsY6x7pOrLpbPuB0/2grP1ukEKx
VVIyDLOMy73IEJpucbN1moO4DubfCzvI6rH6evWkldTtkmvudgIVYG8obF5CcAvw
MLerdA24ornqvDmcde11NngsPak/GJiBia/t2pk0fsoyhlmDGFcaP4ZdtAkmJdrd
h061Mv09jhXTu84Zo/C9BcpGIrT1sQfpoDsMUb8Z8/ho0zEiO10fG6q7KZm5gIhy
Hz8D/Q3Gq+WPQGFTAyjxHbSAPi36pm+Nxw+ORnEupEgFCmHY3wToJE6bM1T57M7Y
56RgNCs/u2i7sR2ku1Gm7Zo6UKFY8DH0/LUwUc1xyWCNYX+3j9T8n+xJOiLnsay2
2VghDKEK55fzxP/Vjo7mvXc53ULJ+UK7NDkb82QRs2VA2bWvT6dyVswpZobTKzLT
ohnWXISWRp7BJEWjDcv+s54CygWt60ZMPIron/LU5Ksf7CMRFjPJWBnFtWPCJ4XR
+wU4ANb/RRmD95rJpQvLFAgRXnspxxAYeU/mg1U3EV0Oo1pTc5nqAlJiyAcV+ux0
DzJbb3HjAUyCyrf69HnfzC1qBq3zEhZxPT4G6NL9AG0eohjXjyPM38sAywRBe3Na
/CzNfX0kNyESko6VWvCl7z+79qtk+wKSZCVtgPPAFcoFvw+QiJXSLMJdl+7k148e
6zrVxL+XWbsqltFSSO2OPZfRKitazBu/ZSxOB4GaW6E3vtxjo5KW2kymuItkiBcB
dLPUXtiZK4CIws2MyRPKAYi4mwTQRsAULQeqjpkwLZwJ4H75Nx/75CylM6R+sxxM
yJrJPjN5eg9jJVvof4FWG6pxSZcobDyJFM9NfwFGO43wjpFZqm+32KzlyYLD65XK
1OD3U9DvXPhwKD+Nb2R2itD5rWRvV7UkGrjcwNto8rYLB7XMcEpoO8PtJMGPT+RL
zsXGeYMJAkhheJAv+a7iQBkgR1unOwIGXAqfqsCL9KV5kIz0G/QSR/eNoqsVzTG0
CiSsH9TFpVfLdUCbIjXXZudD3FB18AmTHPFA2mDDcsVDUQrp7capZRmqaLBkBrV4
r6f2+wiu4/gQn2flXkV/fJVrs2HZxt6pu0atyNVH+NroYstdDAY52o08ViRtkacB
RB/OaVAKZuTPtIcIT3HBC/E+lKUxQKRgu85uHkgEqESpmX5PJ2m9krcPVXj1BDcH
`protect end_protected