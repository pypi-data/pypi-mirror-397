`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
WBMQXuhR3Tp8WpycoLuICqRsBuvkJ2Sj2O0nVaNDFIgq7OmrcRyINUjCLqiqkY9Q
GdK47ZHO5SNE3k34/mEG+QnO4HnTOLeys+kU0HAriwSJ3vRQTyezkvCwz8hcpPYD
8L3zN0K0s9EoFwmOCVWaSaowbYKT+fe3wNNebxqmWE9BI7cbCGlhPXJHnk8M3aJs
kh95wStDPggX1yvnoKYihWwXJ28V63cj7qF8IeicJ4Vfr6d6UM4Y5l/crcR7C8aq
4uPvVOsqVvwsits173Ds2goYsN7bq4jGInfnueyHNJOiwqE+n80HwL1e5lY8c7sc
MsW75cCxk4MgF0fZ95hbqqMT7SVCyENA31oWMmXMAN6PR68/ACo5zMUxbs0gg3fC
0fRrisQoesBwaEXVVIrnzKCre8M5S09iAFsOyz/zZqt/mC0PNsttPTIw1w607RbZ
Qt0I4QgyRIJlxVS7EczYrN3Xvc5vBehLWwbzRYDNoNUaouyW9BpBFNdWeze2BhzG
YOfiA6zj3LilY2sb9/1hNvKaxHMk3IUD+FoI3b58xnaQtELrydv0+lux9ayXex4n
yYU7S3xf3EvtVS7M82Uo6TryWozSKVQ10FDPagIVoYa1fPxa1lUM6uZbFvCpMx6N
EjCGBrYZ/125hF49kItW8j9nbiQhJx0IlxaIucNZ+pPAAimVW7Du6/+tVcua+Pf9
6eJ20NFl3PtC91HWRJvtZwe1Q0DnEFIGKVJ8N/6JCuRj8tFSXT7cUAJrUCtIBPkD
AG7J7mUqDD5XzdEHPzS0jbPW5ktC5OTuxMNw3cCtC+coUJPey1Qwf1wdoGiRk3uB
VrACOZY3ROKOXCc2+XnmnTakLNXGfHPHqM6cNr5p9ym1ZoqdrawPwzznAjwKBbTD
uhdJUCQKZeE+1dDbaGrPC/1XcXN1pWBxmPniQ68EmaqEiV1ej5LpM55UCi+UdwvD
MIqHHZ8Mh5SO6h0g3GF2VrMiSZM/KVRDY3FEtJNFl1PbFw6Khxs8zvhNIaKq4kBC
eCppSzH2+ogkBoQfDAbMEQS3IixHadx/kBGoKtSpBqw8Vh6LFDqNJJonrQ5LzjYl
th4X+scuhgSq2IhwIxRaq+08lWIL0Wh84V+c+c26s1ZnZKK5lqIfWLN09hfokGr5
/GRo5SbfrkR26yznKeZK9/tAgh97toCKXV4uxP7WVsDgGNTflnKq1rAOODR1cEAm
OrDj2N2RWCGHvN9X9WMI1cN02cnOcNJE1TlFfEfQVTZ7rcxFruuhlnWxxL7F7uMb
e9CMZ+O0tcaKCvSnWm9PGDmVpLkcx6exETgwPDquK8LGaR2SK0jr+kD1pJKFXOr/
m57WL8bhIdH8D3uUzRbdRjmBWhiHr8Lp2kLPR8F8jmfYYn0zYIJhzS0fwxnM6tIp
TYN8i5hQX/cZrxFXU7q5vv0OTC+AalL3fCIV4FdwDWDEK9qVsVB0Kv0eQpMfX8dg
ldsFStJ3zApHqPv48cgOYearVBEwjnzN3uPVRr2Zap9s6cxueEyO18P3leFpmtct
UhyanVpEFKQBJ4Kqn/ga6CGaYvGBbxP/MjHPmJCOawqzS/F5mSSQs6Dr8jg3VijF
7vK47aIzYT/9zd1KFGcw2v8KmL868rFKUJHSzXuqWkgl42+k4QChOdVaIZDTo49w
hvBY19PbawHcYmTuLQpkeTFvwohX7HVjL7ygnLAJZUhbBR+uwV/vmVc7/uFnNhPz
/2smvU0ESvYUmEoafKFmthedUDENC3/ubfpJuidN9DAgjXGded/EBwULfWnYgNah
BE7/NmhPzzSWbO7sl8wHJm7fwwc2386KkxCZEMPftofdhnzpUl85bt+BX6PIT84j
jG72DLUKWaOSxheQ9DVGZvw7B56zcZc+On4A8wdu8CY4+T5mRs8dPsmg7+TuLFmz
JiqRuD0L7RlHgWfuwTBz4rrAyPkYX9syqzxv3rxsNfbVx9G+vTPsHbLh4VxVGpP5
ooNRz8l0/hQx7xxYvwOo0OFEv1QYVzx3CpQHVKoC3OGmk85ohL3Idz+C4pdy2td1
ju1VhqwKq6iicNHY0Ca17LHnRiISpwWEhjktaXD//Iy5zQ7xR0U4R0HXdNvEVTgI
w8UCYGl1px3i6aTa+4seLPRmaevv6FcV4ndK9bsjt6/l+IwvcobejKAWTJamfI+F
z6jBhoKUcuIfM8MG75ZGhg3Hfnn15p4SaHDxVEYt6erfkWeYsi96u7+5uVu/oj50
pl2eTlLFuIqbfF1cl3AAfIRd/nQ0akUHytskt2ST694JvGslg2mrqG6KlmPDLRoU
CoSMTAaFeVGT1UO7jcjaeAJlzhz9ydm+sEG5BO+GcjhZshv0R9KPlY/8LbDhw/64
6PAokjCiSDDgmVhS3yk5/5R9fEEBo6ZnhX1wqJzdGjwfl+Ozwj6ov+9u2Ahdl5SS
zAIR/VPkpmnZXwMLJ0d4SAJ9JENLGA0Cp80OqBBDyuyKaAGhpjy3pYVTF0PSQQMo
TViim3yujwtJVxd9i9O6AQS/6Qz3ijBW+1ZVb9szanURtRU9R96nNfrPtIXYdmMy
aRubQszS09s7xE+5RJ/pdmRRb/NctbVZjtbFvzpEgxBLvZlDuI0QyzfGem3iQAKK
RTdA8yLfYYKPGY6DHDAJ2pOI0PHZ8wKLsKAbzSOkHbiwcPNNZlntN6CZKe6tF+Zn
86Z/MgS+XsPuDUMFTdJ1rOuXlwtkyHcqWeYCq8GDYXwDIxLvx2aiHawrNSv1DV+8
cPKQ/EPPHPRbuc9BxLP+fZFedCt472QIcTddscLKXlUTUvDdi4EYH2596+mkH01d
AnOcL/+r8IdflYDCZiDemC1yfvhy06O7zXx6hvvKhb3YvIvYlHM6PZMxA6jgW18e
WmAE2BwfncxBHNT973KkPleeNHtPZ/rAsZLPba2dCEU4m1w2FZ1trCa1KKHBEFRG
bpJdqWe6S+4qF0l0z+RSu+9b3XXPCV3pMh3ED+FiEYsi8ltXFulGqJ6YCYPu1Tpd
d/c4Xs+jPgznKLpZ252pQ74KtzBSCnkV8DaKSar/zwUgpzGaMerjWLfgIF4XZJAF
vksntvIx3r8090lp/Ai9tqgOkWa4p46RTKHf4VDx1VkfAxd/LC2uEJj+FpslAQGv
uPhho/Q6dPIFo3jgZx6bN3LyHoP9+ny2LBy4P18KOQjqJQ9M8m837SjQ8rsLkySq
5nVFP7sLrjrj7gCsyTCjuhCimMjB5Z90scNKeqyD09qM/k4ivMpAz3Cmf2rg7Qjw
PUGWbpM8KzEISs6qOlCiqT07o8sHcIuZvL8Z1OkJ5QcUnsmb/iygK5FOkpgPaOrU
WZpSK7qoivl0ZNeXCL96hMgkQ8HCynFe84QgqzxU38pDush56YpZMcslOrNvknrf
BQxvJKH8RcIFjTTOC3gBHlIVb0Q81MOGIcG9OcmapSyP1Qk30LmBTE+1MgXYKRK0
8IcJ/VBFRI2rFnspG6n/sBa1ZH5ZbJyBZ56pUnhGV1dFLY3pESJfGmZrDX98X6O2
JMVetU41yKqX5RIVZioDxeovtXM5jLzEmV9+nxGp2V/2rTwdXMpJn2XdnxJN2v2O
hcxwMe2FYmzmq83kq16GZLu3b3VN2dHVuOF2iQ7rp2HEDQhK8RffTFf6CRkou8Ll
/F0O5zg+YcuEUNxrJV4vkM2A3lWsbiM2S9fu+xeu5g/ocn2LNMOMPv1aGCbLuuj0
hHTx3K275OSbBUu1Lh1gv8XtkRPpkrGoxVHZbPgR8jRll2aLD1XJOUnz2/9wgP7I
QV1GoQK0wevUiymv0AziteKjX1GHCETlEYUgBcegtbSaFvw4Et4L1GnKEIml9mbk
YMgTs5g6XIyOu1OgSiHG/W+llc3NjuAfEvEfduy74Umc6nJf14D2z0Z3PpUx/d+q
OVM3ON2I/yvm4CjUSAqqNHAL9VJYremaVktsujlmwf/oUvPv1+YeS+yqLRmSUGyR
BVSnc1sk3caZQvI5GSuEnN+j+1dUzzvI5n1i7n/VYeBPyi8jBih8ZNimEq7WpaeN
pKhnvYSSKnxYKOsSKxI0eu5yCp5ApSVwGRq6cRvNuJrdQHUxzAa29U64B9cU5QzM
kQtr0Mi8kJBI2Ne1sqIXIq87qYKehGFJLkrIsiOgwST6tXLluQ5TyoSH2c1RFotA
pCNksJx2gntOOWa4ydcVYyTurumCqzpv2+fqJgJd85w53h/osrOBdaCSNPgYZKB+
vTi/mSRtS7dn4F2sD9n7BCSC4SSgAbHGbJBbdGfJ7tI0MAQBWJvCa8Na+82pvd8X
sULKnmysE+VSEgq5uDmJdXsbYkNRDZvlcXoxEOdHBiwobQW5xOp8WxKLPU94obtD
VdqUpFDY02ovXoqXzt/YduuOhRs1AvOJw/V4N45BzfCwjlnU7FRXkuu2hS4He0wE
dRMOmXgXAikCg/XziSbggXKQMY5U37c1JA63U95ztgyWRISX+ldsk0wg1WCPylzK
TXI2hF8WkwANGHH48ZIC+x18F9UocGwJqr29ygKwSHLBrT90CjDxSot72OaEX8K7
GKHvr+LLWEfEcD1LQ5e0MdTIIrvhGn53ztCdmRHubengLKDXksjUN6vNPeCgiHFj
YyDXSOzHkoquRYOm4vdPDYbKMF9zoATvwTMAaMvVkPyOrLf3reZ969efsZaObohQ
CV2Wy2saA1chO7Ir6zT5rROxH2C8DBiUeTRxuiPCQXHA9fWnstk7POUTURj67oSC
EnzAe4Xcc6um69phk8TR7HS5rMtt8Ni+dYKQJnhEaqOioCEfVSOIf/edH60ZdY+5
eKS5rBMLY5kjy2I2ynJuGmDKcfwDJuzFt4T76p4a6mNEFZKXasLGC5LZSdZsff9j
LH+nPvXO9VkjVE12LJWThQeav3GDiD++KL9oNXwmPqbtbrYoWf52SKDnAa839S5b
7iwfdCWu/rcutddkWlhHI2xCtoJW/0ZuC96RV/0OXQkZW36jeeqB2v1BBvG7qLa8
rRPbCMp5i8GTHTD4+xga/qX519rxrDs5Q8s5tKQbsPE8UszWdAJvNRI0H2OcoVF8
u/GWFaxUyvIqhXxpv4SbuD435ypkRzcEi028IwANDPtlDh3tizbpOecgyZ4TFsuj
PMEJ1++sWB6k0Z05Z+LNMNRz7Dw/DGkZ481wQyOL8adcVtvCF0wbm7x66SbsIEJa
iowoG0EWUEzn/DqRoBgWg8MpnFZl5W4mMqIKhI7rgIi1w03jG+MnMyN8gRjWbtl3
qbpIJGdJSvXFDEqXGN8viqX4xQS6z6KzFOddkoxg3uh1zIvunCCt+77OnvCsHng3
SJHEST6HF89TShIxFuBizjLbjE6aDBjeT5D8r306Tt4z2pcsDqOdrKUIrN7U5zzE
8gr3N6z/6SCQiOlbNWOeSp+DdIkIC4X4TwjaSgB+LxV0EFOL1L0+E+QrFZFeEBgp
cBn81qksodVlVgMSh9DIWeh1FAKbhPP7YVfhEs76wW+mvhM7knn3tWXlIuBmEvZ8
xtQyoHMW9j62NVm6kbqMVkY3RhKVB7Q7wR2juJ/fW1rzKJpTef+q/Gk+PtDdhKQs
QY/TSPT8SPNvz4NRHSKGCAkr8ryKIWXlwMFvSa4t/WdAM1e5ruI1lu5tjWBbFw15
vVE1t5tEKMlvF4BPrSZX69I0uZrGlZMtdQ7XQjX1cY25ux2pUoDfgF0at3pEW7Yb
oI9gc71IAtqKlNMKUxbFuTeYDiGITQGAvq/mpftLoTqiZaBuH81sAZsSrcUg5/+F
qdfuaYiCDMEJ5ERx7RG5PTks5HfeauH+9nPN2iBTtL6EiEIyopexSi/jEMXsFBZx
0aH2eEm5rUdeI6GCCchcrsiFtiDkQJffGfudTGctwgARpYZOr+qEjNhmCxk34125
Pmm84Jdnm8BkVXY3u6sQwGRqDCMQpx3wsWjw8VSQfQ8qRyCczOReqpeHi8nN8Lyq
+3oYgMuRwPmhVsXt8LUcFSlD4K+wn3NYcvp/hqYNzW1tOoD41WLpx5a/C2apGuQq
UB/87+dcUbq1ugeDw2LOjkziMDto2wXwhNg0gOtzjLx/CkLED4NYdHDlumIVY8Fa
ZfwpO9M0Rt2aai4b0hHUbqPnHcYXveXYzwMMWG9dZAVrlT/G7ctyJxUpg9uIcmV0
NRK7jt8dfG8hMFC+FGhu5jY98Tv2tgcTdWihOFwXd9ELdBE5JbcA4s9T1bwNq96E
N29kXO5/Y5kanlEeRP7obExhs44h28odj/uzMIkseMtTFvxwEpooOYbIrqJ1HLlF
hzVTojDhOPWxl/FGhEEzYV00WN9LtJzZuKYZ5r7SYphE6YkTcuO/JY+e26QXKxVk
Ua+sqKKlP30Q10n4AjhYpht2r5EURrc5RtK84l+dNYIF7d0wIFPhGp0GekT/YG+H
YSuPgWAmbOo9ZDSJivjCNUjT3lOROi9P/cpDTTweP/FmZ8C5sb6cV5EIEY1DZSsd
SrpAHpixfwVhKNFKVqIW9rlyP1AcxKrS/l2990WFbr383Bpgbc/JIC0MmGaOlDiP
Z3LSwVMpfOg2ZTvf7+cThFPaO0GzEJ+TP8pa1Vz01BVB+DQVMbvN1ok3OQkS3E5k
1mbuOKLNbENWfAKnESCgq4c2HmHitktkjPHQrrc3hIdueK2KvDaWxbpiLMxcgEiQ
iNTGLK6k+135+vtw4Per8Xd/0KzdblNHqHAMOhupvreupDaLiXDATTiZam4r18qQ
prgwQpQVy2FwHVQul+xJ/BIzoZMVunIjzRO47ZrLivcpWsugudH2NO7PuSak6Qx6
I5vKuP8b70YV4GamKT7xvQ5YmF8xe8EP0sIDO8sXm232VK7ZKXlQkI8mt6WSDaPZ
ZbIjlmaTYthyjxHgGKvGvn1I8Gu/xEUX09YyA4Huoj391EIrAqfgIxSC4YzjXTsc
SWKBoDxPBGz5P0Y6Yy2LwrIcH2dpAHBG2LhCDvOjWIfJtpAtplVrCldFxYKDLOdG
SmvO0l3XaxWAbA44Xn91vNl0xfRFrZvnGTNNKDD4NdMd3q/2kjg/fl5T2d40dXxO
Yo3agIcGvLSlA7vs5NPwbzrFHQYSrG3ukzQ2y78ahWdB3GzmTWpW9Z2cChoONp4K
T4cS50Hqwn0lQohBm54cvAi7GN2sppj41xq+dfntz6uWhyF/tPbMyaewfiL+3HSZ
HjsHY+rRiax3mj/Lt/Tng4fsc7i4TPUhTEYd1NdfXVS9MJRrC94WhrMP9k8LZg1e
ezfeA6vhTIIsYJFxS6agKt6cQAc3bR4OySsCghjUz99b+QjYCT0wLJr+2TMP/JDY
kItEJoMmaKtUc5cBNmquWqVvPTVjinp1yGxew2bfHJhALjYb9QnOkErBQ3jYq1GG
pRKiaZlBxjX0x4tnFJvyeC1V6hx3ZYrCddETscUmU6/9WhWLcT0buFLVNqpfZsdU
gi7xPHug3bGK0h6BVe0tV9/4hO16iv35mqPs+U5h6/2KNzy5Zs0iQsH9nsjthsdo
Dz3YdKa1CSZuGw8WIOmiW0uMeuuz6PAjVzS0reH8ZLa/r8CMlM5QSiXvLJIwpCDZ
Qx15NTN47RBMW1JvImawRi8z8yA/QnPYbA9v98Ui9eQHX2I+iTS0r+Goz52yCKFI
7LdnHh3WvQyi+CBc3FdOIhIlq12GCyaoZVRzJWZ+xMS32cKQkf9hh1oaBpTHagPx
8N84CmWDb0jFLd2gbf3zJD5vhacSf7vjRoHmZwHi1FQdUNubx9OcnS5JSMJmXXO+
zlmlnm/jikkr66MLxHHlR/akbFkhs2O8tnz1uBiNWYL2dU7krey3tWs+O5xr1IAh
yZdrMAHfUTqvuZABNRXMmS2MT1gw6vGwtB3LAy3US7pRGi2dLqvr6bw7LFrcrrQA
1XuGCMIWQkp2up1jxS93rLwHdW/zf3St51s9nlU+YfSRtpyZ3s52m/eN5haCiRhU
T475U3Zo3t7N5c+A7Hf/clGweKZ6VKaspFACPizcAOzjqE1szuT6Z+dYha44Q7TM
mWIRekTIU6CpYQRSWz4D45sWCEW+RptGEGefM9s4SWNfZt+IjC55LQ29O2rSJRCZ
n7QdvrmbfwNvKn6hNHA6QAJHQFtpyBIMElMZSm7NsZdcMlrohl7z7XlClrTC3JQ/
68n68xqQayGbXWVZQcIktdFJyae9WvRwNcZSKVBN+4ISdSIirP6jqLnymrJH3oOy
6BagAd4UoZ7PaTtCGa7lg9ij1w5MzXd828DX8sTMNS0hwH/Bc2nqHl4wHs5ZhBeh
xORy5dLe6Bezg7+Bqpgs+u6d5yTmXJBZZWUBUhpBi+tZjvFCF5pcZAnb8p2IXIjZ
9asbCEx5dvV4B4+NpMUJxf3aNzUj0e57WsRXESxITGLGgCAJD1leacePBAvv8+Zj
S/QX6KVhbsAUoJU0vtQlbtb4TYS7ULOy5wQQ3myBBJWdVwEe215mmSNC9o3s9Kne
GWjh82O3/Zeqv2jN+gBaur8A2wwodQDTkDbWTYk5UHwfCYdDd1rz8ma+puXn1lJW
++u95kzVNk/C7rYYH8BhkEEtd/BYcguBxoFJidgzhYh0XMwgSTk8YQvR/ho4yD30
gL71I3f81giyVOaKHQTn7wFhuWkJZo9HnngWZevdL8wczuhJ2+X29oytPzykq1WH
ymCgv6TIdrFsXneUuEYhz31toxR98XZx4wpf9XrS1fJYtIgTtLCBzDA0RLCR6Ljz
pcWPZ6ymUcNkwAO8juiLiv086CdKCyhxfnSKQOBlUcnnSuCHGBkXX7n+Gwxy7StI
EvmZbK8iSChkMQo7Il7qpG86Mt2bM9iBp+lmfGdeEtZ5YN1PIGFo9reb0SickOP+
jHNjkEFx8OP0N9iJ39iKcS90q4oxFF7StzgYaikQ5xnFM+cBRke4gySca1j2vY50
t+c0bGVOqExUc202tyCVVcNPVDAYnhshSUF985sp7AwSKc82i+Tb6I2XmQ2+UiYk
QWlhx+RYxQkoouFm08L55D97lYqb+8C1sy1bLGSDpwieC9FWUy2cxFpeIcc8Mb11
N33s+JCkkEy7e3b8iZt0m2L0SB2KBGjLG6Lhj7uYZcq2RmSy/uM5fLdFC8N+xjS/
`protect end_protected