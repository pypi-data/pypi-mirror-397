`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzbxWtePNA4xLKWL+TYXD9yilwZ9HLVbLfyGB2cwNQMwo
xBKuyFEnxxnX+FbcuzL6AXT4Tf58i5tI+hY3/fnYL1cn2CDePmo/fWooHuuh0/Zc
wuSN6I7yk7B3YqYkWb4oLxAAnzbCxhkF9kK1zXbj3ezZ1QonU/0/Pn4qY4TpZZBc
FEXghgf7IP4iL9816aHOdh1+7+qVt5gjFNp6Kpkk2LjhbplSrNXEV7g0V4a9Vjdz
9r0yOaZxrskvUkYmipRqavQM48qZaL2F01eESB8P2GwIiyjPY2THM8yam1w5wbQz
juPUrpJxw8xThRM1LaKqq2tu+ZGRb4gyySpEkBB2CdhCO3rVGPLU0+ot8OAsmlMf
yCU0F4vjS65xgOLusX5K6QY1wc5Cso3DqaYSFSHKe5Sz3BHWPQJ6nnWFDJfFEJVK
ZE6ahwqxpgjlIS6smdGMje8bYEWm8LNv5g2X5HRxGWaw5xR2M4I0z/OI/nv8Cvy+
rhENk29PavYB894z6hhMcTtQZHGBWYTRJ2Q99+Z8KB6Bx695GzyvWGuEkFqUxv3A
PVdIZff+H0pNcFLcGISNXu/cZI1DeIxVFWLicAktzOB66HJcHykesTVroM3GJbGn
NRLChRO5RDaD1onlhift6h5S+m6f3+JcNROnufaBcZWOBW2d+mOH6nVsD0NjMHqz
ClQ1RlwQeYQkdruhDJYxF4g05Z56HlvUUUCdH/nUCsjStsxPub+ts2gwS9KNhg8W
nKINWkPptsK6TwHlYlTlbBRmVQMu3EFHn8RAWmX8erji1svigXyTJNAW9Fdz+jYO
7rArbaTSgKwjc0xNHoASTNgx2BFFVQsEz6d3tiwXSHrXaS32Oh1w4wujDpm7gVY9
yvwQ3RBM16/eGndV+275IEaJt73yzmjwmbJRL28yIEzAA4m2hrRP+ci0Vqobz2eP
vZWOJM4A/C3sxkcv8s2a5SQelYHp8/QX/55dDJSg4qU+ML2RN6aTAtxusi+e3TkJ
UB3pWTR4XVlPvg3yjA55i7h6xPV5u54tGZsbBeNTB8bmLcsPlRXlyFeD53uBLf+N
5t8FpKQMNp6fyL2Tm4sbZJjORS2qYdBtpEsgikUbMJFMsNLYh0i5wul2yomYDrLO
DipInUH9C8ftEvBp+cjWwh0p+BH9To+N9qgDTVyL++bJxoVTvdJ751eqMe4Br4Pa
idMjBbMHvPo/+VV8nrJroEXAYai07lN69OLEwb++skw6Aa2OO4DtVyF2FVHSGhzY
TaCqWuB5ZAbCom4n0Xii/J2NRbwzR8kOxYPf+8NjRxQrwBwaozoCfmyY/McQ6jIB
qsE7Q9njrIbfkvrb1CHwZuD0SxgUq5AcNBQiMeetH5YE1kd00sN04x1NctfS75fU
fgjD8G4M2PrDO9UBRO1kREQAPbRJ4WD6gx5B9c2IlYpeb4pgko4ErZMQPNYBD6Gj
kFJOuIP6RYNvUuKnpiqiN4cKv/yzZituUFv9FgpcL52kYRazb1wt1u73cQ4Sq3SR
Z58Nk9WG5+32YLvv4syV9ldhodayzh6ZzB2ydfrvjxkEE/xgOETPAZzrwZC4wMCE
2pwCJ3GRejFmSivkj+65dEGLhm12IhY77QTge1/5KItTpvw8ECCXTZRWzX/1Dkqi
SkXATRYmA+qNYPur28I/Vh43rJXW76zpCRJZ34S37d+sKv8GZ5SZSG9BS5M34Ppy
btGcxUakyVpmXh95MIhiQUEGTJXoa1saeT+McDwtO3ZJfgh4x+y2zV1iy36UfZXV
UA1vObuA8MnGM1n1FGAOi2Gr0elo1i2sn/elk/F3q5ZK/UU+eEbvb5beBgI2ejvi
MrRbfcPF/yjPmbhRqaGfghD5HFWGGlibauNoW2jRq0G1528BKgL+tNBa8iCwIqCx
ImCW6+w2CMzSpTrG5GNgPuNiM6OvsNAbUqoAPAFfnHDl+MpyqinVmbmgDdCzCb4M
NrLA7OGBriqMAjuCnGXf+OizO/EVvniDUR1JKD/SFUnbJnqhhrHueSfEeGTfrfcj
RoKxl6/GJw7iZPxijvFc5tInp+fvYWZm3mPY+VYRdIJznxMVUgWwpVMTmWrupy48
juNpYTNErY1lRcm+9DEz/UHnmJ7Ds/QJe4ZS81a7Dukr2lcfn0rxIb0qUYZsHCav
tr/Bb4TSsUWMiE+/HB+NzGT4hKC2ZqhZD9nxRRRohn9thEUqxHc7PhsjzTfGvn6U
dHED6oEhB+LZR/5dMO0fjEfhCOEmjFhfgLIE3z8B2VhtJcleLQ5Q5hENBjLC6Zn4
85i1sxblKQbi0qT3nRI2/eab85DZoaAny65Txc9pUcwrW71Mp0dQiqonSPJj286v
Qz2OAJpCyCCRWLUa0l452KSJm9Qb/ynh2y3vKMimyrqhJDizBqerMqt9s6j74rFO
MHoIexVZcK0hESwHUJtrnaZlraPOq7/nlIJVU07s33soWgdlBuTyETfHPruOh6b3
y+Itll1ubRZCEmWmdFYsVRBrZ0dDvDZqNAoaJJ8+6HQcUZmR8NnAPzF18c1efwFP
Ub/ynDSP7T3388yC3gbmqHsGrYxGBVcPjdye5ExEkt4dIYq3jpz8/wlIAHKz8PUo
qF1PCj3WY6lqS1S9zIA1G/a24zK20J9hbEYOlHBcW2jY7h7Fh6tWuHgoUrORDlLJ
rjDNriyvNt+/HY3bb35qy/Jhp5HDRGuTvXby80cV8Qvpq3uQOxnyGlDfD7JGTqhE
IdrEIusZxrUQuNhUuwvQHNm540udCVwax0DEOAH058NRGo4HGq8RGyChHHNawz0d
2aHY8wJCBijucxRTYfW5FYlJAbPxsTlfnzsYsJCvmwV7c98NByk8FF6YllkfGzBx
XinMq08d9p6hhOsW47JW8CwsH58/BdmnNU2en/bS5Ja+eryNblKrNw4g5pH1XgTQ
uffH7CKjGUEGHzC6LZlClyESsAjTYOrXjtlRggRLu1UvQNCO0bkx2L+TqlQnrY5n
MQ54OIwpGTnbL8CFXdh9Sh1Byo8YUFlg9gCUdpsnQHoGpu2kr53yluHh0kd/la4Q
w0QkoirZgGEVu/iYWTQPWy4zd9yX4RgGtTNXANQEQObuYYpKX6WiZScdmBzCQTVa
CLzAtjGAW651t63Ik6o9RcogHxMOUWhFcS4TGGB2l4h+Iu5eDCbgqnM7otc8vyIS
6wbr5nSomcMlEPeRb7NgOpx9jfEvEV3Vs949fcyzDCGIkHbGYGRBWI6aeG6IuaT6
aE5slB4r0uuMmtCLmOgv2eLeV2ynYsg7I5QcW1gMx07L9m0q5A5GOpThF0qs9LNM
T3uw2OqlK0AYfp4BcJF1ut6aCDSXK50c9RqcAkb6EIjE5OdXZw6QneNGfxPMyKHi
zoL+i6+UUuBF3XC2zRgvjjZUFjSHtP9w4IMLAM6s/UXk+X712Vs/qg+NxEWJvBTb
/P1VUlNORNAoII8dXFHDTcedIgocK7cvBVHw9c/imWZ9nCIJeJYKcizxL2grTbWt
2THEOhMnOBX7RRsxCQbNUiZRuGtRukpSY+7qWKWGdYHXLkE8xccX/QW60K5iWJ4S
k89F6VN5tRzr3O5u1C6K/FMmiTn/DT8SsQUHHqqbXwNDjR8aAeJqIwa2sHPJhrn9
O0KZtGb7rlPYF5mipadTBYQC2uVaz7u8OhEIQV2Dvh3H4GhD5yZrUudnh1S3Zos9
r8Vp3vFpcZBpvPaRMiitS2eWxTUqhRCpOfi9yg9EjS4esIxP+J20mj7NwMDAvMdR
+yWdF+axjsKqsoUS48C5BTZWESsAmHyXBO9cDd74K5mavKszZTECrvLl9VoNq8oh
B3+Js2nWUT+85DagQ9FAueEhV7wuaIXoneQc8jF+8MusDNyIpqHmgZxqCrJ859I/
paPLjR0jADwfPe1HzL/d99k9LM9cXl+X3p23Tc8MxAg3M+iPsXTZIbDE20d55mlx
zGECMGVJpTGreV1vnqfnPLBErmkTME3kjLkBIjTp1aURECsMFwst5vywEnS3h2W6
/J0fK5Di6BwRoO8l0wccCTUpPBrDllrkW+YAiuj3LGMVA1rUc3jqBOKhj6CK9XUm
7uBGXBEleCKBDyI3JVaitf5UzNwluKVEj9BoewnBk5UHr9q52dOHqZdlkinTfVjq
ShLNeFBIG67IXuu2Rgq2SRarYVsTg52U5UD/CwLXVGVWkhOvNqFATntEecFtuFgh
iDRGsc84+iucW6QSwWcHbWW5qO0iyb0ZOVcKqeEKt9BXLZ0LRC6TvlHwE6VuLWXj
xySxK+4IY1kE+BVBlmyVFF4LO9uupyWfNvfKSQsYEGdMgIQzMiw6nB0RGBWbE3yp
nzlsjAOuJLBgMYxz8UHZbkvvtF44zMD6Us2+VZlXzieGKL9x1UPSmeeraT4g3hVt
CB48jQ9kbz6MxjrG+wwOeIBOSi/z33tqwpy0fPEgHYNHCJwI1iplEkS5cjKlA0ha
qHSqhXS5zwl+Invh2GrvsNEYMbtrsP+0ZIs67DyXFiPBZvMBn5jAZSr7fk1/Gjgs
VGRDhXJtbWu/2GX9yubjUaj/KATOrlQxTPlhY6QX62dyAOXPxovB9uoX5qSh7sTu
zpnsn0s0EMnqMBbQPGtyszkWFyfHsnKT+GGvfwkZwK3dsbNnE2shV3gwX7ERHslV
47WDCYuKHdINd6JcKLgoS7uu0Q2pa5QBA4/zybKX7um+IB+bPiziAkRw51Q5XJAR
zYPCJ5i/36NPdjkL8JNbUS4sHU3FrVLK2JqwlXMpC20CfuIKKRD4PyAOR7BP/blc
P/DHSa6ExLo+AyPdSKjlg48qAEyYzx2hQaB3Xhjz0MUqQRv9/tgOKDGsOnFPq273
F6EadTpm799kaS/ImWjlG3Rg4f5xy0WPZTJEtPO7xNQVCW/2oiDpxIoiyoPrSFhW
G4bSFnScy6ijI5bCawD1Y8Rtb1cJW/AoFUhR1phcTK3kMm2+Bvt3D/C6mVPvS47t
npeX+aVHLjW3FZBo5Ci4BSyxAgnFHdQlOWFdhebiyqexAqpkvFzdTpyVKEAxDm3p
M1hYXHrrWhlYVghkbXgzcmuFjSWI9bf4aQprM38J1RPBHN6Fmw08gMgV6Z6W9pPD
umhlExBJiALG5pno28G+++p6G0o1EbK4XhQGU1YW1fO2Tqv/o4qp267b15SmOGwc
D/S9jLAVDVBEI6y6HU6Ww0fC+iSMj5N8nIQ35VLQoi6F4Wnk/NnpjMavnavvUMmV
1kXlnDzzGgruD8wVknmuR0r/MVSikv2EzOFuKve17iVrO38x8UYEPJYmTmW8l1s5
X88fddUWGlUQq5WpJGJz/Tz/jJW16QGIftjbiqG154WfgNua/0rys3eXdHu51o4k
UCGnaNp8wN91IniEEuQhNJPIdsRQ/3gurijn8827ojW/kvHGVksHz7Tfls39ir8t
vUdrjdrUcWnMz5se/Mx3QxLwN8TkoSuI9OXK4CvK5klxAff7s1fy4gnbJCqwPF9G
FvN/I6ajyKHspiAcixDqgBzSst4ygvlnQjNAfviEx2Ny92k0Bs/D7KbCFHGllZmu
gARHTm4zqrKHYbne8tKLTgCL+YVqcYRb4OnAimB9Xk42lUbBFr9vXW8FdNwlFwSH
4aKVuSatjzdZHBZyIfJiLNiZxDAHgl5/lUW2xIhsJ8tBG2/j63tBbn+1kP0T7U9U
A5+qm60zEf2TLSpTHFZHuwnEx8QS4Oy4pSPv12Uyu7xwR+AXN4hhl9vST+oDDZqk
A4JwLerMfX2adUCIwbhP66zKHZZU9Rf5K1rpmjuAGbVFEulBBvwvnW9BrcaU1W12
CiqkQQFekOuidi07yHUmHn+Ah+szKY8h85sFuRhQ0xswbaePjH4fM/48ioX5IR0r
IxAQo4mzw5kUArl9s38WjTBr9BW1c7Gv93f3zY9/dj1dUcSMbvZ1Flk0Y9lCZt5F
Xx7RLTC+K5x5y7CHhvjTlCe5T5WF+GdkFsZOC7R9UN5U2ePGofP+6l7VHZJMUzca
Vys8tbsXO3T6cHNaX/64O/natucYx7UI1ucE/3/KY0IxlTjEm80mq3GUFclGb774
2m2Gv6Hf+6DBzOQ1nOvQExxfnEPLnDPurW6ovzDdjzf2LElZjcAT8RAu54Wdubn9
YmIJIIsVdRuctdillu+dVKJNx92Gk7DPSOyAkqsQ7PfR74AzXLBpMBHuBdW2TMNL
7xCoWNbEGAaBTHR5r9InsB6TB5h6rm+VPc1MjfLa/UX0Uil/jDrK0XOVf+4MRRyj
2XHCrNvKvKlA3Tp3drvNXXOWL1W2QuI+8OhETMjNDr3CFsDurgV76VrnPMRxxQxl
T2zOz++8ShoL2xRQZ08c5JKYcbzWt1/tg4NrcMUpn60qeKupgWIVFMLPj+eL4FzJ
xWv1jnWwNcf4EvOYEUGFdcqsm+MO0SckHMjT0mmgPYhDqbctdnghf1haRY5oRyRh
rqAEkgnhNZuny04s0Pfm9nUw0teUCxCRa3Bv3anIZxjIFslWp/a4Aw8eDKMAbQKO
mlmeHH1A5VjwUf05+fLbJFE36WSYqNpZbTOBgcdubDUISIwvzrartRO80T5ZuJ0U
Yr2Uek229iQkT1U15+civyzUrbOhvUQX6/gDXgCPk+WdPizdlHa9tRMEsGK4E7dI
0JZx4Z8o4676I6/NTL0PLyCYR2PjYbPkiFMcXkdq9V1mxq7mUEdguSjxVuwdH4/A
utYJS3cDr3lXdrIkpAuuF+sHBN+YSbb+0SZShFFV3IJFD19RQvp1IQkcJXR8yBxX
VfLGpYkyqVr4yvTEKBE4ezo1M0bkBHZsLeaHeCKxtURRj7UzhwNHU2CuOZf4AIGZ
1jJs0sIEV3h5ACy5oHyot6qnETpzKVa1RdYII+QutFv0cc71pEjK6z7OMDiz4wtJ
5HfniCJX2wPmUEmeY4YKrJaQGh+Ynmz258PEUSwglbgyc+gGg+Ia1U/skh5uhzIh
XWyQh33c5NEhlUeNe5OrN41TkXQFAL06g3QpsORdjn1wR2+UpiuZ/6CYk3KBpMny
Why6XivhSwCSGxDNMKhfHiewXWZmP00sAE/L0sSWyCOpxXSSr8wVIc1sChQZ0UYL
oSvEncYgSL/mPX7lCsvt6SIkuzwNIA79j2z6+Obw0h3QGN9tCKwF3HI/wTNOYqqq
p1bRy6+L4A3wSWhwZr3aBNitAB4x1RaFpViffi3z3ADD/AQ8CWpAzqSXgvT0Rfm2
pVdmGC4X6SJ5nWy7bP3ifZjZlVcHrR8BUKttULHYqNtsum25W35fVuz1SVu9DF6R
Yt97NR4Z0+yNPNDrTkH+74dsDRs6CBVi3Fxic3My90EVe2FRHRaftYrBxo0NfBql
3gPCZQA2a+V+2uMu6c8Nf0e2Knk3nX5nk52tlq5gDMNd36+gQDqrFA7gg6tktvqf
+qKrMJkz65WL92Vdc/SzXQeBfQJIeEMsNczyMdQMazXl6jRQsns6RIqNa3oQ6rx3
ufjef9wmwfwBhDHqZnQtwKQQlalK14YLis+YRqXGvxgQV68s1sFnGvrInzJmhExx
xaVwyRtbNAmAFKq40tU3R/FYNvCI7dL3/rDPUJrOsh9q8DafTytxeopE2KDo6Ji1
Micnp8mnBAc5KFPyLzB8KMgozHzL3Cpdo/3O0pqm6bF+TBE9hqs7PGE/rJNQ0/FL
TFmzZQ3/uojSSrNeguoG5/9UIEO5L/i1CjanVcV2KAEBUL1N8luY2Zh/NCRxAp/E
XnU9df7aFhPcz1Fj1d/7L41LTfRaXm9CJ1fAFo2QXyNVspgt5pQziZR4eiwtqUqj
yP/HR1lRlhCTda1i2GFEalbvq8AfPBb0KDL4/2jXoVVXFKAIJ+TCBXaQJPAknK9Q
sogG0+HakHSnNl/9/slibhKU1+PV9u35DT1qLnK4xGkA9zGZ+jRksJpChVHW55eS
un4WuFiev1y1SOhTpchqLAAhZA6y64NVMewAlRG5b6qY5pI9qjRJJXpPTfOSJ8QP
eM6aupekZDwxYogXkd1EGsM9SLn/qx+1GW89LZY/xpTRqsfKRzZDzDJasomlD8r3
B3Re24A5kBfVc8KWzTYSle1ygLxR9iAGhENnpxo8RlIZqn43UUhLj8Q+VwN2ifBY
T0L9D/hetBvBvhQl1emvzPKBbCBu5zFQ9p9FvV0rv04LM1xK4DR/vBfW4xkEiMSL
zHLONbJbkrdI00oNu1S1HkfQXPB6d4cFiDfDOGE/E78Hu51mL+v6T3N18zeTfUR0
SSe/B/gAdkPTo8qmkdHsswyVr41n4tBeDascUFbgxGGxNo4fvFQxNInwIM+YC5j9
AZmZPhCbgGUlf1/Lk38yrrgg2FwsD0xYwEKPlqJ68ovc/BKpCXdCwFwXzRYT7wKz
tbHlQtq6e4f+C7jtzkDyRpTHe3HLnoXZ/5r9pH+dTx/LPYu8dmBR0CdX6pW2eonG
UlQhTfvR1xd647cKRECDuCzLSDr9kRpAB7msosiVFBPBSQwpyR7BzZKuKJQEKBqG
Svk1xSKgto+xfJLsKkp3ZHi4J7JfMCXaI8f3wYy6zwJQtRjIU07zf5aEsgaXGrHD
g8jzzoNAG5R4pU7mYIEDUfy/iimDcPtgoKej/Akakvf+uMtyJv0eGOGpu6dlbjdU
5ZaJEEvrlFuJtVZ8mrFnjz0XZlbMxxv/VcUE9uyT0Jdr0fxzscbztPcHFE1i1BhV
bhsaTKFCl5dUykbVENeOJlNJeYBv6TAVG2zeGEedkqcswaZsKjdF17M+oKuXpMat
gQq2rpATr0ve6lHEhZ7qHkaDYoDxoB2Sl8A7Tv3ozz+vwfK+hdBGAkqFFhxN7tmc
q/dzmMATyi+70RbgnE7OpbO3BbAORNPrFeu7L9U26VBFgPCwSRKCVlziRp+GF79+
282IXzGR9nJVJw7P9XTV8Upq5tfKJcs0PjukPdYXvEn1a8mNUug7b3x5DQnaq419
jCVY+igxnq1nBavQp+od6VfiW/nAwQeARYUSUWkL+b/Q+hdPZ8vY25ISh82/I7q1
fHg/vv/EYymhA8Qe5i9JYUGnIBrxmnRx9kCbiTx+mMyJ8wQeLuKZ14Mo91zyf1aA
3AWz2eL5UnyJAJ0zOAzM1EgFx7YsQ25cGF+5P2pzebpllNkETPx7U7T31YFjfuu2
iPtwwIiuvbbSKcD+myQyexTZ8mieuIvvS89OUEP5RvWhp4Zkmw86RNwbIhCG5zab
FuYlI0jMjQGJ1fPy4akE3qtzQ9nJeZJEpTu8j/gxHv7stiKAUgHDEfhZDl7R8hy6
o7dLDvVtCfi/bumnxo5MHHOKfHN2SIA4mEJzDQoofTwD5/xmbRiaWyUKYKjre9de
5www4WKKcey2lW2m/AB7ivsWSe1LjZmQ7lDX/sHw5Lq/DIlxtsn3ey1Pdxv91JIn
LK9pPhxtRlL6fy6Xzlz9wrQ5tIpcpHffqSsind/0FYgB+otaI6iVBR1Abp4hIbex
S3FPQpHybHzy6TLVBmH43IhVU8RHy8HbjXTjgeRPxtfUbNsTS5UdbZqHOPBVIpeV
yi4xCA9UfSZ1S3Db0LCFz1t+r2O63NQuhPRgKi7lMTtW7x0SJTkt3C0P4xatTA9f
MKmooqInJX/94dgf/4HoF6Qm8vJY0FFqCgfRUFFBkmIVUfjAMR5dsSWSgAuslz2v
2mpy4XMkEJISppgqi3pkwxQGp0F5evPS4Z4npvcqneYPEYD5URhW44hIuJgKkCM/
qwRg3yp3wPVWc0fefr5nE85+Rv5kTSq9IA55uKYkL1hbKFSbbKoWZdOLX0mQlLYs
42tyGw4Y7n1jXW3W0p4B5MY9TlevCnp0se7KTQxIgiqwBfNlMjRhd+TigP1rzjgD
AUI6cfF8TCsyJ66oMi9ZTcoTvYbcMF4e8D6whlgwPFMw0B9IlTL3YXJH5ykBOQoX
uEwualxTb85UkDX8P72Ym1+lox5eHxsLtBGUgUu36X1m0Y23BX54znjGgNdGK1UB
UIAWIikCzICODLisUAu/R1A4LTOf/L7VAwW4DzNu194F3QLgLlyteL+v2vWRsCrV
zR+WRD2jUkZcTQekCmIcB9fg/CLFjB0w0pJNrgVnN2OF33P3ybE4HCN4jwAfFMy9
Ju1jykmtFgMngA5rpF6FlTIsh845jkjREQ0zZyy2FxI/FIFkNKaLTq2sGZaRu9mw
Ik6eYmMrsWsXU01nsf1CqXcC+QSObEtQLF5xzVlK5n9CphcnA2klrBrP6WMO1lV+
pfP86VTxkKSlJMi8Mw5hzTQv2FaBttFkOPBT1qMF8nCp6JiF6WgtC0ZhdFefkZAb
hwLGalTlTCTjLmzvsInT8l7YohKx4DCoDn+eTi9FaWn+lO0pqJ7PIRNXwmICKWBC
vG9af/W9wL+8eYk3rWf3qLHtQ6CRNiyS300Myi3yEU/Ye4AdrDjDLLo1T3yVozVs
35iNPzK+KYt44Nvb4lbSOq5gAu6MdfaOfyqW8Rz7IIoQm1upaYLca0Jq4hjLh6Yj
V3VEoS1xXuzkqDx5klC+k4qgk7Me+A5wpypLVD1pzktZZ5FXNDPAFC1EGEAuU67v
FNF8LKrciIyIyE2DlkkK8Ex9AoC5fma+nkukg4NVospOP/j4q1bVY+chuvb6tYVM
LJ34+iNNJB3iJrrO8pvKPC0n2lBzwdcm6UJrv7od7p13yLBehiuUXWINuEhXMIR5
rpHuvY8+JRwyMaAmq9Ve2dgmterDhhPvgPxb53GjstRSEbZbW+aKLJblaAgVYOz7
p4UhumRx6wCQKpmx6vuNMb+qfZ+gbh7RxPjvFTgyRKvxeTVvGizQpvxbGoUeDlgJ
0mdU9WJJUoz9kZsAkEVJuqJOYDFGH6QYtoL/XbHkJ11Uuaqp7U963WXgYOEby0wr
l6FfEwy5TrbuRsBYVcIwHv4v5qYtnHKlWtu1t9Jtjh1rcToUYj+agy4Gmqg2QB/A
BvAo40yzC4OUwpX83Txc82VtGR3mrgQl1OIyTN9rylQKuCKD1mLg3Zjo82ctR1hD
V4+B7xXcVDpNq/yg5THOGrR6NL2OB1z2vHFKmlLTKZLu0M/TtR+nF+gEchBh5k3B
q90Xnsj2Gfak7BFTaXmjPsR6kCqLtnamONRjh5nVf6tEKf7qoQhhdGX06XOITXE5
njtR+Ua9/C0LdzA2+yQ07ll37POAtrWATch81Hte+x4Ln9ahmyES3MGRoLI+fLnG
1mAJtr0n2CpI01ktuLNi/znmZD+M85Utih2USJH5opYgxKa0oIxm9jDrUGGXGYvu
ieOiol9/auWpXsm5IQV06a74b7YqGpuV9nsrSEx0EpH9SnsInMz/R9TZvV8EAodQ
0TdMOjISJmDpMDk58SjRNUYdAvOA5QXQtmrOx003h0TK2qlBZePsUUhybOH09PHy
CqhBn0dHae/ANz/Ge/QcTSdhtRxl32aW1FrXGSqxDJ/vj4wYGp1Fy/I/IkufzU5P
SDI45e+UWIo3zDqqI3dndAMdT+446l+52TIYoD7lQ7IPjhY3W2CGfH1DS5cq1ii1
m7A3XHs3xr0qy6ASrDGvHTGanJQYD/v9W4hU6uP4BKqCrmw35ZgscXTkA4pGzDhq
9g6cPJBopfsJM1Kl/XzWAtnR57VIHZvmCahm4NWGIIXJaTRjSsvMCqjqdks4NBCZ
Bf4aE4cwiEpCtz3iJT6StVREFbsyuBXiVGgnTVs3lQErpLyB2+SK2B4sk3nm3FMq
zFx8xFi3I+PCgSDjtmJqvrWtx7ZqxnCY3OQmcfA2Uv0B37Uf00A5beT1ENNxW6nm
M4TyrCiy6STZdiSXD66gAqI6Mw0yCnQYS0VNCZ+IOt4CJSOLnWdC0fGuRmCuqV73
5XdKk5MUcqc2Y3/14bwv5t2jwc6gxZJljVqhqZzmxf6qZiEG89illUo5aqG7teOd
II2qMdpIHCjQLp3kf1fYgodE+a2Qx59EXM6hm2X47SpOIi6ILtAr5/QcoXCGcPxw
WV7kimPsZJ0hcst1zrU9HNvzl+k1mcJ8d1q6qFofVl+pnMOWBv8RT+Mp79Z9tBWM
xUTPrM03qPHLy8waf00JvgfAmCP+Ik1IWwu33H3n2K5Uh3lEIU4wOkJWf2W7avsY
Ar1Ct6seaob8rzXpM4XhB6f7usJj9aCFJYJakMniv4fvvWy9PcHcWJu7OV4DiPXh
ZqmLV4gaOz5JEHpH9Q3Mxx1eg3N4/bHHasXITxJmnj3p/j4b8e22qxp3LJsWTLgM
77u0meju+8pSLyhh0NW+4gKmvdy3L+d0Vn2OB5QKmAcOqmErPjOi87vPD7RNQddG
r607fpdZJnIYlUxR2kXmGRZhoDTROPQysFGEqEZF7Xf4QVTF5RmBxLxEIASjJYRD
eCeytjwqjNMjH4yNhd5DyMX3qG95Jn1kl89JGGixlnZb4486itClNCGZhij1Eafy
y4xwyj0yR6jtPm2iNbeNUf+YrNxE7U8ifL6Son7q7sgxf31NzdKxIwb3ZMl3yo5F
9YUytYsvRkYCnG4NikC2tI6wFsGlPJi2GS/71D3IgdAS3kuVwrf+9CsHSekyfb9S
R9pyTXgnfON9K5KblciwGo3kUOkyOMR9xQ9B6NAD5/sXaQXX0XDjTcnVcXg+DbUF
LsLXNKsd//gnHeP/Uenai1DEFg6uOZ03BY3d1Os4q0+t9G2jv1lS/2F6qoGCctEh
O0hQcRLbrhZhGhPzZR9bT9NQSoEtFkwB5tDPZ5nDOyVm8AN4LytJL5IPMxNaEzX6
FGAsEhtsJ29F06s3XvY6C6QXhsow0NKdSe6TeXYmf4J5uELvvEmDsLkpUqXf+ZYi
E01fm7ALMEc5/IdhAkBfaTkNjZ0HNyR9ThAbOP8c/gsp4NzcFjEMg0lVnr3ePCsa
Ydpl9TwcxRViMsrf7t4kttNCydt38XDUgSabNaSz6px04Yqxb6QSNzLo2Db4CaHu
O8hD86LcMHFrCX9AG6LD8BSOYNRDOC8MwYgCcIC/9bm+42MTPP2OOarXg+891zKO
GB2i15T9fyVv5GJO+9w3E17E5jTjpfcps+W55Sk7VVW/RcTwL9nh+g/7gYoOtNJt
5dhFIMXDOMPm96utcH08PukgeUJHfaKDRNHRKelQtepubzodAOyRCC+OLKsN4DEG
kbVIukZ7k3nYUWTje+ZJuz4BDF9ESZHDw/LeUVJjv/peb3mcw5/Ezj99QNxVlb3H
M8xBc1/cqGZnVngYtYm8/xm0ahu7eFHsYzuH15ZndVHMwojj/+CN7kLTQip1BJjv
uCcnX7T1VJmEpeisVIyQSge08O3B4xiGFJD9qQskHx18e8j7sO1cUJ1nfJ3A/B+5
3S3bMiwkzuTEtZJXCTdbBmFecx6FYlExOdZ8xNRHWpNEKyuQOMtm+fIyS0jshS5A
E3wQie2Tt9LgwQVariZnY2STUh3IOE0ASVO+iiOlMzGDLmqR7GaUSR3ECIdMc7zi
KhIqkyYkaxJO0CH7KHrHBKa7QT30vv8sjVCnjmK/wWmDaxGURC43N28fN+846VZo
HD7fmors2KutMyi6EIwjrR+uVtd/eRtFZX/0HrkeKZueH/LZTxH5elvnRgepkAQX
wa1rPWyecw67c2k07/CCA9iJfUUvL37WkBZ8s86jIdhhQJzw7UxORnblzCxGs5t1
m96noniXUXtklDjlGj4FTyTDhmtq4lNtU6QbPflYlzbWP2//c5SH8Jme2NQXfAKn
9EIFCGfwGBNOpFtG/s13+LTVtR/r9Fy3Ov8wCuI0cofmeayS/NLgut856UJaeIGS
+jq/NRy9BS9p4NelYWB4sR5ix3TmNMJkhl0PO6cb3AQ1j+DzGNFuxuEAu9+wHYrc
JqkY9xrrFYhiWORXeh5d4ntMH1oQHZ65NdSkpRQJaZNpP81y4zY8gbhClRz8jFdO
e1xQxZibIJW88znlMqD4qfdgCUSupZFg9TCK+IX+ZPGsx2vk0vE5g8IFU2++oeba
WtlT6x3rg55yq26z8x+9FsREZ2WB8gvymlMne64wVvz57PdkODzfQU8qbkTW/NlK
ecTIJWNDoatm/h5wPIJy65MvCNc3hYy5dG0Q9Vde6AsO6duVSnKTYG2SGlMxK6vS
Bxwrg+8qWSBCZuZ1PVkT5bUsWXJ87ZQ+bWXsjfqH6Ief+Ig3ymoY2SlbeEY4iL+f
v9oKftxV/5N/9jTvLf95/UwvF1AKLd/OCtiRNGZ7Gf9hczC+ta7GKqqbkfWUQMAe
ZF9xUDdFSD7lLMpPtCqBWCH1YMBfCc8qYdEWnC+QX6JmQgmF7OjIn8VVLeQ+8Y12
rlj69khmcAOgIzDxtX37LfM4gRXhn2ScVmJQxm+ufLod7pywc47TiUK/nIDQ0IPW
zUcS7Jm1Xnh+GfRGxWe/+hWpHp/IfXMVP6k/An+OY889M0GBgn9VLkhaSmxLrsyx
J73IGLcStx6GRwsUkIjjzrxnvMxOsyEkZZal5twM+wN5LU8x1WZH7CaSfGL5aB5c
EHiOtT+0HrIf6wOU7cIPexB46QRwAye+gtshi6P7vHwxrkToEgohfH5RPqlRrLb0
LZm6fhw0g3E8uAPuRQix3AnG6dueWcT+tXzsawbrAGIUZrotcW4X/JG0KdomPUGm
3AxyFHG4mPwqzF+emz/RX4Tdb+6T/b4HH5jrrbFX7jg3ksejr1NRDxW7Jex7qHLZ
2qYropetXQ+zmU1mGSGgHd/JZaN92d+tS73FHCUTHfU6WekU/zaoJSAlQZdxKdVn
+LrATSqHtHsP5PPwd431SouS/Ck5avKPJPtWrnpnNGvhizZVJHC8teGmkkhhKPGn
yMZ47SD/oWUQG9xxk1iEsCT9GMMORmNU5IjlraCIpFLr0LAQTJ+/ZzPyDnNVCRwK
p2BUuQhsb8URbDFg/fl70PoohMvHyxID1UzlnOqw+EnO8TMqrgsQzxtzqpNkxBUa
hGWUt2armxS1kM3bV6qwQn2cc+hxWfGJKkPWfqcuGHLBFTqewDdvdyXmSuaCnwt1
BG885CqZ2tMc49bI6kS9B2xnoqeh5glT4CTnDaDrMDP4BwtLR5aL+vHKKK6QlWAB
HgstnNPQcs5oxtOrdmRY//CNb1GUujveAkHDHBeRCum5bi1ECisRHMWipXt8S1kJ
bIBZT8tAUPLl04yng/1BAFc5gNzVV+NdWArf8phnj1rA5MviSom8RINM4LFC09iD
5+08sYia1xttZmLgN80cWMJGAYDkA2yUjXjXetCNCq161Q7MLlOe2KE/8IjqGj8o
mJAJEQNuYut6buqCR9LbPwQi5LARc//Y9bEz82C2QpFQX5rL8rG8ZD7vKb5ifpQx
D4kfJH34s2wdcNHiWFjl1dN5OtoXh/L1tillO6kk/U+Kf4+6LQ0qPqolCilocOsZ
WY68LJnW8GjL5/qy5zCanXaemHRx2PFz0r47C6MW1iGENPhEXdEumkk7YzDoH5Sq
iBsCIGtDCmmTvGyTky5Xs1R4bDcFd/rtEijl+C5snxZkK4sDPLThnbCxf6y5ftfY
1bIiU2H00HSd+ZOGTSvJ/RJOpgVeFi7m6A0sFq+il9+A8a4xth3ns8jjKQqkYdzx
X78Zs8et4BqZ+O6ThMsdVk0HQ/F6JvTKc41uh6GmRcKZTIVOSKU+Mo7DAjAP0HUq
HjNiVFvFpapwRY24WWjAk23VJrywZdWhp7g4h8fcpzNcVdjIUFC3df/hhk/5gs1/
QmPLlbz2lA+BaYhwwlR+anZR9xdHCukiU0o7b9BS51ze5M5SIFw2QxEuFczkw0ZV
j3l70fpz3oiqBTKZ1V7cttLPYwR//tSQ3YUbTQpdcdCjKnqLktMZ+VEaKAauS/PK
s8kNsxOxoVkNPbAEHrlWgKGiTUfJarAc1OkNmNRuJ4+xGWbRKq+ZlnozE0sg+dqd
GjXA8AjOVcV4kxvxqK6GiD1ysJxRwv4MMTWhDERtlga1Xx16MXs29WIbP/69mXhq
udddcGZ86z6pfoHtu2vAASNLiKMnTDTzsikel/xyCd6dZ3tivcIwlAXFOK6ZYOBf
BeyxVBaKX1bwoZZbbpSnNOd0JhgSTPEpbs3nmma1vw+o8x6FbIAA0zQFyqU4epy5
FvdlfbetGQAREgPxczW73aLp3FysUmrgvCa5laUvy5XfVpFJCbLpypnx61QSFJCo
XIN7+ucJ26ZabnbF/suCAHXikRmNCY/hFPCcswSueaaPQPCYRYp4Rw6oJ3F5Fbqs
B+sevAp/H7CRvvQ6bJHqrlbCX6VBKY7hlaQjuO+VZZHegECByj5IQ3PXjkpcqBXZ
ot521tbp3xEaukzx+oTlMJdo+WSM/Joejgn0xb2SXmf9N2zYFZGewdMf7ImciWcL
+h85M4YKdh78OgQN78IBcgc3e04MeNLGzKlESYEwuj/l/Wxr7lD3UX97Nukf9G8U
rWnrENHRhUOJYDVCXJ9gotBaNQWgVfvBUQfNUMEmV+Xwzb5D/5+0ch76YFSV+YDr
JuB8aWBl5zk1bKKx9lkKHlJwMBC0/pAgfYGzlriVRTRykJEgPFampb2jfjvCc6NH
8WVS16jSmEa0dzLnTraimRbwlWjYfK4s4gJTCfKeF8Yz52Kpy4eweSutKhJlJLln
PUaPHPQYRIQ3TtmBAdnlgBAPkKnLPUqaoU99QrJ5HFUL8a6C3JidjCRLYPaVYbEz
C3roRKoOY/swcfoKEmH5BnRuHmhAUuY1dLOYV7E6eE4QeNoTZSsWn809SBllP7Xl
CQbuSpr8ka4aZk1bO0LIl6Rt57Cr0GwcLQqciQzzsW+Etl42TAGpIPhdn7s1p3f0
FL+qvkbIsB0cgUgIq23/e71dKhTQMy0wrsFXhn+/1EIkZHfLjo86ij1FsMzu9aPU
kcHtjLK9rPGkz/uvWSWKKLld1Vi0gpXuGm6tYEAVsYI/26d7sUqqSZcWHZ+90ig6
rehkwsyuVpZTCqs/fyQq3dIbqwB1keNB78jyA2juwY78xliDXTcoeXh+zh1Vc6Sl
Z85CiTKdLqF4ZvNbBYSV/o5aW0Vyv84hh5ub45lovTv4HwUrr0y/o1CZPgh0Cf0k
gC7dFZXC4RxEstxFJqXfypdV5I1U+XnAxMtXYpMCie8Z1QyFUoUXyavrAZ7DHlLs
8SmClttK2LDgOUymXxKeBWBjgdAovUUsLfWYp2eec+1l4M2W9TR6azHU4L5gw3SU
AS4T2Gwt/JoBcVQEKhWB/r8hHs2s6xMvL73Djxg+7QEDSo6hJPD5SSjTUhUNr2/z
Ic5dQrQWGhpqP+jNGHCsu6aXNYV9sXjIEDwM1cGgjo6IaMIPBe+tMZh2Lx6ajAfK
NaDXJGvyqYPsnCRD25IqHZUujvvEFfe3ZTn/NfITIGgjqbdagwMACCIHVSR7IiUQ
0k5z5C3sDA8AhStn/fzgkc4IGp5Qsc2EV+kZCMXOhyUv/HN8+RyXI/mv2iX/lsZ+
7/alyenGsz14CDKvrG1L73+KMwKeXMxw9oQaS6zA7sGcFI4LU8CfK7LBe3FO/qHR
VI8fxvP1q4zB4YxVJTCjWnqS/yIFA29xQzoCgch/98OPjjMjaBbcDtUuuS7JVyaU
Tx6vcxDNHfWKZxUQtQ9O6EslF/N7CsRZDXeaJlDHUqz8ztZMBH2abo6kr3dxwm22
nGmAV+Jr7O4FS1uFIhGnbQs1zjEJrbVOihPrm/LyTShhrP9zIf2QmNEU/jxoBbHC
Aynh/9nYxO/umHFpwcoumXGLumHvDR2jIcD3SiBAYqQejUNhk4A+CXeHOJmr0Pk+
FTnGXLPB/+F2YxjRA0mJ+ZADWu5tIN6sPJasHVXt8dDJn6+3DjVO+VxnJ38vQRKp
+wsnzHomWQdee45zXdXqgDOVW1ZfhQ8HFvBWhzniMuMRf3jIWhKfEbRP5pdKt601
1U3GeQ9n/+QmIfhNki1hyjSz3PR8LD+YAMkdABD3s2PYMDdq4bn6gDuq34y/zNdh
yoeRiE6TTbUlDIyz37+0rIm8lrrEJtnKr8+kTD17/TGaIpCTBspSiHdwbODl3OyT
UQ5RO5YuTwXfTqJFaT6j1/lhlRLxOXG3Y7rzjpJ/hNDfQXW0U8MlWJNqS8PmrsZb
dSFxptL4POUqAh+6tMQtLT+jM1hAGVuBTZFAyPr+vGYznlewkdRLqSgJ4nn5lNer
eWQPV4wy4/3TijxW9+9H6qiN4oI7KA1TDhurEd6amHHYz66kGW/clqWViqTcZGMG
TDpWr1gndd7355YbBU9md6sBeZCjCZqFhFfjWJayAuhnfpzTaA4Jt92pbDao8rvs
WrM+oDlpz0RP/CUo6j3c4YYGyEacB0voJHa0dYs9+61yl0TR5Tfrukl8Eb4byRQn
67enCQvRupMbxJQew/Xpa5OrG+/ykS8Jx72uUGWxW+qiQgLvdT3Xc3MQkbzRSbxt
ggEIQm+62r/vF//35Ho6DTtFLB1g29yQMpquDZpD1WiVfqmD42perQDkB90T7ukk
mJ52KLH4ZKcGWyN4rkwKRJvpeTvnYK60vyGs9pX9oqWccs65N3UhcAq+N57iOxzR
v7RS5mAZcUwWQRAF3f6Q+IiS8psoL+Zds3QMZn4mY1sHqqP+c/jZ/jAyTt6ITH1t
DkAZKg6urierRSFLxB/ZzImpJ4yuEGUtJvJFJhfwXPQKIS0Dx+sjlBeXr2j9M1V0
kwo5m/Lz7rNw5ky5Tj8YzTOcHwn1i0RWlMlQ43mPxSXRKUqPquohVNO2ZbtbTZut
DXmVk6gNQvRMOIKb5OaIOUpkkx5T54ZZkj++kAEl9Ph+259rEnnOA8k7YV4k5rms
inoVhYsyrHr/ysofYhVzC2mLCqfN4nRGU5WtevTUSVrPzEAJw9Gl++x5Sq289dyg
AW1Fl3z8iGycZ9GDrsRiqh4vJfStfY/70fFpKDAgbt6NCmmejYsAYfSXo1+bXqe2
h7iLA2lAWNNpmC2uIGvOT2VEhzvQ9bMAiCVqfosdW48Dhd7zsob3Nq0c5yVzFA3S
IkN+OPe3PrwAr8C3idE9MuyEOwX2Ezxg0jzjyN3i1fY33Dh9s2D/g/Yrv1DdRsWz
lm/1a5SGCflOtqD/1knIAlcAqrprEt7aG8TR4ctFfsI2VIyjQ5/OhB1MiP8LhOMF
ge1WLA/+UgZ+wJbWvMs6ZW6AZKVqPQp9hq/qlLT/VqKy63Vn1HPzLD+BjWSBAKc7
EGGBQ8f2t//CFw5Ys3dec8L9Y1USFNkAhuLuyXdm+d1H2/esM6iI3ROxVG+s/Q+R
knQM7HfqT9bpO8wjwccxYqNNogFMqswAfMwchGBzA1fboo5swCSOLmhXXwufbtV7
AdiwCVtWGCGH2eE3BO8R/HcNXxvzuwL+3RcJAn2a6Ao4Q1tIrVX3tGcSEb/j7Xjo
Qii86o/UEf51/e3psqKg+EdvZdvNTpt/pGtq6PxjOWDIMEyN1hvjEBDVFk0Kb1J7
QQXcrc9Dm/jAjsOF/01bCTm8n21uSL9OENG+WQwtKCPDLKXyzuM4bBGqlZB1ZeVd
hPA28RVoaQFzYfoMcsj9Dt+N3Zrf63+avjMFeagCRGloWF+bMlm/m3nV7Cpbtld5
WGllaImGeJpwPyQTw/DZtb5bp0BufeGGz42o+7fLJcAhYXdJ0HSFIUq/rhcJcA+y
/W5YM9I4wNaw/P6D0whC7ExlcKhiMtPZGm2VTqkG7p/cXolpoSnzxlnWRnr/4uJz
oHhcynsJyJ/GQWZ09/FyZwRO1bIWBty0OHRbvlV4QdaTThSMlJxtbUbspbATlLfj
xD32xOHhq3/6YKG2b3ZpWOu4p2cxTAuQRTBfa2rttCoFa8gH4H1vE2qLRXXM7B90
2Cbxf2uKmRxcUPzs3g9sjmVr0Up6/HOUzjR9iszWrlXZufTjEQ8Adjt6p/cybWFw
fLiPmSQWr/exf1R+yca5skMQ45hx657yl1zfPf1iSuNM8wGtjrOfptKzV0es9yY7
heDXtmOXUtZkDJzNUNwiqTcJXAJYv5MVuZyaq8g9yI+ZgFfJwHmK/I2Dy9Z+egW8
RxzIGLuSUOgPt5tnKFDXaMhSnmr8jAz581mgyUEMmAwNKjGCMXYIoPsOeei1N/bS
cUnFAFqCQikRhDKhmQTQHiQa8MxqUIIYMUa5nO0+eHZy0fu6o3MZ9R9vBBvQTemX
UCDLYNTgfmXUEO/m8xa5ZJ04hrC8Mvm3HkxSwi5MfEDhcpSXw4X/nXAGy+6sIm34
ja5UaDU6ncxX4oQEhaHFs2ZEyLlv/eyB3YQbmSqUX7udAUGJHp2RGObEVNMsvZzm
Q2luG2BDDYrM2aN4nxQX8XoKnfNDZzxvC0WoBZuZ4XKDtRhZh309Hscchgc+FOZH
YpV0LQwM963XNnefzAnuw7MEwbo8XBHwgewQu/6SrFqk5QUNgUCIOf7yOHfdNBtc
h3c+89hR+VYuZR4G4T4mlCSRyn5R4HwApEhU4Co5I1PEh8/NI0if7iJaLhmLyT5f
tR5485HoshJmfWrjZAdUZBBzg940u6d/vE4flbN28P3g4gqADXjxM3HzRJTO0mJ2
HrUx7bu5p6Clzuoo807NHgbrgZr15AAz1MBfGE96x1VWwtLT4uJehKrDyNe3F7C5
L6YAl2nhrO1OzBsoFSqY2/uVIKkQqVcVt90o/nMIgLDptPah/wCCt6y0Bs4nD6n3
6j62vkyn1jNw5oSiz9hRI1jmwF3pgHjyViR88YjmBCvXZqJPkwNDu6C8LI9mLTFk
Hu5bj3yfpr6RpyNpWFB947CTbB4Jr9Gukws/OpUXHrG0h/CWDdo7qIg0EVCwcetC
Q68yi2qsuy6frbZKk8KjSdDrGVOJFHFieuJtHmIvStos7X/YjC8T3kzTl928hQri
CbLWaC4H8UpteouzZB+nKVAZkhXRKdytM0/WKeoLVOaTmFYDfq5UxMwToUr5E0PZ
Py9lSpoeHAdgz8aIFifky5Gu9jna31PrhFexJVPvmixsMZ1qa1yUCHz93a27H4i4
PXwaxDaLRAn/verm/1Y+lkGUDfbF+h9iVZkXBnCW8OMsuwROEEekbMEUkniRUMwe
FLA8Aq7kBoiSGZHGqA0uRlsJkF/05MlNPOqeBRf4OQTOg+wYA7XrpqSDpGdXZGxB
lVWx0pVK5G8YlXWLumEkQvQ5F7n6f7lmJe5YI6zjCCr8yg67Ya11h9kvEg8PusLj
3LobfEHLa3lM4gfDqV18h8hBLetIFOFl6Wi5uSslTmvkOwV6bbGC/sOTK/lcEz6l
g4Ms9yjO8+99fwrNCeNAG/fS23iPb82WWwj/Who/t47zFjZcu82am9TEzvHEx47O
U374eQDsAyQ9i2mJB43pJK8PwUZIwlsXNOrFFGvS8iP623V3s8499VHRHHtuPpcA
b27mX2/m3uPlP88LM5EHGhsakU1MzkFgrbh0KsZdxxR7yVP7uML9ZW+lRWrSdY6y
DcmQzM9bpd4XG/44yj+xuV5btosk3hzgrtHic1DB9u+VKcgHm3h+Ny63u9+r774O
4BJov07hHmN9xmxxo5SJgdJiNoXK4hT8949OYy5M1u3eXRi9dpUIxgO4c2x2f0fZ
MKqORP9bL/Q74bFP/sHJYn0ShomylJag9vzslZaKVCcMCpM/6Zy83InfbvLOo/5G
/+3bsfAtoPBspqrjJ6Tdae/CTONoZofHqYq/lQddtDb30t3kvzqWiAkB0mAAUUrj
Kgs1In77lRQufL+7/igN2sukjvIr6YmJamIRPzX2MEWSAyiJU/HdoYfG27Bz0nfJ
NPbA06DU3S7v3gu01icElXdTmO2H+46qLeWypiFkhshorKftZuqA918Zf6kkNyp4
n1ZyWJfpJIv6QAAvkXOeuv4DpGosxNozNJ0klLujHIaJx5Lkyb4HS+kTR31jWzCq
wSyI6ShK4WS8gZRjEwlywHz/b0Vm36SXW3xzSu80RwC17Bm+CVUsmoAMCo7lnoU2
I5rwVirTYIA5Dgg8ZeYl+piVnaeHJHAzm0FzXkPiWS9HXZCu/wtgaQsccjRB2RH9
M9xuQmshWFueLnFQDTcTLaSwD/8f5OV8jV+R0iqRADqMFVXm48Yuv/mE7+YjUEUu
vZ0xI01qDTciNTBh/g1x3j1vKNg+WsoATBsFnACtzk8LMv1qsYKujW5SS/fiBGrk
ttcTDJIR5c14e/10aLHg6so0HwCkgxoPo600iqq8pTvPhBQWJxE5n1q/dpjw/3L1
NVXZk4oKAtWNjvM7CK2Yp5mWJww1yUBtftXaX/rIiSW2jfcVnMnH1SaS6bWtmrrp
14MVY+X3e+sIPwibSBR78me5b0lJjSFzCKNbRypBbAz9OxIGbJn6paF3IrXMlUMo
QXzPVQeszFHAsRwUehJJOsQjAu1B3oNG+iHhaQJ5DzMIChL4KrJDEfpWouLyFVSd
UkCKpQg7CkcLBGKDeXBUA4UAxt7rchevBZKYZwBtyYGwDY0SWHGfR2vjVbW4kTjJ
zK5BiiqjOikkzVNHbQxbON/kLfCLiggg+Yz2ZhRkTDEpN+9u3m5jxdkcxbLafYqa
en6fyKtj4RC8wdvjSO7RD85G4KN/N8iNsstrembs55lmHTmmMXbo6l1sR1CqSuNm
wp9Q2LPKb/CTY9v24fnXfjBiTnZu7YEMNoydogpvVzuWvbezo5+MNsz7WAzLJz1c
MQxxYlGEdDJx02FGAh10LIweEGb4wTHbwkjNqR2ZoPd/LK59m8do748HZtj+IHGP
c84tsTYnOBbEDO013tc8fRrzWwvPUtOEfJmG4oDvy338BynbQKoGWAhbiO7HyViu
NnxPjsFjcHJbrB8fmFqNWg42YpWigdsYW7wWwI0kRVIh2LvhI9WP6DmtMRlKA1Ay
RzE1li7vUPEuSH4a5ESkDTOxHva2naA7EFxVzJJFrfJWVovG8L0UFW51FBgGTK/3
XH/HPxXJssV/Srbs125RB0kyg93fdBoKOVRB2Jyb9dspDFkZVTpuqvqBPhJQ21At
N7FsQgYGZe+PpvrkUmWryY8Y6RZoj1dUYMNr1igBPwq44DkxRNS5UYKCnaskAqGc
STcUQyd3NpDa9sNdrhI21WFwyBBldKkKKR/EPWo/TN3Mbc3jgPZGycTylR7HFoV0
9rSeBWoT65NIpA7GZhlNU+BeOKLvCs7VFwrLT3goxX5+Z83UzgFNhfoTfZYAJq0T
SCe1iw+W54sGPi1leG3Yz8fZBxCzAkf+ZYfD5QUco8noqAmKpo9qM9oEqUosrmRq
AjNnPrTAPbgbFCPRkmlODWxdR0X8UX/y+0CT1rUWnx7EfObZgz2857bf5ItCOHew
t6TMeAbh4RSHKOVGiYFxWDCqHD17LlNkJQCY7Uh42tbo7ulq4jFbExJn6BMv/KnL
sz6qbxZrgdVlPQELeA1u9ATK7X/zqyPPSRqYFJe+XVvocHTogkcSBWOczi0bLNMp
WRznx78b9XPOf57ZwXjf38ddw7YaON6/kqI0JB6JiXyTYgFe4sX6iD3GQ9AFgsPy
yq6AFcitB0pbolVw0JhDry1f9Gw0jm2gFzvWC8jLDa5bz1zc3gDL9/QivnYsbcoG
O5dYbvWl8yEniRMr4DRZ+JWnYakcTnZ6r3VY3xzqxEAp+5yP6fJJ4c1tPcDdBpuj
ZQo/wpsKSY5rd3YJllJU1lY82l9lowYVuhAvUCfyZRp3lVU+Ai0yPn8lJYRIJPeU
dKNGeE5g6ViXKQf7bfCGDSYgVqJSa8CsWheRaB6niUv4b77lOxzAbymduEe+iczU
/lOQXnqqQmJZmYLcsXdWEi1baCwteOW65yR8wI+y8E9mU60q9W44G3b7dnb8/kmR
NoRA3byR3jzFcvA6JgkQCFzjQtKuxjzXFzfl/rTvJLH7PYYZmLBi7Uqfm+0y9yxP
07cpLxawJwAj2soH7XNIoHylwtqMSbPq+ZAxYx/tHG7MSiK0MFiXKxtHzg2jKXyU
txiS/9C5eNUusk7al4jVP8cDzXfkj/atvKUvbBFJSZOQ5HxY+LBq/VYlyMs7HldX
IizwSbNro0LuIUqs3bQl57ce6/jVOz/Cs1RIzW/YfPLu1NtuY5Pq5y8Q3DjuJns0
aSa8UV4Njwi9UnvKRBV8ekoDK8KqsT26OPAZKgyewdLdKE4ucJ5MVOKHiJLobRP8
qRk4ZJHd1iI/nGiGesKVZHZrlCEiarcZ7UtGJtCB7i7hHcCfuSemFF8jqd4ZoiJJ
ekG2wUcso8h99RxLiG+/ZERu/FeCIGa/V9eJp1HBZyBUxLls+Gh/r3BBZ26zIccQ
OV4ejo+WFFGiZVjNPr7R3BnaQKLjVhoEc4wvdQXd/OyjMAcj2eK9cPH80WSDgPnJ
X4Xo6gfSkob2GbFBP1CbtGbvdwIbkhP1eOcmzWqXafdScEX5wUNplO/HPMNGts0I
vhWV4TGju/Aqy+1Gwbak7KOPLWrR05kUTGPDW9ME/ZDzGFfswpigA/Pe88AHw0d0
hg93WLl0Ipp3CZLvKbUH0Eb4qKEMczu4V2wVtxZHAgAet6G9w/i2GF7wfcAoRsWu
1pCz7km65nBIYdsULeoWAJrRsXAxEcYMIR+fzoHb4u1NP7omA3WuQ7tw9B9HIL2X
nr+4RAnsbnxRnu/5wBqQrUQc7jasdTVFMfTUZynM9yY37jSP8+8VKhdaXPW/pElu
rch/gBu75kD0fDkxfOjItBShhW4udTF8X8DouUmWPHmIDKstyVIwcodaHBXtsany
3JrRxqcZ61Tj595BwQMKX8C3JK3UMzh0N/YoYkWIvws0yQrdImRiT0kNrksdn27j
qb4dWMiM429EioP3Q47W/gwuCzL+jlG+eI9G31HGf2Vmh5bxbmkT3kvAnjYM2yPR
G+IZwVOWgZy6B0RtzsshbnOiaGSUq0sQxLhWlrRGxRCjJQla9jwcsATlzcsyL3By
g/Cb1dOkOA+jodveL2t3hzxMXSrYC53Rmk2Kotq343yAfYvoD7Vv6KZwRdwr8e37
Sv2+Fsdifpsdt6KHYSgWXY5hxe5Xk5DbGueiL6iTb1s6moDN+I9ARLyLQpGj2TQk
EiqWHmbJMSVQezDXi3M8JKR0wayJBlrV1N5MAvYvMe7ug5QS1THtQ0echQ/5eNwW
LwVzTXxzC6VZ1gGPcxJ1YH7Jj23UqVlSrbDBiP8/QBbDL+uTZGVafoKdj100leBq
OZ0wMl0h5v5iSN1rpfcjFAuDLot0E8t9cfs8lXaQdqb+mfkJ+oQM581O0SCDafip
s6LTOvOMkWYyOPBCIULknCE8SWSy/PwfFKJGE3MtJxlu8sc0Dm2ej5QdcCDVVPbc
LThYHZOS6MdQZPJqdOQPkiP2xXlDiT8Q6RK/kG28Vi4w1aMEaGt+HBOOK1DrRPV8
2X3UJOP8cSs/KB+UYo4YjXA6nY19r6whnXcBYisePBKc3exkjcaPezbuE8CxGbos
UtGGIe1/ncgPAB9gybCvTb43KH21tYO7AKU1akF5JyG/GYrADPRSaLi5yd2v17Rk
nCeB2DLqaHCZ3ZaZmp5AIHYHv8ejM4/UoHc0pR7TdbJaicL5rPIfkEjO79QOgjiW
51SHYaM7mPsyuhYPp9Bdah005SoYNxXEgymc0IPj33+r3cGJFZv1Wm3Kj4fiAy7m
UZRtclaJQYA2Ut04a1fVEvxL2wUxcNUpf4mZSeAuEG0JyFs2Cb4ENDyYF728qemT
eZGXutUpoeh700fuAK+0CcuNwtkwKmTCaMpq6VKz8kan1Q5YmQTtxBGro1nU/CCQ
IJkhw5VbJ6MBejhJHtEtHfIkCSa20aLJ71bg7OseBQVx0JrZd86vOYv91fgMUgjp
U61vUHsbhUBTr63hMNJS6Vh95leh6XOGxaVzYbZYgZsS+h85+f53N2If5NTovYyE
3v2Me6Z0m6IDeswdPTiFFN+j4jQASTYcCfOGTb5rzPIpi1Pwd0uU8kZ5SoXFEoCL
1q2TkgST5Ipy9SApIleQpyXqT79mOZAmafvH7aLljNc/Z3MIvf8Ng3aLa1aXJGl9
yaCqerHo4X9XreYY/OETyXZtNR4L6XCEvx9t19ilHiQF7KZS6mNOwAAhaCu7SUsy
N9ltgwov6FVffxajzawtNexO3gkCTEjhvTxFeEG4IB/LtXEV52If/MYMZz25nbyt
QPdAfjBKJb4JJWZ1pvh9tNYZwP/BE00ra/ZHWh1BlBm2qOVuLc6lHGS2cIN5v9cb
qKiaAiFMoc4e0pSy1YqauyPka8CLFh1v54c0R63lxDv6jovqCTvLPsBqMj524vCm
OHVzw0oTEp9gdDyjsjtt80Unle3r7pAmemh2fbximwByyDrlE1VH8wM7kexR1LPL
07Ox6QhuRC9skWFDLeByswq5V8irGcXD8TkvF/2/ghXRtXwM1Zrcb6+HEAgbLBey
ltopzk/BZTCupBg8rd42aXwEpSeHEHvh8xDsPDR9oU1VPJgYgDQn/GG8YoDkQgwt
qmp7qcprK5IZhFNnSpJDcczI9oBYQRQhb3Z0QmSfAkqnBYxDxQqOy5XNyJQGYLuH
mhNdOi3KEyHspyhx+rJvgkuM0G1V4nQgVfZIw9euDvK0Qt3+MEQxV4oXfNYMnWgj
2Yzz1I4FVxQIjUKpxxFyR4kSm+kQmtZNr/IYX+wlq9Mi0nbOgnatCoEfLEoUKIMU
8U0kBvjbYqWJcpP8QVJBHDOkd2RNHzCKQTf8Ya+RWXwjFfbgjGdBIB/Bf5Ko9E7B
hMtjh9LYdi8AuCSn4RZFbxw6Hxq9+NrJymMEb9/KjlWWwcrISiFzZUeOcWYwOkKe
/uPdISKPMT4dwWfThuZdGKtyQKUqr78vrZTWu4zL8M2UYs0LfgGRsR8ncta7r/YI
lT2ft3/nvMGCw8JSANAP+YvsHBxWtUIC/rs/ZrJaCv55mJmOH82V9C90NrlzWG/2
dRTw63XFhUeCEdB9+nTc/WqTd0HX56DA23VuNggAurQk4xRMRzBXHbyEI0gRiqkM
AKjQVJfDz1shqFVA6KPbNeBD9B8IHgx06bmtucVmiBHTkll9rBfLZFx/C/tCyaac
Vs+NRqB8QGsu6smnTuiCh73Cmy8aY9usKo3iGVt3vTJJKNduQOfR/RXrUZnxzYnZ
kW8nlxbm9dhMPhcKvJmeEF3rrQvO8yL895l2bVYHguWUgw7vZAwwq5K+xo9pUt7A
UTJXgz8MoyNzo0ZwSjkJEK/B1+NmjrtvpOrMqla0KIF+pEIZbIZYzmDifXGeWIQn
y3IaRB7gY8V3nxF/Rgo8uPBsfqQ68laJvVr0epXo9HcmK72qF4F15LezpB/nLX9u
h5gstHiwEcwCxj+0H7wOAldCRVH7NXnYPf3osdwpaDryV2Jn3NYubP3RrbYs1Kbd
WFl0LpBeXtWSAnR0O5Kxb0K5W6ps0vPVAIWoNzqYZ4RPdjG1rzSUOKwCtAebh97J
yyxESxr4IfPaZ/A8WD5/jyH/sjJk+Z4A2sBZ7VF2sL86Cb1pDeTWV4glfbgawo3e
QreWVgz8SyhB3S4t2GYte9oVstDWsLN5XkhT6nKcYxlPWJWONE7YMH4EmDynoQ9Z
fkoMZTvH9AQBn/Oz8VM9OHzKm/y6rHlDnphbBmnNpnDPFawtGyfX+qVmMkwmKqD9
wT4CYDG0Cq/gen9TJa/Xvhm5Vqxzxx/OaZSjRWdALzAcRSkM9OLDcN29aGKX3rCW
i/85XQVv3vtq1ehugL1OoI/UojhHDoz2iRbuAHJDszVm5EpxCcfb3ZxYthwG5d4x
D6XRJ/brDZjNUVi9rZoa3iRu2SqCbHA/tK4Lg8r6oord3ELncgKssr6ogz6Eksu0
5e0qGg2NZjnKWBnB/LyLDcpUr6rDY7Oh/ZbkQWx5oXIQbb9YvRpvTd3tzR9iUkcP
+qUzDFEGmFPxy0UMqRwX4WxeDg9cuUexQrwhs/0Mfl925x113iliFhgGOaTeABUQ
DCHwTC0JFJ4a5kgBikxUMwP2oUK0MYzFBhEYOvoYCv12bCZZwI9n6hF/B8rwF39o
bffF4f6NWyyLIE7YmSAK/uIokN0aLz7JFl+mZG9pfCyqoTHavq109MAF8w40rAwA
DXMt5qYKufQZ2+kn1zxQmTBBa7lKzplqAHpV0p7eSNcwFYeWFLCJ1Q59S2cZcnEG
kCCdIEjcetq7v6KtcohkR+aGo7390kZ1pracoPEox+IYeqSn8hzQr8pG/yBj5mMn
slLS9Ao+2NOnU6MWLdTHItR+EbHjnAnIUabJqxYXCRohK1koY7qfLD1dhhcr746e
jfdW665Ldnm1JO3jhJ4d12eDmrDpEReGCncC0ElBDBplqKhChpiqThE5harJjmZp
IH2caq8EC0nLJcxcIELQ240///9gyOiSki9MQAfcv8z6qG5J/AfCmK8NHeF9BVdj
fHy/KwM7Ms/+bTqjOpirmCgYavikkHsVFBFyZ5snxz11K/jWGka0bjHPT6Nqz1O6
jOeFRZ8+K5co3fTSTwQKKYltAJdaUKZXKgWrn+DrO+21jWxKyLTY+9w6hB05mIBg
GAksLducJq2b4XxFK4z3Xw6IMbPLDu7hqCR9WsmOr5ElHS9mr1pdvZgmeL5+PTyr
aE7x78ZtP+7KZL6fukPpWEpU5Ae0tbdCh7h8WZuTpmLW+/x/o/M8sLV4a7zQ05vB
R8uyeJaqIs8DG00+HHoCSP15Sri9X4yMe4unz1JUifLSk3AnC57xDPiC+UfU6l5+
FOfo7rx+T3rZpwR059NRx3diNm9/50tbUvrfPNwGP7c3vrqlrYw0rUdMM9pRY9Yh
HCJvsRJUv9acJ0OILU/QhioXnUxZiiXrEfvcNvYnQxckx2mLXeEC8QGR+OL3emNS
12dM2O5Ewe7EzX/JnT0xlJu1QKxdUDR+lhOv+n77EYhBE1n04afr3XD+CSkoEAKr
7LNph0Q2Nb9tJVWLzaIp6LCV3bYLwCUAszsNZmUtbKu30P9EH1geEqEUq4N7ZcfT
hHIDB0WKi5rSM2cwAugwMwnEjM247gf+fang3ym2TY0pBh9zsmVBgVPpjFlxalJx
oEZ4dpt5OGeQipCiPdOxKMid8XX9GIHA87rFFjJm/LZo4vfmhDW8UymmRueshDua
K3MYn67vWJWEzX2T+nGv9r1fmXC524ajliGyGL4kWBvao/sILojCkUuTxa+lHqdG
OmfE9zRjDDQa/cTgXb02iJsW15FkCHKh4dy9FOPWGCeIZUA+WGMfmjNc9rDPZqYT
6gcB9VLbtetRYBg4M2KWNXDF4p5EV7P8stlAJ0jhqOPydWg6muKFvHSM0ZsJWmlg
XC1N9RAHjXTlw/4gjB5XreUpRcBO1v8wYrD0FiaXSVnsj2gFu/57glnIiid7IHOp
yzBjjFO0k6CEqSvnS2RGRH9l5XRRfLAnW36alXZVLxKWrxrmElKR5RlunoDn5m1M
VYy7IMV9xCCdnLXI+YPApHP6EhwRU2YjH98skDU0xIhrg+op/Ig9D9/sseZWZoFS
2XRqqqwvqnwK0NdzaIbVV/9gcV/va+m7NQkC2blnPSKd3APjvIGgJWH57ePeeVRB
JwHn9sV9ds/ZjuEv0xEATziaO9edYh+GN3gDtnnTrzerzLyI95ykpfbkwC8hRzMh
tFv67g9gFkAFf7CGy9HxtVYyMHr6sZutW0rZizZXK8xwbOhqlCIBZzQ49sT7ooAc
ID2ERIcRjYCvRDaWN6xoZ+nQMxHTLFw2rHQDf+xvXdmhl2YMPjbJZfo240jWz2OB
/AbfeGFBPKmrbKqmRZCA5uasG3rNfwihYQ1+ZJCVC5NqLkWWGxSPywK8fYgi8jwa
IvgOyGCR+WAeOWN+QwsiPFFoi5SBB3vpdQwqeE/yHZIm2mebBxMLy2CySb4A9SVF
5zBbHuC4kZf5JB3Hz6CaViIzc2F/ZZQV+oW9/7ypsxzSu6OGxG1YTc6oHP5pSfwC
oQ6Mmjn0rltNHTfCljHsrdfabswZ6QJ23BOjbkk21770m6uW5fdVkrf+c9c+Tag0
J6dXpZ3Bj5aHL9WrT6m7fD2x93sW58XZtFlQ4gJ3c0LixGGxB0oPmBP5wnfQinR5
FjM1nHgdBODWs/g2Z4f9XDxoMwComF815faU++RQbnDgHES2vEKVbq64YMlDf4Xi
7pVdGDfpBOIrvyAd16tX86Dd0GO2BuTG5SSIxOscJxjc3/d/nzbWpQcavCirSnLQ
n7lDN1QRZgut2Kaiy/2UnAxrzOmi6mhKF4hdZd/taf5NPq0svHdW6WOHMPUSdKMM
i12yhWfpjm9sduHgVajJ6xbz0x07LYVaEX+V8Gzu0tck/AYbuLd2cLl6O8yoCahj
0P5jCS7QY5VwIdHDu/vXlTZvNd/CoP/H4d4ZrhPUjR0cvn0KIxIV7wIL47A361AR
jVpJXH69z9slUreAmt2bTvNrJaImXqm5zi73Kn59xi0YbtvI+j5e1orrq8L1/eZv
n4e+EkA3P0JdgA7t1aWSScLo8oKJSrfg4rCZPcwCQc2HerEo90Z+CthZA4LHOBRT
8MAvZTOCZo76JeBSv6trBrLTtah5AWWRFLRQvBk5TZjDygeMnIQ+iEKdnAj8Hsvr
fn+G+Yr+NR14oEydFwLQw399baCkRP8whOErsvBWe9RoznrvnXzuZCEZUlK1NA58
zSmS0c/JGuCdREBhVBtZNn+QJ9WfRS6v7GnIw7XbjLX5aDU7SIcZ4ijEakLx1llD
SGsYumKCMkC1u0rSZodwVPvDa0QAiDmh4giPyJ/BReLVA2TA28bNtPkUQ75Muz4C
wekolSrCOqhT71Iz5nWT+84pW9gZ5QgKlKQaaQT5pOa7d31CKqUgv5k2EC7MiddL
qZEG7m+pPt+UXuPGCNLb20B6BQrO6U+r20kxCJK/WxGQ9npKOdnBw1whY9RQb5L0
snIjXRhAnPumWQM9cCiZwONwEgv6264enyyZ1EEJUTFTl4h7Mi9+w2H28Iub9jsn
E5GFITj02OQEoTViLdVohKmeBz1Yv1WY3cNMbGMwjRGiL4MaDOMiJSE3CHZhG+0H
0sObTgQSngtm6FWBdXLOuNwAgqS8f+tZCDaJ9Mnw7PvfWBj58t9MHFnegyrv+1E/
yzclQJtHFct7y24PMAV6VkpWB18aWPd8M7epOFq8jRABIBzggofuswzKjRdAyDlA
9iwIRpGyFB5ZZ7w7Sx+725SBh5k9P+27TbIZEnJz7IB0eSBZV9nglSF9LAUvRT2F
mJZ5Dkrsh3wOuSzXBbVcLv3HQqEfce6nwaaUr0gK/c1xlMf+xZRZUo0nUBfQ/sMw
jDXkqxU3PHVER10UkJtCYEzWKer/IMoryxQNhWfnV7I4gH8Ak/jvjYooWPq/uINb
vkU3ouPlnS7JW4tPr5yiTjTGEOUzq3kRJG18Z+5KvQEUhw36nqskUgza7uFSl/0Q
RTAZMVIU+WgoP0+G2Xm1/YNoloGK3gdZcGZ+9yllr8OsrxWQxTwLdUTgNuJe19Pv
ZDXK0uqQolD8lPB9WytQHvsUTRLAYBwE0PEY6hHLwgnDjOO7r18LqyG/IqTtHxgR
GeYFMOgsG9UY9rQGzjU8RmubTWMmkRoWwhHJaeB08h+i4NYFstX35iEpGVnLomUO
JO+A3XzCYsoL5e5jXXUgBGrCkxXDQ1EUCoulbhWT0wNSsipHfZNqcatZk5ga9pvD
S2aL//yFpki4AjrwF8AAjO0Gk97esojMcrQh9j3j7ytnmngONEfabfBJqQknYbIf
To7odBwjIMtLjwgMYQ70YQxT/2YHpe8MmDYBlpyz8XMGgUNKD8bfTFThpUvVkCw9
jnwsDd4mTKc+f3SyvIQoMMyNlIsWXG0GFNHgXGD1DoJ7Il27Qm9dBabJoX9VUG2J
A+6HJuTY7MZqFd8ilFhpJN3owamJPwuttoH7f1+kLcZVYJx+8jzH14ENZwSAo1VH
`protect end_protected