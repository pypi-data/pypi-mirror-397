`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
zZSxD+gXg/oJR5jdsH5AQ2TVPE8YLO1PWtO5IzxrqooIp8KKqLhZRAi6W+yjCNul
Q7RCgQOLxwMbEHUjFnZuKpoua+MCixUftTqKoKorAHF0PeBi9zCO2DLTL/eu7SZ/
UmsaXlgwFgB84Imbdd4/az3QP8XnUEFSHxUfwRVLEUYOTVAxaqWa/0jQaOoGtNIR
4yme8/Wy/eaEjd2bLDDIHrXS2RnV/6dmH9hMKWVpsEhuoHVwxg1w6dOyP/coVoAN
52EGQYaf4Q2JEekIufVVhCeXWMF3xT/e4AKYcPwRXbo55X/nM3CkL9YmW0JkB49m
0JI5/oZq0dee/ciRKO5eU5zYRK5RglKXxi4s9bzSnjg8gcSeVSk5ow7hftjf/O+o
ROjxhE1IjBdL3RNu6lORCWnUaV3aVcea/O+WrGmqoMyeUnZWkVFZzks47OQngYWG
TnpZUl8KFgEuNog7qmUyzPxV6lIUEfsdewCPI56Je76kKGXEY4FxYOOkGUbuHY8X
5YQMeOYQalrYwfQqewNcnTU1si9eyKDNDI4Q04+zs1rql4OAP/dHYajxUI6U2ohh
wsMiU3G+BXzAMSFAUmcP+2jrZoEk4AjXD/s4SEIpREnoq/40bFRnOmNkfj2URTBE
AU4MQQIafOgswmWt9zCdh/IdluzfNNDO6nnx1oD2MttsnsP4Bjk85w+dAWYouIOX
DB5veFOmZz6KSbZvHbNhBg/ZBtzgE8JyyvO8Zt7WCHVczTJCvrrkiV0mapE1SG4/
Uk4Nr6k7AYKq4ZkOk5EoXfzZUS2TBlHz7XmOJseVt1YsX9qiLTrfPmWY7P1Ix/QX
vRl0oXBF2beqUs61AoG6q/de+WmnCOuRng7tztzL1/6qpGIcYU4r9CxxEQBy/Z75
nFg+Q4d3QKWE7WdFZW/B9MVAczABwPVr6M8zLu7tCDIXxqIrFvemKiaHB5vD+r64
tldvVKphp7EYb9zVJMg5HimP3i+j9TaygkxUQmFcR1GWbX+zzwMD4c7Ic9CS07Tc
h/TXPsuaxYYEEEtAN8sxOlrFgJQYESe2COCKZLX0tz7cNhr/neAtgVMvfItClX45
aYp+Ytr3nU4i5hebaq+xRdQVczH8G6brJdtwc+kOC/7dHL/2Wdpa0Fxt/fKEE/ly
7b+CVi9CQ6eZtizW/IyFfa6/bARGrQvXn+fYFU6NUMWnSkcA1YHDgtTPk5Ia1ZrE
Ty7DHDBX6mpZVto7oWYIvb4XZUpwnkmlVpZMVbNEfF38zsxgB5yi6cY5tfg7Es1F
utcpQ5/CC+6T1ESgmzZ7eDOR7G2KVb/vILd4/1ptdmgmjAvevPR6N1+NAJoaGP5l
pXcJYoZCnM0lnnQNmlM+HWXH/BbO1shePp7p76u5urIOObe2aWJ33jdUITy98FNu
MUWPOB6QsusYu5BTcLRDv8eHO9ZyVMoxuS36qwLCzY9AYVoXoMhXJWY6cttfo8x1
nticwDNqqA5ES6yqE18OZpobEFOHe3VmVLQUbpSj9Vdo17QSrLHB0qJT+8X41woG
lYnRGogNeIl/AqZvIMvwKrufAjXRyDUPh225sjZlMq7cesTxCD9X4jfwdO1IBuDJ
FkrkmuKfyM5S+3XMxprGOPOg6JEGzmGn8KA2PUcA7eIZCGBMFYhY3mCOW/5UfIaB
7aFm32GbLaKffstSZ54IQddpW0Up4qfHSXituRD7IUUygbJeV+yE5qZmyWR3NC3d
ZhTDv5K4lLQeGRrn0/3Z6qy65AC/lA2FdW46GZeWEvdtXOkZDeYe6h9CJk0UgZD3
6YCVpdjvkrN0kxTUGzqo6fTLctfWQj7sB02V3PcEK9Fygl8LKOQauuW8quwnP5Jb
+AEeukRZH/H+9+O+5s11GnO77NfDZ5YShzlVpgFTB/4Mg87ud6eRPst0IlXeEs8D
hpvljCmxX8Cm12LwctOh0b8POeetQUbJ/AghfIUgEd21dQlVGMJzlTujWUZ8z3bU
d8JYbY6vMKwHZMMUwd6Befw4JYeXUtqyxdZLMg1PJmYORz26gtGNiMncUwhqaVPG
yLm81zesILrmU6RX2DCocTYWAG33D1FWiM9zvDrSmSHu61r2DNqItcbgI6/hHOZW
WXNAuByzc7oUIab+5xJ5T5D755Ln+et38TcwrZqyiCNgrZR05yi3y1nZFGa2W9o7
uBrkDg+ZjCvRRvKMSfqIr3WeZc4Hp5k1fo/6dtQHKPxdePAOAeP7MpR5u+RtOu3j
r2LEDwhxOOSQSfQ414CQo6ZovSExKxehS9A3ktbnBtBaMcEuL3zbMZvbbZABV03/
fsZAF0iiPUjstp/bHcDM+QAmOOv/9UylOc9WK7yhzCqwEA0MvAmxNwD0s7KvVWKD
zHWenpq2c9pkW5gQrM1BmjofZIf7R0E1TZq9Kk+8XebWw16RYJ1Ly5K3iCIOwz9w
0jZe/Htld6DOnTrleuKEFTgAmmTlaA//xxB9sqyujh8Y1kWU+BcWnm+WbOjF7bYD
Bbu9iXD7nY89+hTVynUSyPaSOnT2FZ39HXm5y8G+T9NdCiWKxaw3C0ouezzMMAja
OQXJihxi2dkkFQEQpBFd60IZaZ05iEK5baoSkr8ZH6AyzsUb0vkg34I/aOsGy4Ds
vZKVG4L5XS9MMYtIlZ/Ea+LF3CplBaJiqeyuIg3q6hj87UOpN9X9G9B75LnQb7Ii
LWIk8s+GLfBTcbewLJI54SHOuYzZfcIJDw5mnHAgDwsbVaWKd0CHZtaFU7AkAZmM
AjlT658eSNtEEt0EZgqaBQ7ajlhAmwQMdc343ScwGllegK4XtF2SlEzmlu6BHC7B
NDJoHhcoirZi/3yrUh2XEseK2ErK2f0bebytqhDU6L/9YVuSH1+D0zOXUNQr9eg+
7ZVAvb6rLPfEM11c82HlPQUh9pOpO6cBVfU7z7MMITYXX4nYDP0E98hJ9splLVUg
Ya8ROyiEjbwglXpuRPnC8wqYqGhI9CtYpaJmYYb5cGe/b+6yR+e+h/BbVmdSN2Ru
qfKCkNaTC9xHuCnRPiRHMdZaqjgRZ7J/SxQj17gI/ssc9ukeBiyMo5LgJFp4q2pf
tbvFsSC+0VFG/4H24+8/vHnRL+vzJbB1mdpRu8rncHb5Vfh1BFoM4NRTYzc0Ik2B
6+BXTtGrJQRVVhvXqc72DOPY93Fj6t+FervLFzGCf1njp/aE8HtJHSvQAktB7CAU
acQSK3NmIbnbCAmPTnQP+f6e4a4om0rIsuWPKGUh8pQHd9HHeagPvBzlbCS69MCZ
6R4aVZLTIlIL52Y0Gu41i2RQ//nuqJjt/Xgy715HLCdQvyV8b4AFaraHFCZDV0li
cojvvCwwBFuQqjX40p5OOtONZVvihIcuAFz5ZiuE0j8vDaYgpX2Sp8BBaz468BBR
qdh2Z4KH6vGo90412mkVT6eL1NtBISr8pG6OqRX00zUbc3rtlLGu4hNg+lb3P8Cw
P1BiIqOXUWIgLFw+ogaUPLXi4/aKmFKw5lQGo4hMJDJHwpJKjTeYJrAh+ZGVvfKN
hqP28oi5xixD4a5YnSFGTKNRdrjGJkzNPAc5VkEtmiYt0gtchQQc4Q2tEhzfNsZw
EeslK2BBg4A4E6NWXOfhdJHrqx4H3BC4zcRz83NPGPWldApfY4pLPRF9nQUhFzus
1hWKlVt4uFLJGkRCa/gTFhBg+gOMJuSdJe3gB7aKDt7Wntim6o7xehjLzm6PcRGK
1/MJ89Q9RMfUTOm4wju+/Sv+3kKzfUV2+hYDVSxvShp1Tfnbj9u9pwLkzp1d7e2X
S/tnCXMgY5k40WIOFJMKpRjMhQqUU6Jn28VOXeVNpM4wu54H9k7nTpBtC5iN/vvL
AnzsTO3r0DWQukZ/5oj4J80tSPH6HROLsj61vWWOCi6WdoM11oJPrDyN/0wrGvZt
f0vwg55k/mUbw8ed/MTANsGzL6BC/kRe9Gs8anVnhfmsOew5oIx1nb8WH+bIx7Np
z/S7hZcBAPbI0yjM9hv0vDVfoVKwtk0yjcdm62UXGYL0SGhAJvWWCdztTK8ICEe1
nKIhjwrp+OsE5lKGfnFv/YhdkqMN4VdOLT2PuLOT/Gpgn3C+GmXrlqMeMusFCPoD
eDy7IFxEjZxQ5aV9gs/LrtkVZMdy3mxDZ8DLrs0qtxksHB2fZI6IPqlFaxnJ722h
iT4OyShNMadj5dMDG/bi+gqcFLl4fjcEKYdSIUoqfOwCnRMSelKIScc2ffkvltun
Hx/+L8XFIgcvh5vOBV1wUpwgS3SXYulBgeCtgteSZofHDI9arnnBwfGq33VjJipc
GFxJNhWPp3z4FPvyofE4wPmlFDH/sT8Q8YpsYHadeP8okThe97o2UlE8Mu0LvSbT
v5FKgMYEOLuo7rmZRWrY9rsJ+rPlmxpaWCixJZd8zlrBMy8nfpqV7GC5y7ahMsyL
qzkeEqps/+p61Rf1qCRVf9/yVE4p3D5xp1OptquFZGYfVV9T1FeX2+1Pk+CGheEW
YBxmrMf5mhqqvwycT7M/HQYTzvNZP6Y4AdHs2VeC33cyzVQ7rtIE5bsBqE7kMh11
Ku87yRdjuuXYfmwLhqbWJFKcqxGzOYDfXNh+H0sjK0fVJBN0ULYK8KYvQzn4FhNe
NekOANJ7Tggn2wskASX7UJsed0ScTh02+o0qmeHgvW47QUrCiRIvUr6y89HWJ4D5
ptX0wJHQrPPRu/bt2BMuGKW5XGEVRNJaRHgv7KJmnGXAQN96HCpUIbf/wu+83PfZ
Gj99O8/WsXSWu16mspQ+REQwERV6TrY/Xi0fE1nELiStCmE61FFZUdnYLTii0ZCA
1RmhL7uqAXStlMksjR7gVAKMfROUmyLbRDsSLT1856xKxACqp6iEXN1+FrwVt9X9
A96D38Wb5TFCU9fCfUHll5bCO84oGl6NjGNc3fhrM1GXn4YB7jNDGGoPVqONpHOu
LH9sSjNITRiIWrKHf4HIPuJW/OCIJ+BHzMXCrlnL3A7vym2Hn3loOQkSF/6iOi9+
bSoGf51aT/23IKw5PYtRxufykfxpMN/n/UYFgNrvEdntePkZbQvpKYsKD8+P+vD2
RkWjwfWFOWSkvlxsmfcICMEIwMPbp9hXkA2Rj1w/lF6WNhrW7xx2Y2Hu5ynszzQC
gYV4yFEn/Zs3nwfadWMIwn/GmZzE7hAhS+aQnlXhVX5J8JoOM9d8kZ47RyX1RZcT
6jr18FBTn872LmI0/EMUp/Agev0zB6rykayavoUncFsEJD1X4V5nqrkOxeElHtiI
iLebndQOGLWqMacm1W2i92lbnRzu31pan5jmupr/WJDF7vbwOOmDA/tnrRTCmv8s
lEKJ3V2biWANOqVpKflDK7ibbxqjhjL5lvvkTJ9WqyN8Ng3yFw4n4lG6WC1HRQEH
qD+0USCc2a69ow/iCXDoMDsYeN3LInWZ9rSLaB/udyJ2z64KH0TeSqqwBEsA/KNb
hbp/0y1hbvcHq4Mb7cF8h8A8sczC+H6nPpBJ6M4mpUpfyWr0FczORM0EFWJ6Q0B7
WOFO0MtDjwR4FxXUs7yLbBWJhowVMo4kTexjSOyVSmGLqVMnPfTBf120wmcdmKDu
cIKM8Ry162tGGriw4GrhUialgs0KfYyNCOhJ3hKhfXMdyVXsYQJ+6EwVKu7s+z46
RvuQ4AB/ZuflZbVD2OgIm4JmKXCqjee3nCwZKcH5UL/3R2O1ELc1ilHdQnDaOTnt
TN1Npxkfz26VoejkLtc8V2HM1ufvQJ6KFysqO6OOyd/q5VCNGWd3V7KepbPmNQb9
fWukho1T5JpmDQH1eVoGEeXcHqtoJb9tFYlg/nzE7OIZJFUIlYOk88XOwYVRIUMK
honkMe+ED6fuDJvy0vCYD/DRzsNvxesepKUzZHnS1TNimMIFe0vanKC5FPGmClAH
NtPs6eGF/Vksfnk05PWSolx1xkSDJlwU4F4/ZsymLRIsslud7PcLiU3VgokdpASu
ze0wFKoT8tAh+IW+MHtr4XfQyi6xXlj+MLerUi6O8L73bHOm+4EiTh//LQlEv4PX
xIxnfaORo61/JNLZkv7Z3Z1vCFn5RQuCNBWdxMOjFCigroPD9CW1zNGCF0altm3O
d/hYavEEEnaJGA5XRK/8ArcKldbi5fONqvceHgWPT4EoBOxp7IMPGv/C4YzXBohM
ql1t5sPOgJ0fnbBqSvWdaOIcW+JZ8KmGnA1MhIUx6viJcJlbzgA5KuWhygZ1Y0gA
GLfHbLIvg1svdLODW7KZIZCxe81lgvna8vLOBwK1kY/Q8xtUh/3i02tX7vos3rH+
drla7MKNvKc+065viRuoNLtomZ3eE04xVZEbSeNuoRijLm6W/4zcO2YKlbrqmwHl
bpqLLnUBLW6E4ELCiF/JwJ4969nklxeAIR1hRWQwo38DVIbxjWFEdvbCefy2d/cV
K9gW54yaiFMB9vOeNL9J9Oc4zva3aeWzv+hNieZ2ziA5sm0GVaEJaSJ0J8BUlM4j
5UcSt7Ef0xU89IW4ISlliAYDsIJyz+U7FiXf1XCKXlttTy91R4Dbuog6IgumOQS8
bq/we3HsZQpHxG22S1xXUttmbvY3ROChwmtfCRDn5w6qPcNd7Q6jBanjTENWyyZB
LGjL7zJram70bdA+QmWCeIt9oqot1ZriywfsZqsoZBp8PAXMMESmHzzUI7ndxVWS
5bPoaHDwKRLLIrrEoMkxNuiHqnVLPAtyMRO7i1Sz1RrqZOjtlg9trbcw58RaKVxQ
9aZBXFpZzzses/nN+o2v8h1bptjH5gkKXKiwDc0kzv0kB0rF5od2JwudZIENKnVq
66EaRa+pmQaSzvznkBpxwoEH3pXMEDD62JJDeH8EmiaNBZ2xQVEEeOKVRDM9qa0u
zyvDqZ6lCfgkpey3Eh+ZoRUM/g6Sf0+UhNiqZR1VRGGJmfQhFkK01+F8+C75IKYO
rF/tVtlMEEoDACKEchJ65PKaZFCEIGXDVBSWj1QZ3eKj3YOYbDpF3RDLrlGtXuDM
3AxYZS9w/ZRlLyuD9Cia7aw2cSrJ5krdKN+TVWDOEh8w+8lEOlwjKdNmKHs2VSJR
DKt7a6+XlA3MnBKY4C2XsvLgQz9EdxhOcofyo1ohJp2YYEO7HEOJGB6DqfyNRFQQ
iVv3P3du36v9tsnGlTlyBkZVEM7p+IfOJRZVWyWaSwaahPJ6XAqGrud2OvG1fLFl
lRXdU+Kege9z3bOm83T1zRVEMhXQvKH53rqZ/kdgbmni51S0CBgAU8L1LsKC6Mdw
BO8SRmf/ZthszRafpR9sGFuXTbIy4pCe3zyRM/a9z58uch6ZmeyOjELpksCosmNL
7VJSOsM6qBQ6kIlhchk5aJbsuCJ1wzlSb6DD790e9vk4KQQChO6NUOVLg7NSvnzO
FHSADt1xR7F/tZkn2GDdQw3P91nDlG9cWxPg4wygdKICktTwbZ2Y32abLYxezl0b
oLpa7Bu+7KmtxJh2N+bTYVYzSA/qjLIJyHiy6/0JPTexgHzR0hwenxMEDQ3FO18v
yvbv5Uy9BTxlwV4FKJw/wIHDdCX+/k+1bhQ/Qz1I3Zk12Ii8EtXqOlIeVbNb+Gn7
ONiNm7Yf/F5yah+7W1ZniMYPH+CRcqFR7GbdFj31EfCnZj/TTMGzgwJF1wXaZva5
OJIaSDzSy0cJHUuLCkc9qjRrTpI2x0UyRTKXXkYQgg32vqmhrkEpDJxu8ONPxr/Z
4egH/6WjY0I6p6PmLbLxIPC3siTWfzx+P43cBuZ157v2dG+bCl4ZNU6/OQVFy3NX
DSKV2CUe0jx3bI7aXvGmU5Vxo8ylJ/1oDlZuodVxWDsXgr46czI2QmKTnjmAM1YP
yN5dozdBQQvQDp59CUo7qIJE5erN9817dB4lV5YoZiI5UFDUvur3SvdOZk+lZRND
OmAa49Ot9VyWjzmMtHfGw5AP5j6DMKZzjsmjd3C2VeYx3EEz1SsFGbANeCep2UHy
q0X4cMQLeyqxG1dY0pnCqz9b+AR2aoAI+aiSOqB5AqAkoaOG9fZZ9cqQZoHA6Hnc
2UOGlE3nCWIqahluoRzy1pkQ/R/pBHwiTnXH6Se6MqOO12fdzbi1/jo3fe9spmuH
vtlN4n4G9UB0J8JuqA7ZvlYwMmU1uuUaStF4eFL8Z3yTspXNN/gXJUaAGja13uf9
X67jxkb17EwB3nWLBOSJHRpVI6jCtzll7bdFwm1WxExTZPFX0jnWNInjlg2XxbQx
4rRs0iwUJi4uq33wDdOAo2Gmba7YvdEK38anbYu1BzOc8JbeTIvyOdWSK3GYdAC1
SI4pgoNyXNnC2gzK95ZCnCcZVlQ9kElqhXihSuN0hMAMQBCG7vaVBbdqRfop3PBv
ismYstgFfydJMEFiQS1uNkupbU8SlmtkksvAX3+iygAf3rYKPVO01BEd+MDSKy07
9dGty6upQTBo+g4iFl8jUL3ln0UzmzfbdRoj9w09mFJRA1OcpaXSeSdUs2A6LpGt
Q/AG80PeN5NCU5rbK/iRNBBb4kGDd1+btcN6aJoYQLrxVcYY7nvwXGn+xCo0PxyQ
+X9PoXofRscMOKedRDGIm7jDx6U2BI1SCBC887XHL+NTgmI2YuOkv17pxkn/oDS8
MRKMqbWOY8DSOatCvlFo8L69eLuk4Gqh66DQgSbzO4ZrOb8RV/psyG8p7xs2GvdH
vj7aA5lxg4d+LwPaWmrYMdmzFpI87OpfghLaQduKZZhAjk+aUJk4713WMC14I46h
uVwmGKEOLURHLNhr/99qCYEjsiX5aLRSta2emAb9kka/JwmWF1aoiLj7JiCSOmae
TnAeoXiW1HZmkUv2D1wPcKE/6PezJlHrgUpwKpxrOkCVHS/aum7WY6HEYpBGOlat
dNvneELOzFXEqa4sCk9iRQMZVutq7xrpsAWoQfjycdJIA/d9ydtTa093ToCoBdl0
EXI7aw87IUKMftZ4unNdbAkZBLPSwKylnyGBri5XgKI7umfnWvEpz/MZENDxjKOX
uQ7f6oFQUbMheKNkKGZEIUzlX9uCZbOLsGnhtDR6Xagysg2a0gWTtJi3Nz5w2MmI
ET0Gm5U8Ad064hpjtyB/TUeNWiz/ya2Sju0uJ6zKWQ+LRTx6SY/fVTOLCKrBms+c
Mmdo/v2j/vSUqiK99rWOu6XMwQ1mgPd/47XqUVeI4tst3PFmk0XLF90RoVrz9/Ff
rI47bLjTeYWeOOfiz8UFCb5WfiMXCpoGuGqWjfIa9sKVtWvyrlpBTpPYQ6CpzYHd
ghYXHNjMF/itd9myk+TaFok2tAmIWO8Fp5wKX1ckF3c7/WKHHez+7qkRjS1SGwXD
osziwZM6hg2m/iWSkVh/Tj6Ex8MtS7WjcAXT47xwLbdj1DKy3F12eenX2kz7jgD6
gS4lRUaGWEPS29GCpy3qBG59LMzHA3M8AIr7YrequPm6LEnyWD2wtK6odSJPfp12
nVHQjW7njUfKp0H/Ezky5u0zsecLp6mtcsloVxSmto/srcapTW3eYLbvC+Rgs7Y6
aAZ7tK6T5Ld3eDQOSpri5hBKHQ0wmFxPIq2K1OxCLSfvYAsY9piP4lnqUx9Tmvn2
vGR8mfl7759WsqY+eosYxdZodGCk9eQoEqtjojBgi8IEvRQ1GBz356IIzivbyPzE
YDsZelEuau72voWjL+gwq5N+jTOsprH7PxPfuzaPcPFh9DhRS4f7R5mEBM9gIv9b
Ed8TvW1N8N0DbRq73G5A5pukWagabexexgDm3A63t8P5ekn//GBpErShkDauVpKM
0rgMZc9+V81YqQZo0LBCEDwn+/32czaidA4R3mk79tm2OGzj/OZiZdyxyeHPhz75
/S4v3EBCsfw+rOfpmf2peYah2GioCXeca/XyRhPwDu3vfDcpBZ8N43dvlKgTu7L1
7clo56UBpGK/TC74j7RrYPJMXeXxZ24C2JqxgQAYKs7MN9+SNL3jkSDkGvcqCK3Q
3q0fUAiYKgiLQOxMiORcFW7o3DT8RM77+O2qud0N7V7r3A7wBynIJhQikmAew7vz
DNSK15vsJbIFmU2Tl+YdLw9WOAcFm2hKEDCLWi3DsgMscmPBMK2cVCeDqTazyI4X
C0vHOdXbe1ymgocy28cwpOZjHLQkQRB3tpglI/8wEIHCpjaovBB5c3+VJjkYSzAK
tjdw8Z1ZLV9Uz4bOdtBT+dxNJ44HI4cgGcyMfBZAv9jhyHox4qSUaOdbD/iDIuG/
Rp/U0VHIswbTk3dtmR/HioXSE/6H8bFxDvD8bo0ouWbgxFqgiSQgHdO3iXDY8s5i
NXCF6Cy+FBS4PoCIpNOAwwk2Zn/EK+v3oQl0GF3PTjOq6cJayGmkMWjJAe/VP3b4
/m6MIPiY1fhg8MN/XF+HtB9DjO8qFSsQned+pjdvpRTzF/edC/lujEYj8IkONB5W
Q6t72oeVpT+xJojnA/SGTyyAiB2/D1agoRsMomCzNKqjPJfuEbB6a38PJWZCKBMl
lF6lXWIwhfm33Ne5VTULUyLbm0BbfNHYLevPTyLz2tD4QiOJ9yeozF9+cozW7Em8
9QuUPjqhSPP75WBmqVtVZ84hs5XAShY8gfUahyTGeCTBT0Du3lYUax2wU2ZUBYGX
AkDxNJpxMVn50c+Dn39RFF2xJwY0B1VZ/nBVJXCEPnB+WjKJ0GzCLAXn8lYJ/TSk
145Zc0WXLbdd72XhffvBkocdoifVBNP4+GW4Em30fNulBTd5UAnDrY+YneRp346Q
vS+PdudTCfQCGZEJeH7xx1ebHBzrGXYHtL6560TNpqAIicJo5C4dJ8gGrhgU6i3P
OaW9I4wdowZth64nmPwYtCJyUyV8RQjxwz4HA5tvGZkcccyRLhvqZkHJSFodsQ9p
VCQeSfEa1vJFpqT04mVyGwOrH1AuF17hGi3Kc5RQ71rCxZ94BSF4BVwX1JY5q/Uv
Iwvh1uKK8sYMB2ppmX+83pWwOM4De4bvXCK0qgmMQcKQzR5F/+0DntJ8IZ3nn4bO
Q6YXY7lNmNGqtkv5hf5MN3P/V38XLta6sBuae6oPvE2+MOnokNO5Jxw2u1pP/3K6
YUu7liVLcf/mtykda5URnsBqI0QJoByTqWrxdglr0MIhhkGMue37KCLCvc0f7Eav
75pX6FF02/I3e2XbyVUVNxwU5A4n4qekKWxF2aMYeHoUfzhk8DJBEV/MxGsKBli0
zXUC0u6xjBKIruT4+y8GuuLN2RF99vl8ZxD2jtOm6wPJu6lbKCDOYkxPH9uJugUf
J3Kt564jVJiPWAg7cYnXqFFRVYhJOC+dUkAqzbKxv6xMiL34HpCRVwD2BJHZ0b+p
XrBCSmcXsNgOnNblQJtPTK5uJz2QNVBUYJugDnOYhtoTSdy39hrCCYFFfiKEqN9E
zFLOkuz7RbxhFm+GNB5Jn1rZ/Ae4H4WhDhObGES7W0G0uSMl2409+tGoi3dsHSJe
UVNBv6PjgYUt2WndKUfcXRZBu+6Y/wBoh+WW8pZsfOUkKB37AtNw7fqjF+cY3z2u
+X5JZKRiZ4Y7DB1kTZ+NVe7SzTv1p1AbA3Sci3mlWiViSYv7P4B5k1SW+TcCjAjI
fsROLzZqVCYD7+aQ8seX8CuCBkKkKbqVh2pPAvrkrnq+yGXFhEJzowm31g2wPkdE
qPl9T+oFQPvjPBntO07KsTJBPOmqcbg/A25iq6ChRNbr7npcL+WO7+cVwDT5J95z
WhMQiULkw8nz48UtQhwF7B3NDOp8QoibwdXCnegECgEUG2rJNfmF0jzJdxuAXx6s
GcuuMvzCaCFvpEnI5oDHtZ+VS0GNoGyHCY5Ianxu99quHA+U1SkxrIA5bNMyq8dG
ra4VFOQWWGpdgx9b+OsVMcfV4D4IHK4p+I7RvHsrG4CgGuksckm04L26iH4DZJMa
H3RmLkbLckxIWdfSJdErXuO9q1jZkGHW4/3aAyy3R+W9DRoOJ1qVbcyQseYCLd7O
d2jBK0HZHM9DHTsZoDDkUNNbLfkA8eo7b+GHNzWbSZC9k4SZ/Q/EoS0SG+v7Dr7X
LxQRZFjn9yW+tbCx1IFcB3gItEfPwb+hcZTaR+edM4573qpzY96pnxNf6Rf/dcc/
SB5GzJKgHQoOQ9wMQAxt7Kz1xNokCVyLXAlg4/V/UaPwubADjXoz+Sp1KRd773dB
Dgc2fmMDp5VtA6exmfs9nfkxx9qAXP6/ix3jXFNEYdmFTaiH+clpGjF5HC11PLVq
19CerFYnM0QC01x4aWGvng+n4DXPp2/JfdOPxObLPlTXjmwGVgq3cb7kIwmewQoz
JIsg43lLHXJ6PPwBicxtJumj/Y9TVoOHEUmUeGwAlNkXZmvCWJNyasPFlAByHyB9
kCQyEfJv3BDcijamV0nJIUrhXyKFyBzLcl1D26VRtFdj1pMYueowmz83O5Fx2MI0
UbyO8kTVO44pAJigVZfTmlfF4KQZXvzyZJYgVIS4GoNNMaJkGVcynz9MKGdsrxlW
it/J9qX2z11qgyz1ZjM7zMZD+FvjfyUDqP8CpoL2C8B9+KCH54uFimDeWiMaYUMl
GzwgYqvtq+V8zpQmVcd1v9jIhExbi4RsRDov3AJDaNqkB+EnF7OpZfBIsiKNWAKq
dnjBuEwzIL3KpJY8GnCV6sv81pEDlMwbAmbFHfIPbCr/c+NFUnnbDkVSBGEHLxjg
TW0Y8cTqazodQnnyyFnAsoJNWuc6WPq/laQWojK1SoMvWJ8jQzK8ZThYJiIpNgtP
hq2upaa9wvuL9KMKgclbz9iWHxoNtmQzEtLsBTs7VqqE+l+thZK4n07Q1R5ZlKeA
Pejoo7YQnKjJGnnCZmR7FGqu65azbjp5ZClpVx2KJCUHjoFt8Ep7Jdtmc9dm9hvc
fYCjsPEJ7mAYCSk2Wq1Sn+t9U+JAoDkzzHM2w+xsa9hsvY5FlOu5jRmEsEfgXmkA
1Nwznp0rwuUI2k6PXLyWM0c+aGPRfuPbkrpp4YIKNBd/aodKGZUVAwwzS2ToJvMe
POeplF0np/nA1e+Qvh3DtbET7kvjkbuUX4D49vXLyF/ups6s0NoibV0k6nKhXIZb
l3f8LKrtJ/K8kDvUa3MtKxnLPHuylESbe7TnGtoHeOaDCYBWm6e2F7zHkTWQ14CR
1P2XytCEdxDKRjwKT0keAtx/2vho3iLEeLTxVfr4n1ore8ulZpPlAG0Hn8ODpMNv
aZMEE2R6EzuJSC+H6JEu0diXh2edkVRys7qFCegsBNYmFUwN6ZQNZoTxgK5G+5AF
T8jwZLo71wSoZ721I00ohh6Vj1Usd+OIbpPWDSzEB071IU/069Ip+brpJFbSbwQI
j+ajrCQemsDqI9fS9xDt4cd8vHemLzwtrYRn3/qDArGN2Xc3Zg61Kp46zb3Ve6KV
Uav8iDR53vcuXzreAl58s8brT3jqnFgCmX+m9oeC5yFmdrsM1IEmTv6l6gn5ZmJ4
HbsHVBSSLcrmGU4M2WjiL8H1kYOjYzWCzIuRF/BkKOOf8wcsHoIwiAcCjpker92p
I5M4gA2iDi4u2w1979vDsIS40B5Fbq419RRaBANo+Hht43UEEp8CdJScPSOQTkhB
/Xt7pk5EZ4vBxz7j7nEppbg7n5baGqOqApaML7LyfIdViNZ2ofvXfSuoF+r4XEnx
TCQ7QyzNpNGRGzHh5uZ8P4fQBD9DgVdZT1GOqNDxpOmFe7T6ol0ATyC3yMNyjVjJ
921RnWZ6Gq1ir1uP3pGJAtWJD87pGnKyEcUet+uCb1c0MHmN9ASpZIZq9abG/3LD
lpYeXZOKwJQkhFQtVdl4mG5Z3Hrc+H7BKBsvceqfz609AM6zEVf8TpqUh0Ihij5Q
FYy65UUwZ1Zw8ShyE65opBBEE9qlI6pbbRX0HGuQvCyCh7fqlXFfKsw8+UBP0ZMq
yN/lE4iLSzHt2BV4P0HXjb1VOyu5hR1OYolQSVgSmasB4BfaOUIou1FBEpPRYm87
bDgFi6ANiCNgOFVJqyhJtnDfzQCUIHos4IwbnYfxvb58MuBfIobj3cJxIAyiQuV+
aX+Bd+WYanioudbdaWXZCQRrUQhIaEDLyyTd+ediMc2ALX+OR9Mh3mlIM9IB0H9E
/N4cLBOVEPq1RsE4aHf0QRWdeYgeTDtoZNbtFU1R4EYraKXw57Yfa02BfP7+fvAG
QTmSqzRfCFMbG+KHgME3IIn16DM7yOMu0wHcK4pGF77wqb965p/ilSZ5vZD6lfpM
aTVVYOQIh6nZEltW1/GIYOnYqyl+rA6O7a8v1bhNQH5qymlcE+DE9ozJSUYVQ7RD
3yTaYvJsp6NkaicBrC/kecKwnPfYhWhZEKBl5uk0HaY+oyswpI9ioZo4v3T8+2OV
b/mgTMDlfxjAoxGhUm9Slq+3rGe75G5UcvGmtrjqP3MFgvh99DqtsNdYidzDltEO
+ax6sNPxmyfniUprPn8WCtxKVDNRd+zi/aEE1I5WJWqrPETzEMoqc7KS81H9yX2C
UsWh8ONx4nDuNr/2bGre/Crw3w5TklWCKEaiFxQM1YPuGYkeQNq/9wuYOsFxH7Ko
MbCi1VPOeVSQ4AsCSoWzSlHdKtEzPRjuC4nm1M1osGR/UNgdCj442SIo2YxgMAxI
feOw6PBneexQ8EcBQmpaiehSlPAtpdnC8Xaje4czvg/piGBF0TDFYUu5MmX8+7b+
a5X0AC0v9T6JfiOEraMoYt1L7+oOgQNhQgK/1zGFya6J4U5W1eiw6d4Q7rfbnWEj
rjnaKX4Muc3jqiQ+o24CAdebRqsX6IOqto87CxDu3wXZC3hBTfeS0n7zdjITH508
CRv8Qgq5dPAwxQEV+FpY2FKlO8VqD68Ofbr+dPfvEPloHKnz1vlm9XLLNq7mo951
1imyQpG9pkUANErrBgwX85h+Bw1+cCjCCUoEHETFYn66DIBZi2yBL3834re/4mWf
6nE9Kb2IIfGwFHsNm4AEAjDK3yrKfdzWIOv5NM6JBcVLCKpLHKwZ/5E+88ii0Udl
WDU5CoEAcbRmsS3AUU298EDetHsPtvhKI7Z5CXyAfnuukyJkLlNGWOZQY3uRzCzx
yF/27U6KZRV/dEarb4wCYLy9xYn6CHgujjXvhxR/XSXfssE+RDpdG+aKanPe/emn
ewuS2RlTcsR/MSV7cIci8b7gRgSp6KOwkSp324CngkmEch/2/IpEFKtQF4Ol0phh
bUjqKU+S3pmd/t/LT8w+HwfRqBd3t8nWGhlwHPs9I6j7J/4owMpxRcq1IzORdLY/
ybQ69YRHUBYVRUixY5kSJD/kj0YmbDM+HDbcynRHqG/4tob6OY3ELEAPbyeA+flD
/bcCVbqRtHCAtsaWl9Qk18SSPuTusR6rC9zifDLTWt1K3Uvzq6Q322JnV07mexAz
oiGlX5qfoQRRPazvqkwDMATi9zDwpNEixmvM0RBg68xYvRdYc6IBtYd0DlGyskWg
VODew7LYQcC4GNd6/H83t3TbQLvQTpjYyqfq+/jOC/npCDZWWmOdlJ8wgMkLaKl/
84KIC7lgXHmUWeCu8ue4w4imJ4r+WD29OSgcUyX4UX4+IrgyQTEaZ3Ue+6EtE/Hs
G28pPheARKuSMF6ON6fiknRBnvn9CSgzB04QBF1FPKF8R0FcKTEQxZKXJOgOH/2n
2EPo7IEHXHuvfB2mHKikVny7DHx4kfm5FcJoSJB8dR/fzeqpyh4psJ9TH8sA9uy/
OwLLrd6wt9jt15tscJk31zNLUsK7H8qysyeTccRjxlH1QJSHU3gcbkbiyLYuFcsE
g5+1g7XNM6gM8+yj0dIIPyO6CnRYIgTiZuuZp1leBKmAhCC5MiGoX8Y7+V49ZtJr
DFzhC+Ch3UZsB4MWevnsP/PQKtxd0CA93ibz+AGzhQY85RoqQDUpWbOVE4RcJWqO
EKs3YnvB1f10PvbB5yjpcfKfFShJyOP3cRcHbp3i+M1zEH0iLR6m46vem9Uq2kaM
u9Z5cNzedr0GXZ1TRz66szFhZL6tZrJEaW8375C25HflNLZpQWbzBM+i/pOaZdZ4
vIVE16JZAbGmAfdtANFxOUpgIUXXZPfyI60EV4CAWgOIqJk0IupkCrHlprCTx5gV
XQar1/AW2mhdmfDf1oDeF1RoGcDnGUxuHl3TPheDHyVvMO9RNBSWyBFdTdaoBL5T
TfKZvVz27Gwm4zChH052S8tQMaOSU9TpLACLAPoeIJaxP8gym3ThMJac+tzAWh/Z
xWiK8noIBWV57BsZw008ytaqd2I8gGWyFHsOiZeJP+f2Ev3EzdGt86csaxu8ZuOi
F7TM2KWYEu8es924qb3dK4NgCOeCKPN5Bj0sFGrN1dZWibmj8xqy8vjSvCSwT9j5
5Zh8tWDGs8G+2sr8qV/Ds7V6qJKtknsy+KUGDcLkAzg0izd8ujf4SDE0yzfH6CFk
lPS5evEAEsIWlEWvrjjnMWghOkG2R34iSLcxAWMdFb0pfB5kHp1tyhChpi5r4/uS
IPHP1yrbEZWxQr5QSFJGeG496WTzYKmhIw484p/5qpSarJV6iyVH9feMzSFrf+tt
gb3FAt5QY8iOSSBelgaQ1GLUIEsEpmYvHSpUCwUI8IYX/jv6oXBUD3m4hcNBr6dg
uk9F9aFoZ76J9KqsD+hvuXkSxyNwRkQoWj/YYUNwNNWdOGsUbQ13zZObaRja3qlb
08rtWhM/Zja6X21nmYH93/IZsr7BVsG2nZHR6eh2N7rQoQ0VMiwztTVHIrhWWfHi
jRRpnvQXv+E6krijszbxaeZEn+T73hs9bfGUANTR3grWkw41i6TnJuMWTXtg5V53
8UcCZhUS6rMEpU620ENYp2E7xcVk/nlSF4Y9khIJ04lWWvxgA6UF1t9hDXU5Z9Sm
nxqQMBMTJfFDgGhJw+FNHsGCK9AIuOV6QQsrJfgzSRNNrgMHA23KHJZ/n1KK9s71
D4jvv6mu+Mc/8q0jxoWvo/6ggYSIqEwylEduOGuIVvFnJCFIdlZ/5VVV5ljoZIr8
gdNuCTnalulfzkSRWF/YprZ3pboWcyWsMOtS+DMfKUBNpYQgZEnFcf1SOwqN9b4U
LesI3yV0AHM4TCs0Da+2vTcSKcLwyd4VRdUJxXneyb16IY8KYOtTTfN7iDLvcxEL
qqCU/yYsIxxhA3icw4d3SJVf0WgNkr94B5aFPw/b6IhNt6p49J5NpwMh+c2Kid+c
T1tnfeeTfHLa/OO7i87nfFIm3iej2Dr6y+ZfgVzf4e3wlA/8hc5/idyp0LlCMjfo
C77OiT9vIZ73pdXLQZ2rTja1fYnJ33okEmUz/eXmHYJZl5mDpKbCQKFVWKosFhOI
xrl6Dvk5u42gMRqEqEdZCJmKfB86nHzViX5q3UHTj+akfUYt7nJ37gshrbuyqxgZ
MTo4gek2x38bSDN1iEuQyL4cgiq9tDq/P5fZ77CYEj5uQxV+yuxrTffmTjBK0EDn
BiGlK7JwU8sWRn+d6Uyz/4nuDGCa+wl2IFMb5fosS9zCMOZx7YK8K/2Td0yrKG4w
JS+JRYSyelYXtwrH027dqIfceFdmPyEl6a4M/Uymy2YY6BeU08Ux5zJ3DdaqIPvC
JTrOLnGMYM4tGzNk8fdfOpTb0vut3BHOl4cWL1t9rR2rpBrAZV7ktbzcvtUTk3h/
ID85iTf9v+0139wSlKnCdNw13IUjh+ouvZlcUCMgMQOW4rRPp3CWJBZ4P84v8ts8
TZoC6Hz+qsF4UDMek3C8ebHwHjgykJ7TTcZ6v7oQELvdFKJ2+PolX/QVZvri3aer
Nwr9SspeYlSbvKRcNqV5x4GOXy2e3e01TmWUjdrczPYafNKW2tby0eoXADCXPOm9
UxV3SVOWgAX0K1pbKBwm0tRVfd7AcHy9kHYhwrc/w1hH51ORgAFczheqPTI0ksEd
YYL3JRyi1MQduWLuByRDEAlVGI8j5LldKLIAmA7cd/71agHWiL6jDj10e0JneSSE
DiiVm+rrakskxx+0CTWYaCG2KsyzZLW2ztaM+UN+gAZBucNxAprlPFTfueEMwsGc
pqZkfs76FXvpZf3fQM+t89cyxQzAE9I2+uLOzj/ORasT9pPONJEy3TIdw1cVKesl
7rk3/ctkDArPYxkzVFKdKDmah0nDygGGJtLgJ6IXUWChzyv9zjfde6OeiJ5GQYRQ
/b94B64lo16/dIsugYmm49FEUTiE6C6TYwi6gnNtTJji7MKlpETcydhfxSGqgjKJ
8L+uUHERHBx7qm6cDDsskTkNIwoX2ksG7Nv8O4U2JxUiOwqCV0CXR2XN+NjO9hKP
+ReGqSXsw328uVdXMcc5ciArZ8GlFozafu+h9igz3c0HucfPUViu0gc/Sw1V/RjV
RbnvujbvwNFeQNm6Rl3Pu6uIYfwmyOXDeu6rIFzWZBikzpU6SQhvrvxGf6PC0JnW
PRbJhkAP6R/OjnSdkj3WN1MVbhxXoP1W1REjWJRb4qPmccLnGSvN9ZvwDWG1gZIB
cOPq502oloSPV4SMcbwJD5OKw23BvNeUNO3g8YCDiIPZzSm+hIlUZ0Et6MPFyTla
wFC7T3vEAFhvswcnAS3X/TYWzxpOTyizn8xnJ+iZm9t6QqYG79qsbm0yN3wrvNTX
IfyQzSDtc03XnT4xjtFRjrIAmMOtfqvSMLzLlE4DYLG3Q+qm/wVBtcJs/8zmeVkM
p3F1GAafTZzrDsdNKJCKkKtTdBVQO5CZBx3j4AGY9s8QpxN7Y7qnAobiOCjI+zjx
BJYvuRnVitGRrVYzwHjMVo2UEq6bLNamC1xX3AU42htpJvrBzKtIbA8pyPx2AP+u
7zc5BNKsMar/nJqicJjv5wEz/1fxu7ncSMt53nMH4VgNLfejBpUyEkRKEiwt/nx/
zbbmIWUH6LbFxh6uUsd0J4z1sWGZ04AqF+esB6IN66VBSEVlSp7uystxYqmMtqFm
ZCHVx0iCrFjKazjP0kV/8PkyBJAMpaC01UZckNPXkP3sQ/tQxwnHk4btrHfx/F2a
h8l0ZvtJBKZVGedtULyx53a3N3RqX5XhNj03dyctoxJX6EM+gewOa9A0AAwxGpzc
x3/bySjLTvXYQPVEEKNnRHPkrO/vVjpwpwDXPaSLLU/S08FUN+Hnoc2MAgiXeoHS
nYADgKmJKTdEzi/IR7jCs/6djgoF9XcUDFHymzQelp6QevZvOHwrof+ck4lUa/P1
WzIjgIB7tTpnz3w+Gu0OycgbVIDb7/4hqtSchNEux3x7dqT23Wuix2ABmk6jQcaI
UJW1cheKFXM4rwge9Ragd0lMYLIjZcLexGD8ERkuXPZuG3sOIy9ebiRg8D23fHkS
UsjGTQj8E0z9NxQfV6xnjjEjHaWU/WK565ddAEgHYHxD2Zlzq55HX44BgTBw74X2
m1EAmn2r9lHmYw4Yi2oO5PDEETCOlOStq7QEbX5m4SOK6QWokPHjr2rxa8HrU0Jk
WEPjjBv0aJlAbQdc005k8B7NEqCZ1Xy8T+sjNgmhRIxc8icE5xn1x/OmP5L5I4Yf
n8jdyadavbWfelXzk2c+f5OCElCBECEgzma43xVjVfHvPDXFP36A4bWlMIsT5DHE
sNM6FLCMx+JcUxLgweO1DDZzbxhEe8qknTpQw1rF/HcLhWRm4bO5ceW2atv2rH0W
oUufsWUqzw8JaAtfYeUUAVJXk+64goVrVgyvmtvFg/bZjyMraVUNyYJvNNRz3MXj
t2PqInWEHQsG31XgIva4cy65laYsPZKe7gkoqZO10fNOuMXdxZOgWvBN/be/OMWC
QpQW1jPj+j+8ZOa1vl0vjfjjH94qT74Ypcn9BeT5nP8nR4KL4Gyh2qYXiw1mwezO
Znq8MCLsPPpxkJ54x9HOaGXUJ3TfYGTwbg3ox2i6eWKStO1mRgCKyURpAxTcNwpA
s4amvEp+4q2OCXXY6wYTmcHGoPHyK+obJ0ZDklGUzkuL17HVREFSZ/St1/SNYiCj
q09WBgYWeL/th2Kz/6RF/G770OBFYyj2OXI4AGHvkRX4GiBLYYu//69Rsax4AFh/
BSr9mUdPtKh4Kd8no31TCqU55a8YmeFc5QXJvdPRBho7s78fWpiOPrivgF/9rCEw
PvJaZ37pQx3ZKSqSdDxYRhChFehjy1VbE4wkfLtutr54DW0PeMx4lT8hFnW5Bq8j
LYm2PMg9nt2BFD+tVXbEfPwPIvbRJrVQY6K7NwJ+xmM96JtuIn0I3qY44uT8kTjB
zeVJkX58d4Wb34WokLBhcg89vlARSS7i0Ny6Qgc6dYe4NOdA8sGOR/xloRdtB2r8
R6rg3s0F9UpzcsQYgyT3WYiqiCYf/J8TsBi1pdxvWw5lJeutsdSwhbxBlj0bBTeA
fWCwlnwJsSl47lUo/jzQPNsUgqPBChzR842qnF9K/M8Wi8KJ90R/KQD4y4bOfJzC
2pk6J1RfD39wY94oNNTtPPFcMirG3hFeNWI8sW5LE6i2tDa32caropW8ssM4O65Y
+quN3jf3s+QepSoH2Efzcd8bkQY3uOQygy7P1iFtxa+oe584GNP+clQSV8oCKS1v
TT/KhybDNsB46gqoiS7RxKAuOTgNlivUUpRV8s3yEiX4BVLzXZPsNTUdqjSH4gaS
Q3r5QQsf+T0z11MLtRLnVR/qQkI3hjQ2m+tZfurdtygE7r9zglJgj1yD+PnrPgcU
+t0gNnGfwfPegyW2UiWnHXW++LGiJdX5wyN81l4znUJQdLZf1di29awLr4equ7A9
o1px8AQWPYsDrOhYz/tEG8SrkrmYMiot/1vfpbqsGjUBfTYOrLdnP65A4qJO9Yky
LP6AhHiPS486fOaYFJf2Awri9Al3gxfbRv2wGbPMQ5sFweUk9+7a4tUKl3vFYrze
/DD9sKv7SOK6EuKYF20M0QT4AC8KASRuBnaOkvUlhk5LRVndcG7SEzqtCcxGI0Ar
c3dckVHG8HyWAlHaLGZffDopgWZbieBpWC4SrIWCO5lBjy/df1Hk8XqyTSNhLOZW
me+FY50946Kg/cDi3DKpFnyCTU/OMljCVjh2WZYzs6oorR9S2Mir1DIB7yDr86Yo
rCT+zonRgbTNuhrCDjcE7BiDVv8I0N/pAjfh6/Oc84Y81R1f0RWHX1y9ulmoc80V
gqpSPp6OFVRADI+1WNXqDDzc4dPRoR8za/0aZy/bYKhARtzM9eMBcHa+bxwMxyrc
762xYtess6rvomzdQiX2R9FjNzu/7g2mA8T7TXXbEeilDJrroKS36+FHCqoG7lDp
166M8NVFhvg6Rg+3tN+A9Y54g2mT+Bif9xHTqCavZ+tJpwAxokqiiSfRVqolWAvo
wSmfX88HTWZmXjTBfAxVQQwewvB6yvnq71hsFv/554EC/+YvCep9kJ9M0/0jOVxg
YbZfexl0kvuApk+s87tQpIdQ51BYJISQx2/ELvo4ioqenbSBynJQJRS8B/+wO+mJ
qLR6kwj6Gs9wNVpvxQ7bhI1nlEmYmml/nKo2ugOFPUt10ZnLo6MvYqXiQvyn9X9+
q0JYPyrY5i/dQ3IwShBRqi3SoZGEUjEGk49lq9d6RlGi/lY/IdBmehF39XMXmJAH
BfAagNtOfah6XhnCLR9fQi0rIXcrz/FQdqIIdAghSt4i+p++9bxe1+QMlBPlGjqW
7S17Ab7GIveqnMK65r7Z9iMgCuHKWOdU+tS1ukJmTzJ12id58i0bcOTZdLKpbl7W
4rQ0P7ubOpoz4pWB2mPZExfzyEbXhjGncMJolZwOdVJp9uqcNmlbdmhtmEaZHo7e
GKAQ3A1TNv56H3Vxaw++r9QO6z/1p6NjnBxyrK2RX7yQfoAKZ+wSBZcBNH7tWhEC
ZOVDAgP83uha+y7Md7HxSB464Z49x10Cm/TJRcKxghV3x6LG24aD5qq5Xs4EPL8Q
EuwFGYEW9NiiD/PYq0KNr1QGCUarnSvAYHWmbBhvzJdUeP3r59dX6Gs3XaRCtdrP
M3w7maS6ZJJJSB2dsG0Bi6KEUGjfZCovVXBdy1Jtp02O0jusRAmVYBg3vpjbzh82
ysGuYCzlzR+n8W1/HglGGTUgOwPOC0V31i3Ld7C3aPo9FB+wo4N5TDI7Wcrm1qu9
9Wvwu53SClVJXQlz+y4+SWPTB5WlNZhh8EJFVoD8AzRzcCE5XPVlpQyIRqOYIkQI
hTGTuqQO/hYE/flSRF6MJICsKFJYDFOgRYIM2xEJxq1EGnSy7H3OoiP+IMHxK8Qt
6fRR17H0xLF0eH4LK6obpgY3C7UnO6EXNR9stiHCUcKDgRMCObZUpJFhr3J10+gJ
Sk1c231wagA0q2FS1yjLNdsId5fr807AkvAL6KxNPhD7jWU9vLxNKTZARIA0xp3y
vXkbFeRBWH2LJ+wzAnhmfp5h+u+ItDh8v0U1SiJbw3AgpY4BuPAYDSlYf4SvsICk
8kXBTHNobWGFicprKxaYbajj+6cAfRYDHRjFGpYptmtucUQ0ySsDyxKIfHreSiHy
WEvozi0pzrsdFGtKtDp8BvW+LP9WG4tDJ1MurJ0G9YPQJeyWY06eIN7l0ToO1blK
HdfL0deICbbLO0udNKg0kHwAsDMm2Hb0BmRxVNLSs6lrM3G+er3GJUAZ3mJJccSh
SsorZFXShJ/3tlALJJqXorxuTaMxFScQsUiTNg01Zck/eINtOCAfZIVwHQ/R+uME
6vaiv6CWYxRgJoJjETJXhcwUzLHo8CT25y1Qil52Q1kGYiQcdRXLNH5UC3VW9ABx
IFj2QXz7klgKilVqnlJ7wTBkZM5PBKQQZC0QshDgEGJronnmuSpz4ml39YOX3UXu
3qePTdCZQYcVW2bqes8hUnsbWXxX8NWGh89KG7U6naSH73V9E1c6/xqrkGmpCcA1
usY3d1MIoEy/4NWAmNY1ckoFHkUBAywB9UW3cURGBe6Pcu5SAcOOPoDEvE/7lnd6
P2CeSdCzDQD3BLMJYaqxlYsv0UQIx1FENOa9PXstpG/O+DY+79qfafnkF2Zb9jnN
wlw5ENPamEkvRUOo2s4nrWr0WQ65nJXVQnGKZdIAyAMUuHmWDHRE7a2slo7EJrbJ
hWX6IsSM/L7vyhCOa5YCC+qorolmMTzq8zhVXt57kSxLiBV+bYsppr8+pwdRbg50
iyVAB8ocK6PY1RGlDBs3O4HZxVHiAwJD18vvnMeRKF304URBaoLWGM8O0tNMSp+6
aSvr4gDJ3xoDB2j7OK6d9tJFZeiylIgdfJoLtgl2mAOPp4eJ3x1hEjY6Y51NfLb/
WDaelS/QAI4BLIgC0JUXZS78b/5gudbMjsPQi8K2f86btnsJcAJEzubcvcpCP7K5
3WEd1AX6UfIpUfgogYOIXGRfZWQvrbYNxy7sLkWg7iMyH6sigjUy5IKs7T6B62Q8
SDkkqhNiFVvtXNQc82c3IH55lKr03GPhuyRtrJIJ7Brw9LSlAu9a5hkbiAbR6tFX
F3O5MmiuV2YpBwT0tOYRSuXIf2XLHv32oDUj4qmmQUkWdW9rOmudPo2ncWEteabI
MsjWRaq5oK/otFHso7vHyiKXUQxm0khnCH+9jC3blCcucL8GE3F9nC4oLcKpTTGg
O839Z3j2gnOXVZYjTsd3MIluTyYpBwHHbxPA4WNctzbgvyM+297qzbRPyFM4Z/7L
W8GS5zsSj4pQdJP4T2I7H7f2D8tpQmTeuRAUGY6OquwQ+CsQ76sBqVoB0zeLG0/w
nYYJHIQIYsbgU47E8zrRgax4TKi0A1YBvKN/PlRGqjPwb3xMSNZ9g5HdVj1HxhrU
+E7mRGddZnSw9L+AY3ZvCnqFRBza2mAoJmtFckQhlwgRuIjtSd5z6oeJV+oK+Ecy
4a/ff1EQ0UQWSumQdj6pgBDbbLamShXl781E7+hx+PjLlewbHS+IireEmRsql8AH
ulOkAY6SvYetja0jPSsXhqFli3vRLZ/FzFXFYPZ386YVziU30vB9wyG5EigqPyiY
Pt0jImICdfOdL0VBOptKAQnrKvtFbXjwkWnug4p198BthutocDKk5XoohNKX2yI6
VORoDw3f+gFqxnhTTaawSR3MaWXHRII1KDSAk9yglxAO/pWlBbEwgbbraShVW60a
m2BM6alKpRiRQ/+4SErAaY7Af1uyU2S4Xv0+VVLYrMWfWFYpGSZWlJ/hGzdmsyDy
k4oT+75nqAJBHwP5Wnj9h+iEyg7ZLMXzHe4UCmCATvGN1FGO4wgXRz2LNP3xc/DC
DW+kuSeR39wcHcYj+R8yqJGefN1cqx9kZzfDDDTm78E7a8xhZHBqUsu2OEXGFn8O
BO2eg9wlqJDGrICA0svsYQ6QJSYEvjergqUYyb8QEqT2Wki9pwsCoso8HSM0Aw4m
ERFQrV6iAlHrtqy46AClRVeHWbHYc6O0Tk4QqFLdRARuZNFM3Q04rBNbJCF/6nCq
bl26kEq+FI1FcL8qzsodqZBcFuPY0wt+U94gyR0jVKWVqTeWfhoASfw6pQC3jH71
Q1X2+oWzJKXGk2vcgFVXv2fRfaYfgR11kAaFL6MToOfI9y0G/GaFMLZzVPKdUD/F
I+dncONbSHMplGJXDCzcuvYT+XWRq3t/v1hD5VTOGCfjnnV0avAHIlbG2offGC1J
xtRr4nmOKTNCXZYd4FkZaug1X9HNUiCPa13e5OZK1vriD41k8IwL+mkeI3WG3M67
NLpAPNCwFepU2p2l1ELNo80UDzlANmkrUHF4gjvzJGLgHGkiuYMcyJ7XcvaHRItG
+91r0vukdwRBCSbVccZfCnkNxHfnlI26pU/FAHyR8sJAIkt09kcBroieDaKKuNNV
pGLBnIO+d7iVcY9OFI6uS/G9mOXyNQ2PcvuUHgABL4Ij939EDREY97uZdYrw+z5o
Oc6FXn5w8KAZd/eWT+GxzRhXxi+wpSIYVwfR9VOjQu1fsHga5Dm0NkiTXSQM9gkL
5rZTSitVBK1ZAM/Nd6B5rJnPqwlAfcrVPm8cijD3sZrdOgipaXP4QyeH5gXwgXj/
uZiAWQFYIO//o+PP7T3OUYHrBCSkI1xx+DWUHtXRVrLbMYtjG8gmcCCUGcElSdSK
ejRsTNi5hcMJpQFjcNDtlIwn543nc6oZFTzjybaTmdI90VGmg6Zgjdlub0Q22XdZ
7NQBW31mO4N3URyEJhEGF/s1KoiAFsN/DpRjK7pRy0OlgUrcUe67QJIHOUZFym/F
KzUtWgC8g4a6Djnra+DH2KPhEn7j+/1SwysR6ojDn4w5+AUurnGwPf/07c06/Vv7
4sdhQ2PSM5p1kSDv6NXRZ4Wed385GaVDNyO1BO553BUkklKceElABukaYnIOv7DN
2Uu/oDEDn71+Lt3CUZjqkAydEVU8vRL/lTX9IbE8bE+USBpotVFxR/jbI4SDO5TY
lYvzK8d8oULB1tC+KW0sk1R1su36ad7SFmMIheW2M3DNvptuTSPZhDHDDBJT4LXF
JlkjWu4uUOVbNcumCuoitudT91cu3dmaLs/LMSImEI+IObKOllNMPrHrMhNtwSCq
qVb/28gCYGLShxkWYGDMl2RGls0gb6F7nqWH2tub7su9zSntKAcuTSQiGMSeZJTp
gUyoEknfZK3LHSyNxWSPqhwJFulG1Y4QWsnsNius0AxVCPS8n2V4vU67Jg4S/X2q
uIENm03a4k1jjznb8hR3ur6OGKqfjbs9Yp2fwVJL3pnxajmYW4F5i24yA5o/hBEz
jpVmTHe2Pnq9gRD5irPoohOkrSWjeA3Dem1kIwpnz4GobrYhNLzCRASrWhrIxcBi
SI7s5hGy4Rj9HCDZK4utCYB+ws+juSnmEprUe5Pm+36MRHOIXLclufLOrUxKp37U
1k5HHkFbrxPFZUe+tixchxCEUEIoubBii4g5Z/znQXK4H4amwu+wjnW4dxuNYiy0
SACXDQ73vUQPORdtepKT39H9ljjQNQqu4BlUfgokgq7iF5Z8ldZq7PVMcwbipz/V
bMYC4dG4Js6CqIPTqb1CiCGpDHx8W/WwFHJjQYhODjImkzvPrmwyNl5BO/N/EYcp
mJp33vGnNEOe3spGBhmizT1eMf/xIhTmtJVjjrYYAkjxVaOOu2QSAZfOzW4QnvAp
IToQvJ3RWjQVWO8sRCoZ3mL8YuZM5kk7zFMcwNMsPfHPu7L5nI8eh9zU2S32yU4T
hdXxocrWscdE+/5eFfIe0SdbIrbkjek7mz5yIaJjVHABHSlbuVZuR7XnfeOK2nsx
SFzliwYU7MV0V050xTKBPWEKmXN3ZmH8XWRuhwogGYMkD3W/qAiyS9LuN+S13ZJ0
l5cXxtF0adQHrlQBigUe8jYk8c6BQpYSqBX51bE95/fPcQaVWgxPGbhA13OkpLlI
Vf7zhs82/sJKJTqA5eFgl/vQ7aEAYOmWp+YZS9/Yb1OI2apEbIgej6z2o9OOlv8Y
ICAA7LkjujHUkuDX2bYF0l/FBLq+2twuPmm5gNCtMMLIGOztXElMub6SME15yUM3
nsd33tzJgSDzxtoeXRGh6YhAmgaRbZJwq6cECM5w+hrrsQphrwm/9p6EYNrE1oQJ
lPlZg2BWLjYpDso8YZ5eJF+gcLHNVfay98CkF9+vWoaI9O7dRZoVpFqy8PDbz0My
IX4m+j9yxREQQyAmfvy9DCVFBdmnpfadGH3hh4ptXVXD3jIQOezsP1e/2acIYOhY
lK6kCNl2v3aqD4pTd6G3wcQl5vGobKek6lM7nqc+n9omJbnLJH9SQWsZ3cNubBWC
TdhoQxHX5QYuK3eTJJv0Bw6NDpg6DQiaXbV/X0kJS9oDm8QO7MVjL2aC0Jd1lk1f
7hXT/he6spOKPTE1EN5serfsk1jUqbRPvrpcT2WN5BA080mMdDA6HnTqnH63BgZl
kjKd1tjetyQHfhjzOXiGZ0ysqsqz8jmUmgaVePO6tDjxetVC2xNuQ55oUFutrPrw
JDr1xx1YoucSto9yDhJ9zh0i57fbfU2r0xMZg1LDEAHU2uqiO6iR1MtloSC7hzdc
1lUL2gHMtWLCwqicUjg1+Iw9pyq0slLdSHIvkjMSY2RSjnnHJ98/CWCE2u9YWNdb
4zZt800mspAM9FLY0mM3agFC82w1o/Jct+J8UKKLGUwsIrCab0bIbNtQ62zt+rJd
WMduDQPMIc7hus7gfgJWLOXcvbWqPRlWYQlqqcUEpam1+CNpImxltOBC14YQpstr
/n4bF3u34g61AJROitsY0kOkT6I0DjRyETmd0r++alTt+rXg4tsG5o2nzvbXMSu7
P4jp+I++R52ssKUACWVY0IdtxD4AaTuNcJAfhXfAzmaqyOsQg/y69ypDFPrISXGc
pjUMsH5NHQ/ZgUeewNIvZjDAsNFqxsLsq7zVffads2ul6Kyr+1SYvXtNKb/yOyLB
5slyg5c6gluNu16LT5FX69IC0dGM7dm1F11kyB8gqICnsSJugiLqmcRAVrKHVZn7
DDTLfqwLdm04uju2Xo+3iMkjkCyT2qasPpiMtoP+8S57LP7qvHf4w7GXepnWzLm3
wPSqH4G1DwAmw12v9doMrWP6oGH363/6FFqdz7YtsdiieGG06mC1GQOyN425m6bk
2A3b9BcH0caH3z8Y1kaxS6tvgNaZlBzpFiclEv4wZz/6A0ipiIO7H4V1S6MrhoIt
7DW3XPNBdPUCWyJsJ8+GGkgn/Fgi/188EzL4IXX3b+va995qwEQFopcSokmTOcbw
GfA/0IeaLIkIQJo2+2HlJQ7rG5Be/NRuXpZDWf8WJWmNzzmZMuh/8uBpbhhnmwOb
J1+BpvyMTuf6u/mPJuzqANQ4ScNrXHVyK6h1J9+ONIiH9SfWudODVQ14lDCzALBA
Zal9OXitZVc4zJqr3H3jVm77KACrq5C7AxWvUqYAMCad3SCEKUtndaVjAkOl0MyO
D9u9WSJhkrKd7NqEbdJGJ+FcEEm2AQ0/2YIv13UBdZq1GN5vtwTFeZRvKvf838Da
Laot/MR84Vr4Gc0rxNaBXDPGHgSlxYLY/M1sebtgLTLl4gyMYZIDKCsx8GMg87/R
bcyC0DuPBVlEBH6p9m54G7O4Dzi21hEm9EfsnxkbUhFpochuhWJ+BBN5RPyVLkjs
5zRlOH21C+B+ups6AT5TEH8WF/yC7sCSri4rHKhU6lp0rBEU8bfufdddab8EMl5i
PbqmqcNN5JEIcUEm5zgPY9i9zeq0hSP/b8ogg+0ZaZqtRUgQQ085TOigtBP2cvbw
Toze5BnH4OgjgSuHSntDqk8hKeRoILY7eCupfFmRIqNkWOa36oXcGzfJS7RFZp2t
fvJrz2KDwGOtqWMXSxpdK4w1vGcyTG9++BP+V3DXveUV/9XsNFZCRFnBad10hF8U
POPPiMkeUQxzmWzU7e5EhCFxE/fOD+iGtB8fyJAJ3Debff+oObiKdSKNNh4EDwZj
T2Wb97N2L6tCTu53t2Eg6evInunBZ0/n94e+71LzHZp9sKfm1ebcChq3FloJbbts
Fevp/bi4H8AzrncO6rPoXf28ZD+8oiXukNeFFjTrnIMisaakXnE3Agf6PtsckLVe
612MtNPkvB9j7O/YukRQdRaS8alYcP5y1Zz2zJ/NowWbTRW7lTv6QZV5vhY8hgef
mBit4zmWm5g1EEnxsq+ZDq0luvqw9q/YQ2D4oP1eRbaA2780kLapKDc+VOHhkf3c
cSrGhPXMC3+1nX2AWkvsHLzszhj88SgIhOqj6CqpB/v9+PdKz53qwECguOYqg1AN
cIKnJHNFj6AlLGj5CfSzKtKzE3aEsppa9+YynbZFsqQ+2uTrPkvdhAveGqXKZtFP
Av8dgJmBOmle7UJojzosLF5AGO7tje3rGUdx2QE1uwH5NkAH37spblmTH2n0gK63
1OLh6iZSeXIUQYVNMkiwyAhapmfcrURlvVc+KsepmyjWTupdCY0xWKzxyWERDY1o
5oHXLzalh5QG97TVVL7d0cc5sO+MvPQb0TZIrYPfbftBzHOIbilJMv1OA2753/k2
pZpAzpZHsxnJ3lYFr2wtX3CBeecJVBBsyEWBtU7uX1nNWK6iMSFKvUkNpJcNeeox
WBghHp6qgVHGqXVpbZtMACUzXYgiBO6P0rpwhgHcl049xAnhd3hzptqQ7hlk7Uc5
ijAmaDuNryr5863Y5EKK0RcaPPwqL2dDsGvtH8lkbzTqVu0f6ZvkRXP5WAdd1jw8
MspxCPOJy4ShKQEkKt70QT80BoXhn9u0qCfYXvIiU4cIWDdglwZXaOuKMChWG156
O6xpwjnGUFxFjY/+McNBzzXtquwRGayNADoRCqt7GOLgbLLRr38wFCdlLeX0aB/N
JvCa4apAs4aqQi4sFpzziCcuub+hKSzx2rgJj2TvHQEz4/uKYVlg4gbTCizOqQed
8WRB+tgvAsVY4xYH2aNScp/+C3ydmGzu6w6EswmGfn2O8lRdYNhG/4YFzEodWegj
RfqaUJ2cddbeCeGCiqa/Kb6wNOymhNVMzP4ph9LsjQFdbZXj5WS6D4sBZW9sNwEc
aFIsX/lpaTuYtcL6a1P5k1nVOp0VGhjlfwFnxQNNxqJCAo9qGnBT9PcyaJiT5MK7
AzQbOxCtR7WXuO9DSGcgAmr5xU6AC2HFjIJAgULKtmJMVYfbPJCeOgPSWCZfk+eJ
4EMR5CpIymnKkssMV/6VM0GH46Nnw7EKL6kLiomkP+ThtkrIfLpQ9mKSBQaMEndv
IVQMuz0hO3w4HqkBXU1FJajFX4WxKCJncEKRY7m81eL3PxQW1R6ocpJNNbutdWC5
MOyBQctVHc4ISeW+6umrSlp2jBTNvK1xptoX6ioMls8NwoZEfoelpG9jzBDSnLGt
hTdS6Z1rNbhC0vEMNSHd3X1VMNw8Irb+IcByCQ1WY8judVVM/eZPhAABWaJWjTuL
HJDydWuVQioZ5zlnvW7YPiWq85wc7/ksXbiTxXzw4UYripUryOA3CDkuJfYqYoOs
Wyjs6B6vp4xrrntowjDTjnb+Pt1XAIz5BidGaZzYztmDoFhYwAdSErmCdTGgV0ZL
hxK43EalhMnyQToqaW7O9V9BYpVgApdRDlxfy9cC3NmWWk1v6aRy8hlaVtnRS+dQ
Xl65jtxEBfvZnEi2SbLNizp9oJcuzaLN8sK1n1hqQ0usHakc+hkB3w4oVgcQZ4tY
Zx2CLdRZ/RpGlw2K9JWo1HhM+USJa0kaU3lwd+6YCsMAACFTpVcdAZHcQcquN8g5
XCR8c2+ijtCrRz/8Qqb1p16W5yreelwu9z0t6dJtObCkEQpqtuOTa5MLv81zdCaA
OZ1yfuNJ0yEOSfH/m60AJkmlHxMKKolA1nC5KlrYqUemGn+Wu/CRLi55yj9dekWt
GptN2+iK20GG2bAZBEJ+U2CenzKP9s177MAJB3+SQ5eyuJ+Vt6vcoM4eb09paQ8I
HpfThZnR/TiyPYdLDd/g8ojt0s8nIf8VVC4hX/XHLGzSwSfDOZYErvGBTy3wb+C6
I//ooKKh4PMl7MMVMKFJZnlBqnnylktu7uYo4NcjsYClrXKLCd82SnR0a8w+qcYt
kdRN3FfIUt2Rh/m6fQ17JUOqEc5QR6s0uqe3JQOYxDIx8GvKSe3IyZeXYG9xKRhA
qX6kxChMStAhN6R3XgvfvbIMlAJeG+e1GvdeC3E7xNY8/r8ECAKtVswrJ2BUhuXH
iWrBpmsA54LL/0B7xV0ezrVdB3VirwUd4A5IM4WPgyy3S/JfOX/S0M5yDQJmRLmD
lQ6d/ygBVpbk9LFP1S9WKeKzAHkoGJVmUhBvTP7fbeqlp/KAFFPV5FdtHp/2R3Ul
ZNzQxOLJSpH9rH/+NxacQQUBgCBpLgFqyJvntIzBaOcfH5Mchw8xGU8Udf7r/fuK
U7qqbIFtq+2s/qBpuv/tC6ro/FRd/ZTCXX8HW2BvSw9lQz1V+KGMRqPqHo3yKMfR
aKO0G/xiPF9P/2mM22KR+B2NhDH/ri0sf9ijxxEN4tjkMLrQP4OxgjlYKDFHnm+K
x/8Eg1IZYj9T421qNzaW+WBnOoBbckbKxuKqjj8aiI377KJ7Sk6cW3RWNV5AetIW
hL86mdTlj/KyNz7gokhvMY9Abl0wVyGBt1LyrwDT7IAZ4PkeuKriXcHP9x/G/7Uh
BrG2CrdWWzR7qHTURcEl54b082ZV2BEzWgGDpCt68bak7Lz5SsrYPdHCR84ceWNz
S9MhGgsK0cZ/sRSLGYUjczydsBE8TOqOPmwET6hWkorilY5RB+pwk9oqjb/0JyWt
6skl6ommRPbvE25NbZXB7M4bz6fv9/k3ZIRxL81lWhX3VIKU87fKAZr1SJc7VGHQ
QUTW3lSMAS/eud/H3jEMJVH74C9ayUQB3sAxdkvrzSgSQzXKMGVTYS11UMjF9oP2
TooABQ6KYIAxXhk99eGJLcet08K89ZljgbyuzWuycDDqt95GoSGu3zTQ0N4ZFPWs
x9JXXGEdBZ9u4Dr4Uvy82PzM87l4SBbCkPt9601OHxnSozqhG9kzUuhG4CH6P3qx
AzFCdEh7qVW1qxIJlxPKOc6HpbWCpZkxcj7Hp35lhO+NiH3kJg4B2NFyUOrqbG+2
CbZlEGiuM3m7FFrAY4pkLKbzuv1tgit+FioqBaTnwpXS9iVPJ0X1G8U/X9FkYQ6C
9rmkd0hWVyM7/zM41G2aBOhQorBslkBpAwRlAZTg3+f1bFM4CmYHP0mFSlZEFQ2f
/fa3EbiU+flo/pTVI1zOI2IQItgxaLg+ALfx2DASlI+Q74xQVLS0hcao+pTtWScH
y+TCJI85OrjCRUIT4JhuWT0Z7cD8htQUsxjXLhHa4d1IvZWtXYLIAUd2CngyufRO
vOymZ6CogGuhXbc8nb7dhxhrfwbX0G2+vfEZJ1JlocicBzHnjr5xBGj4bt8kAGk5
Hiu1JQ3SekUkHADoaKqJzI7mx41iIylmUurzWCoBVj08uc7mcSQgip2x64DbYfjJ
JT7uBHVw/Fkr4NMFSQKF8xneA1hG2cfI6vOedAsEKbCZJe2xSNumNOrR2wCxMiHt
eYTw2MMOCQD5ozOZE+L2sozajAW6ZyeVlNZGHmOFGHrI2xBMHvhERv2jAYN16FRP
556cR8MF4FOOjnczgl83/Gb5m99YdIF2alL9gvEC/zUI8gvQUFq5XTEkvPNxn1JE
x4Z4R2LHNiUjO3Ci9wsaBXjEcQTzP2MirDvfKhpY5ZsgtcGBcGyol3+4ijthSDjm
EDC+jivZgorsMdvjZ88C/m6SzcinB1tA7AGH3/uwpVocNmUnF6yuLOgnkwnvQP/F
jsSBGhnak90EPYYJYg2SkpuWApK4a/JhfhOZ62q8CFWt/yuQZIVLz3+LMBwtYlNM
8cUZAMq/lGHi24GZV+E+Cths+D+5FkJcXUZk76MJ+gupNjOj7xYhu7COeyV8yq1T
T6iUSx6jtjpclqh9Dzgqgjwo37QlELm7JewGmJp6+DoxWu9mmeWi3fyH1A0+wUE3
XolGdyUHzC+S7H25C2VCd0LR7OSaPKsIIEtaK0CfdpQ+40TKTnTs1twmjw64UaNz
dILcsBHolwK8NnsBiymw8qcgmQAf2gluIKNWWE9APt7HPSSxP1FN4fYfH9BuqaHf
8kg1S9I590IpI/rJeaRbhKHayzpyb0dXy4NLPX5vr6sACor9mkpfIN4n3CTdn8LJ
6Drckzu/qtZSBK3YsTXQnDeOj0vx+IgDAaU1GeKJOxaZBXyJdy5jNajAbM0BlkGG
/tuFOQOlVSbD4Zm/Sdtaco7m30CCMr3W8nqZYDOU23vllcfPLhAfIj10uj9nTkyi
ZAIcbzW7ptkexrTcBAfoWg6cpKwbOyH6IhtTdGPtbk1YXpTRKzOfhjTFJ+zAkCHX
iytXxTNWBo5KVOt8TwLcMNg+fPQvnCai2MW40ZVGs+U6mtTO6CPw6o5lZBPETrIW
gPwevAg5Mj7fhOJ9A8ZSpdGooSzHAqTRetjXjTpQlTFFg8X6zIwq2FiiG6AFgOdZ
uBEqJ8WVcVH316YJ/qpg4VEMRMDIHcCC5AV92G97mgLPsRyafoGNxzB/z6BDhI0Q
64fASJtZ+S6G8BZWtDzvhGJbh4e1FnbwsO0mWBokpeaTqXUGw51vJHWYIBDhX7ts
tVY8JZjAznMXecWZINZe1Q8otmH+BorqGEd+xnJu7EYK0borwHyiUa3/mM+vTXTv
/Vk6dFZNCm7pnnuRdu/Jq8w8ru9AJrqJiCM/i2Tgfu7DM/5xeGxaMqs5gKR11v7n
/kCMGoRLqOKkRMU2zJABH1y80wuRgmqJNotrr7pMjGpVj8uZj54pq4Dq9JsPk44O
Z5ZBeoTdnsTqZzwpcDl5gKrYgY7VDoYI7opHonzzyXXpsUn1KIKUbTdP/L3xoWHs
wnruhLE3n3531Q8iBZpb7dOVzmMn2zVBlqvn0Q7iwlWIM5yAR1IgMYEg4PrvfmoZ
ymBB1bWKaN/zZJwhy1pcjHIq8LnQpzIcpJE+O2DSkgetxOmwsfCAokbepnk5eYfJ
N0T0X+0ZDKgDekjHZySAKbsmY7LHErXg5UF8ww1TG5/pLrawZrBihbnSFLeQqmlV
FHHtdWSVdhIWfU5bC/0K3Xn5Uj4TS+pupXkwRXRPVh499+FmWjleaPmJWeMxYK9G
TipCf1eHjez0lB2YxKuN7NfHqXHZ+FZV2yc321Q4C8LOX46Vmg1Z/pKgM9iTUkhR
IibO/HgUQKHQJhaaG7ErNZWSBcS0OanjPtytjVtP3hOY6xt5UU6NBLzQbD7eNY4j
Mg70SJKgvLPTElVZSuoxj2ILguDtBv7ZspoTGPdnjhukauJFjClNxwFX1GtB9uLn
weXZzDn9RRB4SANHKHV1h32VJA/4HMs2voPsc323xGPd8+afLl5KEYdzbUistrSL
drXfQAup0bWYfl18Vq25PE4QOYoBcKvDlJvuHMl2IaGUeLi2OHNHLmojeiuVZ4JT
MdFaY3ltDUGZm66kOgRJT9N9KDXBo4iErnTtdIW3PHdpbR+ydlNAilmIglNyobQF
NbWviQXeUmg8j5k9grdhipacIkMKhWjUc8tzGe8dVcZaNuibEZJHydYbkAohLXQW
05n4WiAZTbSVX2K5bgFQymhh0EKkLdq7zFKJEhFFH7Koyia45bW6uYCPSFwguBXy
LE85byFwsupD4v+tk7ZWHVbTXbCA4pI6VPzemU/PZmsy6Eh4uQeqLObMpVDXwemx
pwUXSz2K0emqEm7w2J/RF5fXoPDXGJqVA87XPOwyNYilwGxcyBHesW8wlVSuIubh
GPNyuoc0FjmSNiwgr+j+7VzfWOSi53q8o0JX/HgYMVR6UFj9PdhRKK4ezq5vEau+
z8w8B+zWIC/zhqtlJGKsl7KZOuU7vTWph/BIBQez0KwY+uK14ujghfHw1hPTAqR3
qVayGPU+O1Rs/vQXty2XscP5ZptpX2NTZgdO5qcKA5nCvOIGpM6ykG8SavTT/Yl4
r8O/iHJec2UsHGtCbn3crZRgurpFnXXP08NxQ4AT70Kjw7DYRQiUI9DGILS3SpbE
vHx84ZP2Hu5vKIi31HqFsYZtdcierSRDaATRBlNOMfUKVD/01cJ9igVGKTsTCDRV
QUO6vwtuf9IKXL/FskppRtNCsHqI7T10TAZffY0le/cLWq5S3Kbh08YuidK/Runs
tbVdRzl1FnbYYxhqaBSV27qivldY9wv+FisrQSvYLEagrxwNSlB2/S7wLayOWwKL
DNSaKGEFHdG9H4gISnU26tJnDMWtlqSkjCMBvDFkL+QGi8vRqRAxmYt/I7dCXo26
9fQ/ovW/b1QKJas/7QXW96dUkCmXydMW96A9/xQsxNo/2SYpBILE5j+uDVVpa4TG
mA0nsOnuIgTHBWc7FI2zlirbWpK2kGl0mpULR8Q3/r5wtGhfWGLZvJLE2tUMFrCg
2p3tViojv+p7BqOwObGWfwoiuyZ4OH7W4JqlpMyibMTB8858wJO5LBnR3ELNOGtU
g0hX+cLVxniB89eN4PchEYZu2ykY6Z9m9SIo2Ncp3+EGHrP+EY7cIYSfVZYOfxUX
uOuuuMZFTeW/vArr5HnE3QNPThdggXCOPgXrZpssq4AzcOsJIfp3ZONk9VOsZ3I8
xzMsiAylxhJLLVvwl7ymK74ZlmvELv/ITeU54cn7dHxlZX034Tg3dudGvBA7VIAg
TTHLoo7oAuvwWMZYUG+qo3NvrQsEwHZJZNfRpDRYLB0Fz1W0/tH6YJnDLxU3zy4n
X7nBhfTXGgM770hgjmuILmVpWCiuVKCESCE3AsbWNtsq76eqz2r7Z5BvED0KAzCU
gbjcEuORN3o8kLO1nVBCyZyEWkh5nUVrafd6Bc0w7Ouke+FnWhUS5FuoZr6coeeF
CQekgoIGOTsTLSMphiL+CehFEJYZKVgrIfyeSvfAtiS36n1UHKpzin4drStAFN7t
F0qgYESiuN/x/3LpUnQXcQQRxZppErJzwrI6mFtZYzfmiKWC57/M7IMXJHCilTvN
zvVj9+uybP+jKp60S/mUjAX5tcuHCZUrJU4bvAp2dK8/0pcBjd/ooLwswYY5e67s
slpLRUEI1VB1iZKYwWzYs21O/hNWnSkcNeob+QRf/2zyj5XBCFbbIG6EtvkZ5vHa
I07BG0p1qyxRl0xBWEWR3qU3eR4GXxPXFpRcdBquxByC4YlDDipq03Zeb46D+Ffs
hBNrRWhjqk2WKUCoWKoAVnnk2cLFpNnhXwECO363XwaDh4E7jEGgdfRcAex2lanT
DYiY9EBDR3S5DqRIFiOM/1kc9W6nB0PuceLE9FBtxQ6QjbRqvLUQT7RnW0Cdp/Qd
3i4mwpyjNwI19E9IywtqoK2pApvLy+Xqi5t0YFTHi5DKzWWRe6djW9q7gNBZMmhp
MpvsfSP/iuksv7nXlpgHVqo4BVrt6bM2VwsZRQIMEr7mxHWgyJ4IcwfXIPmKqP/W
sOy3TN1QhDobU3UtT3XP2yBJAmmwFIMwADGGlu1xkAkFcUkPh4ARTGBv4uWqKrZo
CBlMHTm5PhY16Xvl7r0QNHkX2JlGmg+kdixgsMb8va8XQj3+L7HdjVvAIDzaagKY
uRmkl0K1ZhVJiue4jSGQ5ArBJkpnG99uZOzgMcAbaNIgmxxfqx/Fo6qi3d+jZNKs
iV1jO19tD8YRCQYX6SB6wQc2nWCfP0Op3JOKzgItj1PbVgyVhfziIkcSYBQ815R7
SQJj0t3tIJVuRTrJnhKh69A4dJmg5PsnMK1YQsmEvET1x0RALPRvKkZDwIbAFRGU
NcD4fybk57DrCLPO9J45X/5TNPhzzS2e/FioPYYTW+EZ0CSxVJvTPRdjSGP5/KP/
IMyYDJyyIV/v0py/rMxmVFF34QYi9IcYlI+ecZM83ITjPIJfoiECDj3xeeYTTXwy
v5bSM1gkInNiBERljLuCBZEVKWnU/SsfFdcgr+rlVZE54JJWaFcmHDEDV5Rracfd
0Qpk93h96NKHAeRmPCY0tNk2X3yfo6zdovYHkdC0A1j6Jl7+RWqxTf3965Fs/b9X
BvDv8Jqm4dvjoTNh7IEVl877lFYI2yAli0NdPNnKPi0pYOZ2+9SRA8juLI8h30QM
8aXfJJK9GQoLZay3ufqe3lVBiMVPYwIz1MYBc1wuh1AFbAFHARzsgpexozian9no
5lJm9LbLDE4hzoBKHjNtCb/ku6jUa6fsBbCqkj1cunl1JyBdhPb0N3q3WH9Dif+7
g/d4bFPKvc8SudXyvxn5M0MyYQ5Z5JrvCg7hIBJd0hBVZ5Mb56ygT0zhS8+T2bLZ
fxn7BXVrgu/YqxKQ8m9IQceJwcnHXSGbE2nZZtEM1g3CYQZzfHPpQMahOE/uKcW0
7OVFDYcnUg9V4BTvRj3Ed/dXAryXraNwx9Fq6/FQty1p/4WcoczMsjlv1ZCKCWZt
ZlP0lvST3GXDUMNVoKzGuOkREKD4Z25230sxA0YLu0eifkeNH+8dtFVUMCicYsWx
QgMyc0eRxCM4bGNtTRoX6QRjDcaAV4IzYXQ1p+93gLOieP1crJLnb/W0c/EiPvpg
ABBFHxU9RQUI1C8DNfidArSmZENRMiNiRZ3+OQDFDh3TD8i23G0thy0FhhIYv0J7
yBy6mLs8ESWBWpjCCmrm6utbBFUlwwVqjzIEd5cQTHyhgTJyo8hDZP/IYBbFvl8T
klWSNh4qeO9TD9KMfB2rXkk6gz1H208VlEBb0wtouqqz1HvbGeCtseMJAYs1FJp5
c3/vz3cH8kkHVE9ZK4ouPv79rdkzDlMUv06CsrQ3ustwCU/boV2Ap1TCVp081mCn
5U1OjXc5+87hI1c/0kYqF7BD128JJiV10l/Me1vNc9ZA17uYs66qqoLO2Jcc6ijm
S6C4TctE/x1mzZGgNSDinAkm+k08vLNL4IthE4XDEFbVbTbtBwBSoO01vjYPk0eQ
VC5GKtxpm3S43rAXJ5OKPlpO8pYPAuZReAimOSZ70D8j7Cb63K6QLag1h75ZnNc0
xVJoecAKyC/SiKhBB939H2SDIB43eVYr2suFYc1dXH9mP7+4IBEs5Hc/ov9ADoaK
LM/haggITndQvZpELVVQqVw+5S3PZzmHNy2O5VvGogcVfD8oIVyeuZTZa8Mru+oY
j2h2KptKwQcz508TtisOQBlQhNes/V+ed9Gmi4BfhEsi1luSJL5X58Ak1I07WlMZ
9Gvek/u1ljjZw2M0KWW08AImUqyrbUtXl+HTFgp0XU/hEOixsCdeipHqJXdFtQgT
qOYRnMCbuZHtX0Dv+gSNBmW6xSDg22H1D4NXDtJaJJYMyS3j65u09I+OJmLIEHTG
7V8saURzQrnuTmXOdQ8b+C0rL637JmEwyi0sbcdQ+t92b8vFmMFEY61RGLBxxLEV
Uz+YgGDgOUskZv+oN6BEjE2vTKJ+HxJW85daWuKZ+uL9ylgusOvkcCGOYBLW+oVh
F+2CC19I9jzTtQ6J8fropvHwPh8iRW4zRtNbFxyzLSmt0p/C+kRhPgZRUhyUYmZ9
RATue6y/cZzCvGOCKgA3zLCUBzvXh7O7fI+mFem8AHNQXnduSeAdRKJ+d4JWwkLt
R6ism173fa60sRXGlEhbusVwAcWMW7mEwJg479JlI4p+U0EWmLpv+jnuJLr4lnxX
TC0qNEsHgMiW8bWySTiTliKkNlU4DVP54utl5Ddm3OJXjCJR+xcK8wIGJfCx1y25
zEQF/WSylm+mOhFSDpCl2+ApZ0T7VgD9NFb2gC3o9az2vDOy2fAza2phFo4eIz8g
EjmZu6lqB3gYEpHlZo1L92/lEaVnJP2VVoRbz5iAY/EEOqDpuqcpRNtrd67DVWlV
rTFPfeK5IaWxYULF6xk7FGPv4JjfuTISebWfZnMh/+6nqR2sMPFGkyXpaIlNiu0j
rgW5kx0scbg7QwsqqAVfGRrED0cDsTL//ejLwkeacLCqki9CM7C+34xa/o+PlNSM
6xUrw4IAn0RJEyowo9DkpXTZVZ/Zanvtl+ufa9GwfIbJwxWu/sSs70nZaee0NJpD
C+TODLMl1GrQM/HWDZtPuloib5NNoczbLWSmvvZM2cIIvIKz4+LPMadX3ATr/DM0
hE7BqVnzDdO6PjYEXw0VwhqCiKe3UBty4fTWn5biNo3NKZ3k86gxDNvOYVmwhC9f
veLVpUi7nLmTe5OUvSPOK7vNXkXYr/PpHsvfj7PA7IK9cD6VBbwuOFVLDS0iaC3g
sxO4UdN8NiWC+hhPfIsqo4HgOtT3vuvK68ibTo4NnRWaSuYIGP79BlCYXewOHWEa
GLR4VK5tAvxCiqrnCzAimgCs656cA+pnuQGKAwz5KHWF4u+35KNM0KUxSTz3rWcY
nD1jcBIfSZ6QI8gj62DGBSVvRUqYUiSsIkuDtvaEGhOPi7FIUMnvRDfbF0fp3jbN
zrjI3gOk7fj6/8YKEin5JgSlC03vva43QzbNHEPswBFjE3rcHBSZQZlp5cctj2Vz
JbcilAQCS7uL5HI0D8oo2MnmHMJZoFp04wX3Z4hYI7WyF13AQDq/sOGiwPY4UB2M
Z78y24Qb8IFaipvFgRD+6TNtDG/ULoTPr7nmufelxB5Ew+Ktnjx/kRCyhK4hXVDL
NAen7WEMOBAUM7MAO7QxcuNTlJLeaJec0ePSsS5EBbE7lmw0DV+eBq7IzrBOZMAE
1KpvsFollQ4B5zCssrSxGvBGP3/7dZ8jYyYcb35g5kiDhaD+msGWz81vruBR4C18
HcbZUOYWTOrjW1Y5DbfPH+b6IbVGpZgi5DiX04fJyp2eq/VSd04LG4NUwceCB2xp
tQ7G12/qTpwh7HgNpCkedhkxzp5Yzg0lkjFEOgjIeRPdZ4K/OfIOQwxMu5aW5pjs
ibtgAYOG3o/07A0Ir3PTCZoPlwHigR0sJk8Luj2UfvR7TW8JsA/RvU13Gh0B28O1
z8ShtKTTFXNVYKWlh33HuQV3DTgphi5pIg3PZU7oXFwuWeC2xiGuEYao1qbSOGaV
qEQ0HbF1GAR0NruSA8kidoj2BWsxS50n4R20JuFGkK474cSxqDB+d2+wpbQRmwHe
POv/uBOFU/Kq0fewev8G4+EKR0ZNO0GP/4c8lvkI8gVprm8kl6uMcmlIuZHJY1w8
ctMuJii9EO6EwkrxYPxr6mQvkC/eCB7xEsOy07vSC7cGNDu3lgZ+2doN5fJLYoGo
H4dvRep7Vp7lmhSjIjbg/e7zSp16RspWzHGkaAnFHNknXKXAD9CY6IFiaVXy3kJr
qdHh4Oq3wiiY0jPgXG5MGLa9jdtM2fx10gPXhMu4fv7BZIzyFA4JNLy6S60uZRtb
+CAgoYE5x5eitdh+6CoB1dKnbox5TCmVTwCYu/PCa+9TL0+VlWoU00Xv3Vvb2N5h
PjYRmIOG0yDOYpT/dAtAzc9Kp7+BoWgx+jFCV75bEQZL8apowghISttJCGbAH9WC
HKcrnpdUeGQn18htLklFgZaRGr/H+BM+r4X2JUtvwB8HNfbInghkckdsDTqC8qRK
ADTAWUDPnmnljTkAgd1j03fUBSpYv9vLG6xoPhQQtBieYJIZCPO2qeUn/YSdD6sN
z8DZOQTLJgAVqKlPvZphCrofAasMskajuM0lrQxJ0CMfVK+uVXf55gfeUyzAo4gJ
TfgxdDQgpgfgRlNXXjkhv2OVYRfXXebVgG3hsn96RQjEdiLXmjpqe+Na6K0Jbbe1
aMRZxgEXTsa57NFiqaiVV4ETQ0tEOW/h/lrp78mUpoRV96xbhJs+Ghatu/vfxyFv
3JS7oGgYjmjp+ucn/+E7VrfsPUEE/8aHvMolswX9qLnE2kgvr68xO8McJUHvS9u0
xXYF+0XneD1IzP3oTi4vAL2yOUYUkCnq7QjAwpxGFP2As3A8jO4xIDzmmuJmO+zj
KHWOv+PBb7YxjbxrKRJ3N9jrWciiwMf9puLsQUlM57XuKs/RsDb6pF6MB3xhHqF9
bSE4Smac6yNRT9/GqZrzRGKwTIG6A6ztPbD4FNUTvSCiMtvwCg1FEmO3b1A+zGmk
sR5WqCSRs/4SslAXBqpEn2E5zm9mxcV3YNk+Lv+tU8+rOgmStrkLCT6t4a3NLZHW
e9f6eJ9+VEPRU7XoC46xqLUdAjEKWslRW3ZhkVNqeV8AWSRXz85mbPyUQfwW7MeB
nMHEtdt0/ohOpNFDgSUTVZT8Eij/JgXm9shnoyAN+GbKMDwDgd5O9PMGGYUcnPiq
H3jac5NZpi9YRE99AS7DfrJpvpdwAcMBhfSs2R4sAAC7ZqYj3DLRrZrLyDI6ssC7
B7rWxU+TxpQUoVKmHsyitw2BBzkpwRJM3db7EjBzsMAjUFJxH/Oz7JVcROJK5vXG
XIgk1MWL9lj0YpYfjKHE49hy1bRNQXjN4AGieng4bVya14Swg6TnM8IL18oHuQe6
v330PSLaOV20pYsW/KxQjt1FJqSV2dvhzTVKDy99Nf0R1zGJON5Y9uCGJy5XM42O
ahCbiP7idL58oddPgBxt2WMD4J4QzWXXdbSIJOpgIBBsFsmv/bgVxJcdRpsGuwZb
28D+AqhcrVaB+8KV/tivGBklW9KMFjaDlQOTu2yXHS8a6mv0iaQ/lMFL57TsliEz
0GcQlPXvrndyx9YWIMh9A5y87NVzh7339LbvUaNUdtxzL5bbWpO5KyLmPPxVZZCL
DmxsqkgfuRJ/eUErlyrxUjkkxzXn0HVFpqEGRohFwhdKnbzezZ1NKxz2IpO0FdeY
ylJKgRrW18CMy1/pGEpHJCuIf/w2CIRzmVaBih2rYbAK1Cmib4EXBAyibNxpkZ5x
ck+P4sLDXhDWXF3zNi7n2qgcB1BskEx5oADJeu+q9Ilv2httdsRBRBP/B9jE0chZ
DDZ3nJxihIu/mqXB8OUrBXuvq1y5Bl5K1T0lza04GDIYfntoODiClcGgPURNj8QW
Zu0Nw6hxkPj4jA4gRVP3KXdPyseDzDsH7ZEd0/ePf7koCD5U58pKHf4tkGCCjS/t
1iKwRS/Sb05UkG5mxJxu9mMRSWJWJs+E3G8IdZlJKcVoTJqdTRozaPooBvcVAbjY
JHzFnRm7SVm4EL8QHaxLGwriUIv78ZjYV1MmseH3wP+PVD6PpJSqFqdGocCE1gur
imTfewoiRaRGjy+cyvVUO0fUnEz0ad1fC6F6xYDqIgAZ59yBrlrW50Jprl+rBZ1/
6LzmPIgK31em66oD6aYisB/d8zURbMdyV0ECLW6RI8MRQFx1WuvYfXgn5tlO2ugz
e0sPmjk/6RCyb9Bfb4bDHFfb4Vk9FXNSf6GjyntnVCOg1FuESb6hzmf744ua9JDt
99fziSp3LjGIsBhSPP6+7m0Am8piVBm+H1KuDrjlsZ5ZWjQbQ0ZUFHdWgq2+8YMR
FhqpqQqB5s/oc2xsuqiMZBfj42NPM0UQfY4XpH77zObzzXKoeA8rilGF46qqSBVy
vFxKuzbsOzn9V5M4aKVMRD1WIuZzsNbP6aebnHzoaXA9jgM3dkcgNjGeAKhBY7G1
LYM1th46F4BJYzGVi+g7K1eMTaGdeTIemJn7+OdP0LGoaVqydtEnjnIQ+xhLCtWC
MKzJHP97WgBy8l4WrjKykgNVNX4CKqxUl91n4rDcmWLDeQtYRQFGbljsNqw+IAkP
u/hom3KfPIfe7ViCc6GSLTvVkYbN3876LHDvDsTgcZ665zAQ+Rx2reEpKO/KGojv
wgRhkRqHw4zjIIB9g7y28CjTMrIPPcoMh6qNu6sTI9PJrMNvCThalCr2PW84XrDr
Y2Z/A2GG43BNxivO4Kq97CzcXzoHSK/CNYCDSby37Apb5pFhxnCp1drZmaHzgYOz
Qvvs0Hm21wRo9yps3bk1NnU/ihu1eMrImv8r4rbxnmfMxdUVmyjfSmnmDe+l+USP
DdO0qUKRJFfSvCLP/SW2+B4foLQ1ckjZgojIX5fTBXGa6YOAC5h20wFbQaqWBc7N
3ecMJiczLx1tL9CruEciz7jRYw6KI14pfjs612O46GaoyFIz4F8Wr1IsUSYay4ck
/vxAfOofaf3dLxQ0YZOaktK77RU7hO94U4pI+IzUvSvSIYAK4qP2z0BrLq5W2MSy
BVdQIp1vxd1QcskWudULPDCF/TGQ28p9qJm7PS4Q0Zfydo1E2fA+X4Gn+z3rxRbD
XDlQaR4j+OTiGjfdcEnt+92J6GV2l4CRemju5KeWxskBMW5+AIhVYP1BCPrsanLL
klE8Rd0OZ/KT3E6h+WjQH+cUPDSlDYraIGwdhX04Huuy+IsgEuuhiPHFbUgbuE9z
k4DBYhB+38OyhZywYvjtrXwC1Z+D1fC48QpdE8Q7dwGVp4cfXijslvrTe2kfBLYa
Bi7HPwiuiy5f0t6RR/BgkuUHVxC/flJNr2khKay5BI+Zbu4StZBD8FhDTP28jNBK
+Ja8uV0dbPh5doDEHd4adiNhNidaKlBKbW3b1IgNisVSACTXE65kjzIlaQxWI1Oa
6zKULQ0pMFb1nkZHHiZlQrBSvdcuG4Ll+UOeM9IE25yt8rHe4QLRf0GM/U0K2oEu
QCZmrBiHu0Gg6mcCRmx5RIESyHEUHEHYIddeUTN4mpsHUqIxgcg70OUnpqTPwbsb
PMU3H0IT/LVc4AK7jjyJLe3TMtsi5X7spHNeHBbtzsOjM9jtfw9Gx0IksO1ZtbGI
O28qIEUKn/w6iSPj8OC/Psl1B63MkY0UmFPmZAioTIQGNXwy2Or/TctBVblAvsaO
Iyjq8iHQynZwRMsM4ccB2WF5PRKExqP4HDpeDtd4pQx50/FCljjmTzGaXQBt9U0S
26t7J0o9WH+17aNT4HEVsU6ZuUgJUgmIRSwLZamfrskZDr+fbP7BTTOkXyLYVEaS
fY0RYC+Mh0W4bfrBS0DKQpwZ9VYTscYpOIIbdQ0hoiVmK9mxdO35Spih9kp/loOA
ns8wCbEOkh09Ol3tqynUCB9OqbUFnsazsvNkOI7kBzjftb89wlIXfaIJ/UkdQ/Mk
AhYx7PGosj/U721WTF6VsHgiuuNnkHhOVHvppAP0Ze/DWtraxZYtF2IiTSyjnPn7
a9ch5YNx9i+QsZGbbG79jMCY+hDYo/KisqqZx2Aar+fkwHZYnpEKjZB4ruZsA7Qa
W73NDUI8vvXBgZQuZfTZYyP34CGDJLWogD1CleTjJrHdWHNQ8YxN8Tzvm0gHRieT
kMhSp+TMweV1MyyUT/UU+hCy934i3MwMtVNieNSO3bG6ogSc2STpWCeqnYJYOgt6
sgERG2Y0pfn7sGdPT4AIKAVyncEAvEXKPkF2tofOOwGkH2RRp0ngfju02Pwt4F6M
z+5JoAlLTGBElqTjr3E8IgvIsS4k7DSZF2JJz1JZxx1F/HzmzOeISMRBeRpWu/zT
3daUz0Sv19Hd1dk9oqksaq2xbxBJJy/axCZSiEphINCCWCB4XKfcUSrBu28X1w+g
IX1WiB/Gr0O2KHe9xX3TtQAOTBi4OZc6uIZ5/OiuZy3xAd3k7wE5m0OeTfQ8sakD
aNGboNYoMLXvnYHRMzJMZNy1pEojirF6tMOgXmizJEa5WHrBfjSuHO/Sxduv10iv
uJWZ0Oszyyws+Zn00VNn6P+seqnrqUoR/CTDg8lVlagIEh6l/tdOkH3ke8kPl50j
0aTlSt4geXyvqdRwwIZcyuaCyCtje9dl+SroLo21OltsvdMYycqX7FVH1o8tCCcw
4MP4yg6BFy2lvybyHZKhOEhofCHXWoOdcT8R52c0OEMl3ghEDVuXY0NsEDyrFM5q
RkGJKs9KsxdXzQVDP7xXLcoEZeZ4takRsLFywN/iOXXDcX01kuwp/1ZTaHsgkzz8
LNxRrW9BFtuMrX641fFN5WKXLl9rdwL2FFKQ0l2uphD2XBYxRVmEGo/CqBsdDZod
3TDfTzDaVhThKzmppJsN8wF76s0hE5N9d3N+eHrHn2FZ+Lgw1GZ/S0lJGSNrdsuE
TD2RPe54627n3jrDbjO1j7tynGEg+9w2oFTXkm8jpoZx0EaPOtFxtWVbfhOMnEOd
3RXH7mgkWFoQ6NEfHUbe6sYvKiiCtYCJbVQ91l7egWF6dBgUcct3axgCtMSNigFV
s5JPwhTlmLR3Vpsjt3H9SnqPOifNJNRH4bsYLUuK70lBEgCMCKYoj09vF+NqYP6Q
tmT4pVZ9PGtvIwyHN+Zy+8ci4EbcyFF7l8ljPAFxskMdDvqDbSpq824Pf+rNEOiC
bjmytm7IPSHk3zdGZJMGFUvsyqYI+hc2B2o3KvTiqzL1RzGkNU5yAFuBL8xC2rnu
yQ9nxqVpOGJsPcJdbmM5fx2FI77erXOzU1hm9jME3AbcNaODxb+9LGfm37DR3oaC
JgPPBxJUZCexFC8iJGEfb1nJmwq0095oZ8RYjf5XmExhKasmCUDKE5lLJKsHPh0N
OF3if23WYd/mhny8Eh6TtIFBnYhMRSRMhA+TVnMGbVqIvRd6BFULFMZkWIuVk5VR
sEiSm8BNva1WO0Lj7Pa6zTPXAlvOU1ADfv9AL10no1oTWyvpcrp5A2M2TScOcYhK
SHicxXPaDpi28Y08SuDJCgDyNUYMVGx7RpIPWtajW8gorP1AfssilVL/FISFj7sO
cD4jRk3W42UDeY9ExKFTzqmKrwCnAfLLu0OjYbitryHgNIaM47HVsy11KFGREFfH
hSNRJi5Z6sDgze2DAEjYBxdiV13BNbSVLqd23QnoMFdXYg7+Tqv1XuRr2ZsGN9dQ
8K5P2H1fea6DPSEwzvYkHDmYRAb7ADkmc/0D800r9vWgFLMYnabfT3FU3WL29xL4
py/PsC6fyeG3YMHjvXz0CKUu2TNgeUFn3sUPuLFyYskKz6AnbA70PYSMjgivpB3h
5nxajchD/D5yx2smyo3pU7YAkRvRlgKbnClZsXv4PvKSxbUTEkCvOXjkqi3QjICM
19EFzuy7KX87pAfAW41NMTIy6aJzmilHNfKQvuVNyMJuhvRs8tfND+h/3OAOXR9X
7tP+JMBPgX+5EEQz/PtP/c/307PfnnmvDQcTrXD14hfY4VIVuScYtK6H2TNtzPoo
OucrBztPuKi+uRqfDDxRzqr7XrRUvEmWoshaMOPSsPru+0OitYCzse1hq/QM/jtb
tSl/N//i8OWazmmsNVkzlpOaBR7R0pOctec/HwC9ZR8WPHj3SKLTYin/uh1Z6v9Z
u+QIVg/FYimJjFTX1hV+T5Om2nMv/L/m9IZWBu5vS9IZrHAft2P9BYsCgYOSycgF
07GzIEK9VRY7JUdmk0pCu1Fg1E9KajnvK/H+5mGE0+F5jnZ/tZFEpCayBRPv+6iA
lyR+txVBukjvNo6GKtNHk80pgxWpgpo4A/2A1P30RTsjvA5fDdBupmx3SijeHRbR
79WyMyddocP469PIDVKqzuKUsj4nXlUJQy9F57kAAM5ux6F5sz7/44BBLwT7NRhy
PPjM3+3vm+Co+0buOj5p+YA24BBkau1rpIGUurFJQdrZinXKKwXJ0vnh74P+YyBd
YAR5RJZXViTF9Gz4rYP9vCxZtdGIzp+bTSKjjRUJjRsSmUXOl2nz8s9JtPol5tpp
gwn+SXLli9uerygvrIiGfIRV4RKKU3PLqaX4tCuYY1XMp627LVS9ABwYB+gtLa3s
IZL3tdY7mlTWPUevlFInPM/JQMmvIs2CMY9XBv6d19t8uVUFZYM5dlrH69fE76H3
l1zfWLvieFOk7UhVdkZ/bpiSG7FcxmjSs4ivwYi1AFR3pAgMWE7bnxeSyRowc8ys
Gtz6p8h6UjVnz8ycxeTR745yF0miahQIC6ZHsAmqKo4sKDGpoXpck8IpTmaV83QA
N0T635IhCvmM4cZ9bog6yb+15FpcUVOa7pkJJpDlHNofK1yWE5rwG7yR5sm8Y+6R
RKs3mADIysS4J2pnz0ds+5+Mt7HSm0HNS5HGROOUXxdwW7ARuuXtWjBcgP/vmVd5
Dztsm6VE4vG/gvN2hBnsuzef9k2Bm4+0yHKptrqS+1c+ByTmIPOeGrwj9DZ9fvOZ
`protect end_protected