`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
xGdV/Ahjc8BxJpNj9LtOOux/yuUFtqHwE/8PuD85sZ/laBXcS2EyRFN/0U9LYZVa
3I7lhlcRyWvrZ6E5ChYwqq/h1YR1GDVeAJGYvlQ68t7aFEP3jIEsUXVbwKMKfyMU
z/S45mW9rhKqtoOizDNFgW3hHWHuLzK7lFGo3c6GyDoiA4x3DM6QtEKjVcn0WRip
R3N68tl7uJ/8A9WOW2RwVE6XVCml35DfMlIeH44xxJ5JByVfxiAC7hmfST2MYIPV
5sSaTTosjdvv3HQz7VHNnWpsyKPZ2mQMFng6j4/U9dKQ4XYtnaBjiwQbUrzzXGbG
8V0JOCr6t18DmBR9+hwrghxa5tgn5mU9VUfYXqlSRLRonHJnvD4BhiuQQ6ckCurQ
uzZDN7NtUkHSOhp/mNdb74ZKXsrVx8l52C8x0ziVs3aMlQAy3N1ZsJpA0pZO7CQG
wCDUybzKhg5l/JDX7o7K0wj/+S2rOw0c0Mn7X4R1qa8eGpCmjkKTonmS9tnj+oL1
njCNsaYBywFhR210RLdZf/8UrGoEGhtoBN4NI54kWHZqZaCOhwbM8G4lWnOzUDxS
BrJkm0aefKwGG/YTUXSnHSLZHluBc+xbcMhgJEgDnjeL8ICoVCD1TTIkPjq2+6af
z4OiKNnYJmQeHlkTzZPT/RE3L8f6s7fsQlLwroCCdSEu5ZqW4qdx3Elqbc7gHfDN
l0pIuJFJum75yPWgqt2OkpMC+LgIPyuKDYOQrkOPtg4qGl9fCCAIWlQTLWMXq0cD
EE0duSihmwuaFrBSs7pGh/EtAdJdXiSdmGHHTFoCeYjl9bMG1ZZfJ5jNxdWki0Aq
TH4IfRto+rOl/yipN3vbg5Rl+DaxnJvVKHvmfZEAdhy6m1GYgTwXT6/lSl/gSIhW
FyRq8hWyEMt9kAGZqWy34f9oC9KchaSMnolbu3FW5cZJ0cusFdhVNClg/pPFTm38
W5dG9ZWlnqr8RNBfomb1P4hNIs+2MZOoy7RdOMVtxcFJyB93BM60pXYe7meitieQ
2DPUiWFT+b04vzLbJR/EVySQCANwJ7/ZmOcbrfr5EJ/Cb98gMY50+Iea7D4NMk6D
LLDexxR3Z3soZaYk6kS/jt9HuUvPpMQW7MCG3ryezGOPkTIp2jaFdowE27xPvkws
YheQcI4ov7rgpKjICmmJU/N2o1NGQw2GzxLMT8bjp70kxwtlHSXo6LuxgC6fBMpL
BXSBYZN9UR4vtg82YBgh4MMEDHIcSflvFAZbYNG093mdZK2B5NCRdZJ8HncUhpxi
6TecZfG7APDUzUC4e3JIQ/aptVzhc7oatF/ZyoVQW1eqYNp+bDPMzwrWRLC2el+J
dZOB+cmjsLObDeT/+cT0TPxxwPd6QTMeWuA99ERVQwcLV6LS3O+rxJAnhyJj09HF
cg5L7QhSVqSpxuwbxAcjEBZNU0mp44UPlxLHqHmhY7hN9ripbL+7ntbLgpxyG3x8
fvL/de7Rc2yCSzFcWiY9QoIw9J9iv3gH5HfSVb18Z49oI3DgvjZbQ8NESIz8IC1n
KCDisPDqRfT+s/HThRgjAnRB4akgN0VsU9LHqR4iM1CBB+hNmQ/dweL8QPPfrEf+
yeaPPKD4G+BdT5z2WADEFXVJuT+Ljm8OPPJniRNuCVGqkk2LrUFi1cD0uPx2Iqyr
GPKurmm2RSoJAtb6vAq9hbhpL/hKDvOgDkbTIWMSzUTZmaCJnqUWuMq9yrMJzpXn
bU7j3ZcBufVKN2XHO7+uthoQNDoRSsk2zExkP2akF0ONl9GMT1a04LPRJeX+jfA2
7+a0fJ6dxRf9hKBIZ27NGSZ3VCE+RcSX+RuH0vMpz/OerTnxeRdtuzeSsaYCl6xx
5VpDZMAXEr2VxpTiTPdJZmB3BhM3Xq444waCkmmBMVXkBtJnYxuMG+jnDX+kgO7a
ihzmDMH1+6vpvRRkiaaR/iiooa1I9VqMx61czxPehWuNvJ+luUNTi2+2D+mvBTcA
0Pdcoyv8HmmWUSjIni15jj1KGSUJpaT4YbKhSRa+Ew+zn5muEZ8KHKd56YQRQktc
Tof0rS4WlHgbY7ramE2tjMQfrEdhzR3bmLGz4H1apDgf+W/INTDFSR0SIdAPOvAV
Fb8SdY+C/wSGIpGbXBGXPhqiXzKPG9DBB+BkJ6Jk6Be3tEMBxQo6jZkJVeKqNt8O
jZWjQQXShAGXsgywCimXE2mm+1IJFXTSrOc+WA7tx8GZVFETyTybDrGYTpmBxpO4
G4ulWM9cPwMNrd6HEQ3Lv5TKUWF+zn0okMfWlvUr0fv3QpfxJQS7ybabM5T6jEOe
4FdfNYhFU3dYVyvso+v59EG1iE/CwxXgwno9Tw8MjZ70q0YgOr2hWZNcMgfu1cdV
HbnmEGXlwwTiH1L0AYwFxZBBWwLN1dUR0wdkTyWWWzulSDy5p/OggCGNcOBapwPE
q2IXTQwDap06rdfJZfL3YQOVE42AWYCKaLc4k5KCyVN3OM6uApqc0Rc0viF4UhIU
Z1Ds5uBwP8UZuZgIhWXRx6M6gSX+bRFAdj5oyq59oGE45UbzVc/+bdmMtuzRRIiY
YrpYOxEdVm6PM8MKVB8FW2NKBFHCcLVaF+C8U0KXqLRKWRnBz19QOwV7pbN6GYuk
qAYz3/N+Vv1tcjI+7eDj5qR1cMq+3YJ4MEMTn2j6hKp9j4drN8msoVfEdZ7a3ltG
D1mVyC0F1GElENEpwVl/brhh2R7CGY4CETguPH8rOu9x/QwRVwu3pPmlutV/Sz8v
Xtgn45HhlyMjKgJqSkzkx4hvb4NX+QNDfl2FXN0U3KGOEThlM9evgtXEuKHJ4Aqp
XuodL/f32rpJkDkc9DtRJl0yPbveGBdBSMADxkq2HfMCeF81CTFlKo7MUZ/c24ge
EODBSflhwyCMNoHqwUhuNZ/drKD4GJJHoPDSujBb47KU940q4Pf4bst/fMvHmst7
ms4u9PY1vCOojJEfVXaDlYLixIIq14Vha4oES0CZiBTSVEBBHmKB4Pbx6sAaETbE
ZRhPGniSi6bxsNT1271XxsTc2dMN7JJXDuEPFDvJ+h/0jJJ6OcO5gEVh+0bFNUY7
tEi+EvkaxqTHOqbU5IArpajlgDbUYg8Pue4SEWPlnbHPNiyziZ+9R3lpdan2j5D3
wT9EpeeGaqWRKPMM17SzabzkYe64hj6ujuBnl2k7k8ypB7rGVGI3N7XoRi4FWCpK
escCgZMXQ+OLboUnvEqyTY9LR2Ejaq7xKQXfe1E/6bzI3oNF/JnaCWERKVBJcpm8
jCY3mG/NVevwH65hIzmsYHLiEcyjL2dLTK5ceXy9cQRbaCgNRtzUSCFw9TeHJOzM
d7FyT2sUtvzaOSVNN32vCLk7I6mUOrFKYpKvMpmdkeA2roSv4uEdJtNC5ibLKlbo
lGW8RHS+nJXg0bo93L3lFNRIDr+YRoNm7goUCXLNc3V9ouAsvDSvUr+qJN0b3c7D
Qdr/VkA/2jiwhzhWG2qH9iDKo5mC8MHYtV9zjUMNIw+ix73smNWVSZP4aOBIrr9S
KIoTCnwKd5TVbijYwbrkYl59Kwq/NSsRSOruSXYnccpBowSmybRTDQu8TghuNAM8
/CzTfKW5bj8bhuXbHB9oYWGH3XWgQMIZSlDKmg0tRJnDVn38Ydl37m6hkzQvDSqo
N1iS0uNcSfdo0za1bUjlkRsPssOMB3vn7ZtA1tGr2k2VP5P1vfPPtRlcaRKifddq
IpUkLyic+1DbswrHsYiMgT+tI7Pf0xufBeoJbU92UxVKBCPVBkQ4Dg5o+jlaRQYx
NJAKcqD1cnjKEW0b9k8UuCoCuoFutdjsMj2w1H4zp9sCXpwTmDPanWBvUBbOgojn
tpq71aiTLmoLdEJd1SXcRr93exictMhzrwkWPe/XyY19f53+BxbRx40N/y5J/aTB
XpbQkDiBCFS/8sCcWEmzIJNbt/fUROZvN4d2kbl1zu1C3/TR3qsuguBSEEkMXUCl
d+kiaHzxJX855VDjvNyYQsUdGoUjfoUJkNVCQmk24zK3n6ijLG0FCcVIGXFUb3Ie
fDTgEl0zC/EiI99drcVqk5X8tPTgpTLoZjaIAu3yAckeM2k3wqQKwRd/lmgtC496
3qyJ3bOvj/S3EP6VRgnnziwqp9ZEPKO5MUzfjtOV+grg67IhjNXDzuxGyff9dbQA
ZVaZ68gwpqJsjUKxHO3GkB4i6wq9nN/NhKN/NTbQwG4t07dseNjeGpmozwcexxn7
fj0SrW4uiM6nvvd4b1APiAV9ki5s/U70UrRJ5iMyyubowGpyKi3P5WDuw0BkziYm
DkqxkdQwip7yzlIab7PCkNgu73Am84fG7mk3jUTL2+oEDA8Z1cdCAYorAUi8uSSa
b5xG4QNVmlYw0IEbV7YGkVzqA2/X6J9ohSwio2mILZaCQHkK1SSk2dsbWyT0V0G6
m/liKJKElBsMo9SNMszCsiWgDOR+lpqm863N3iLB6UpVtK3EgTl43iOg3Uf1nbze
VZ1yT0VMyGUUXFEgtBZqyCmPlepUY1+FPFQR2Gwccdc50t3+Sb8PZbe3Jvmu4TTd
JewNF/kNgLRvsJEFLUTBZJmRvK0qHb/Bnsk40i0e/Y7E8ClNeKn9Ne5l8Z5Syrku
TQFzgqABWJzT/rOYEZeENGU799/e2yU6I4on9u3rUDigrcfHkbArZBxZbjKJNhB/
UtrUosCXrm5juCbhifETC7IQCBLBt88HiqP+iwVvQdRDGUqRK2hMpAWF+R2vcUyw
yABWn5kaObkcMMS0Dh6NorRrH/D83xszS2leYZfV8vKl+rDQ0z/vYcAPx4S4P8vm
FznLba9cEQD8JoEk+iey7CdlAIonit/d364AGuDZMVhKBmkJxtYHww4mU/etm0wf
XcNLraZwK5l8+1KeXtOfPejufvFiYHaCjrxeOoRsVJPC0ifALUcp2ninMnSUGH7o
eUwDzNkSYPnR/Ajyge5qKkOHSLR85CVLXsTrsHTh6ycpO+7+RHb5mvkASvi/Blc3
lxovAf15zaL7iNyoXTM74aHNqnF/p6VHTXlZUpwNb01ZDC5Jjo5fxkmVvgHgZZPE
jgjbTEaHiR4vhH3cGiC+iCrudj7BcmiIm5D8qTrf2Pyo0ON3jAXj0N60nIaQjh7m
SlC4T0dSpS8HkLbZRfxujwdA9rTpoGFk2l77qE/bZve2EZOYfE75JnPEV9Eb4rwD
nVmc12pX0aQsEYBTpGak/z7m3vN1gOuS3yFinlVZj+1N9/4cMWCtAKveH+qeTr5v
Fz53WJkqTK+l4C6cefm7EgieTixXcgACkIwQohKRnhnltXzCHVI0DQnm5xr1pq+S
PiQZlZwxfuLVbdYvsqVNvsZfLjPQjD4++IMDvAfkdZni4zUwFfyuB6GEcZ1gee6H
klTR9iiaAO04VP9byHQ6VTKNiIEu5TjNXczSRt3i0VpoY2LdrWYupvLwBnPHz+BE
AdolVY0lzBZaCSnjYVajnPzI9s0q6Au23EJJPJXNqXxmamndsU0kG9jbzke2vpH8
S7ZIo8zJJzNTNAvIpmh+3nHDoc567/sKMd6WfVKvWHF3PQ0P+stKaOUJre0Vqaqb
ynXglKCCICzja4F4UYe165Vf6W64YD00fQL8bFv2vRlG6vdD07ZY54HVNblpv98d
xgDSQ2i5vE06Os2HvFknzx0uwM1Lq5VhFn6uSPPXiH6W2qejWx9YUsWvPr8CnKem
Ryk7SwIXOcyb8czo9Hi5OYJKfRHQI/JTbkbHPQcbEvas0RGHE6daMfr5JbNq0GVq
+lC44TJ0IykLdBcFOD7zqYDrYlQR3Z4lL2va1EqMcJZgWvCVRH3zeZhUpMrcuxzc
gCknIgaJoWU2+fq0/bwIfWEjO8AyDBXl2erwqXfabEWVSNXmgxsq4QHZ9O2TifP4
ToAcfn87VsKv6XrwQ5w+An3ELvTk1N1BBm7h3YYVf105mpRlbVtac2aU2VuDv4hh
guhiVll7hLFAS0IsGzaE773vRAq2SbfsDVmOzxwhwVClYMHwtSs44LSmzy37peft
9QyYYSNc4eQmXk2loGmtdn7los2d5rItJdjkgKckwl0jVF5/cUWfnrnUYAL5hQ9W
ZDrbNOY7JxgbtjW7zA1o7aNEhXJCpUHVjs57ZHsuhmiT3ZSRW1Qhi0XJ2jCXnaEt
Na6TkXvMKVWJhH/plPVytzSASI443EQx8tQozLe9cvGTyRd7A6Duj59S5ugzPttY
f0DLpZXtPhD2u0IQFGSFf32ejFGrYdfSsjgOx8Dcrgz19JwjCbtCXYBDHBguxKv2
v0Qq+ZYiuh8SM4oOmtTnnuVXhMjmEQlQiEBL/ryAdZIBGDxKgkXrs8IpBkOPBWtw
PwoIEcYYVnZAuwdVdKDjfIqikDdYjgIbJf0RCUGpYB+Dd37z4NcQFs+kNbAHDKsw
4STu2vgjo4WchvZs7yNIUTQDzmhDqPC/ZLQoOHFVEGouFF7TTMlAQtl7yKvZ2VgN
1tSlZfatM0jaOtV8gZsdc6tKDVNORqf0dwtCcRMkH5ErmEiFUTKjOZpBkUxanuGu
HtR5oANhVpU+8vUahkyMzBvQjtMKLmLKtAdPFFGeA7pWabSl7Ic05qd0kToUV97J
CR/PSxHXgCjxTPgOrHohwJ1AmaJT3e8PtIVNb5RKZn2bwkHOtXdS1uIzVwFGRACt
hZU4McVY2toQH0tYlb+zbhRz+ZnHkacH6PbnkjEyv3bWU9VDCZ+Re5k4SPefGF4Y
rw17PhxizDtMrE9BW9APkLF8ViduA+2ZaQvHjjKsQHJiFZI58BtqL7CuAY+kym2s
xHFtwgegryZazrLH22q8AeYS/fVr8eyHpqTHT+xAtRoiXc/Wyh1MA99gwWHXCFf5
bDRbAAuWCFj8Ug3TKG+AiDLu6Z669rS7JIy8RwK8qyrTwK115M0uS3JBYhlbvxk4
TQkffhFpbwBzEieFLVrTEDqby/pDrwzBn73WfLOrV50qHHmu+smXcl4/lIx2IXfY
V1f5duJbjsyzkXHkyG4LDJGqXU7KpArC5jJknsu4Rd8Hqc7lyMdhs8D1Fgsh1gRV
06OKbfd2Rx37U07baYUiPBfSS7kQ7rzQk/c1HLb0uizNj7CuFbY7b2V+Ejw3SQxu
gd/MGA9DZtoETlQbrtHREkuypMWgNWWAM159TsbSFsBewEIVh3S/UfECqCKWYk7l
kNExBw1uqpDkcwbOQ4qSYqspq8HCoMO7+QNpeVXoeCSZcWPj8FW9JCe7Lkfst7AY
zXxZ5uv/yr+cvrP9+B0c2hUYY/u7syYk+42t3j20BBREObcCBLeNdfSTAWKEB1s3
zF7eaMWktaW1p/X56IWwvhab+ElycQ5MgI6ISLZyQjPBpdlhHqWua/0tRb/6KAC5
CWpck3tqFULIVsTUMakY/4dT0j1+YflT08KbMoTtCsWkL+Rjgwz5+IytmkFzqIGc
KhrdVAYPCjpdQLiWT19okdyDNFkotHolvkt2iR4L5PyP+LZkJI9Jno3OI4wYs+rI
OLCmQX2va8Wx1HfbhmDOtPAZRAbiubdf7grrkxU5xaNQbgarmI4DOFNkcpqUUp0N
Hz9MmkqTUrYrjCBGzjyGebdqMpDcQ5Tieblj9vSRL7SLlEbNcYTlSkR5ip2vgt6V
O2cm03WghRMA9EUEXrkWKet5j0mVG55D7/Ch8Yc2rIgBZhh4DGsBZjFXeYejg9Xm
6bvRVpmzGA7TKw09ADrGdTbCdESOOwG9h6suGxeS/c5gy74rxBuRcUdjfWatFyJB
Uo+IM1kcONVsJlufZ+FyY1VCicpYeuiGKfIYqlbA1oYpSN5GDJ16mom25qUH57MY
Dm1EWBi6A1Zs1QVwLrThgKJsacwhAygMetSHNn7bpQfZskM1+fcOrDf1UOp9GnMJ
V8WgpUNrR2s252qqR5v+rUUuzSoC7KhovH6iSzLd7BB36D+DDbQc0vA5+BYOVXFe
/9+AYxhBPkchsAEodeaVOJzitPgXWWyjgvDvwMliiXYIH4jli8E55wtaSwPLKjap
8jhaLEMi8MAAMYkJsGtySI2TgUF5eXfkv2wLo+VMNDFQuDcgSxlCUQ84PFE0zcNO
txpkJoip/2TRJjuPJbO+CBp8qZkQ+D1EHKTJeFjgPt5EfJgwUBu6S0grxySFLv7x
fc0cn9ey+UGusKOAVj8NW4EgARoIBuR4jjqeq+eMQRj9wQK4fPtnc99hWFKNM+t7
edIyuS0WUuFYAAK6PXe7a6JaKhfARGkdfApDZJLgdHSdO/hvf3uwKlrYnlY1CN9p
7+GAa6d8KmWfZkhyYiFd0eT/3cM93QjubVJ5S7k299sEob0IdHxr3+LgAWBh7Q6Y
hXxXuirHgwqKPQVjASMnez0+XQpYJ/P6y7KO6cPdJsDf7BUjD6bywIpyj8Unrbd6
9o1oB+vdE4W1IJWemEKtBUcvYoGIex7aVYsk2XBOUvv4CjXIId5r9BBDIQZ1crge
D07aggyviwfdkvt/XRXxa5HyJ+2mUPpKO47A+bAXzQMYK7lQVm26b9x6ymVBBg8x
Kf/+fLzSwOwz01ZHcy31t1mtJx6KzBFPCMmG9WGVYYqjltLjAqvxk14YyMKMj0/N
VmJgW+rkTZiopHV91Ur5J9UMimD7SdanTYeV5Ej1gUankmAE1cmHuZWikUfFNl+l
8tpX6pmBTfcQN3qeCJ2Hr1EHaR0uUXOIzJrBokAPZaU5Ptb8oQ82hT9CdYB8ffJo
THqfid88e9ln+CQxd4P8GdGcUf/9n0+ZLkVi/nSEmov2JEJ9ilrXW8FFGsYP9ZIk
EL/6BEe3LuNDKXHXlgumCfMu63ncTQYaWZriYCNND0Xr4LJnYOucyM1zgc3wNX0N
cOHJ3JTV5pQ1cJV3IhNbZG950eZMj/SuHvDWh7jB2vAQcMd6fxhhhErIa68UBIKd
JvcevxZH3mAF3PmKWJ1Ch2qit5Uf/2dl+H6w09YvKDQUjjxCXYLfQzZwmQL99Dms
VtjXG0sj8omaajZ/zVWZwRKlqK56aaoCZ7ktwWzCr4jhT5SPodVtKjgu2ECVMrWr
9pTXtFyVvMPlrGaXD7GqDqLLl3w01xeyzr3nIrIFtcZN2OMaj2abpaXfVGCEc4Ql
2JapJxrHcfP+woFRJeOCIFkoINVK/dUwMH88Y6ukmIPs0Xx1Kxtm0tCtWst7sKtA
CR0Xf1WCbLehtEeAZnUrP6rcwdI9+cCD2nRAlBCrmBi3x2eNLKsqHFkchRP8qr2V
d9xWFia1bU0UJGiXGU20KSmfdEJafKbJI2tcu28OpCsgAM9QZQ7guxe13wi1XQ4l
7Q7iETYWFZYJWrcypGgiJtmK/bLG+mf7Dxq2gZv/7KRW9anq0Z+NTT+mlJnWetK6
TUXdv7rzjwXSyTOHGIoXe2zr6c2KwHvYxpvPr1dxlt8hOZ3mVnyumza/m+1fnbKs
Stsc9FAY++oezQbcMZ0A+0IDqglzQq5mUXYTQVR7w/DCCXnOu16rPbqhOhEHbz/J
K+g2qhpv2xUsSN7vHxYBM/TXvgl5BRzRooEfEluHDTrOGHkqdiT8Ur6SCT0Ng0uZ
YxDpt+VhvJ3ICYBKm7t0pQeNRAYPxvtLoB5TJktBa5Sy8TDZq5Axy7PWHGHCP9IL
bbN3I9LqHdWc346Pi2tfjbTgpYok7oTE3baBEce+1/Z1oQucs0HnlQdMVC3KXcbZ
/CMk0VzLg4i5gfsdSoBTSMNux6qAgBrHFFpxc0gnGv5GVyXnzodMjnGFAohGFEKZ
tEkXLct/xWC668YsTvfCUmdhvlnAK0sHg5PjxuDlPgSxPTdMz/sGuAP3G9X0Fkfi
bP9goHoppL6IWD4wk1c13GypCYxN64atWbtEj1gPh6pY7+0xEaTujeEezN7Du6nd
H3ybgWVViRXHXFZ9maGu4aEFyMgxG+MwLOXhidbAVE870J3iDTUW1PfR6i5cIf2O
UKhRJOXAzLYL9iICdd9SrRciHKDcmnYesXxqJnj7mL+AGYeOGvqeARtn3lfgAeZy
W8i7OdGOsEaiGpfDah7l/OPqbvep39zjLfRiCe0Id00YzoMDbMQ/JgMv5+um0kdq
sq0OK1iE9Pw3F35oUjoJv90NrHUjt1VhMG1SXXyk+3kHWwzWD9j9YVVoszQnsuKr
jCsnDU2vy0RpDgj1tFyldykTkFibP9kRQZx2Jx2XQ+7tlT3ww81YGQyQaHQV1ZRd
n2IkmPeWqPqteQkel8HrYT+0caaNzu4tON1XYpdLGjYCWHPIXeQ+yruhz0R+vAKw
1x/RY+GiBV6FnCA5/6qwQ9LtTGiXYJ/eHsfl8tS8gFoHCaV49HczCCa5eaTjSkKF
jixRavZYBROGqb04Ks2VZW23Aq4N7tJOxYdW3LwJKT/3vIDHDw6eXi0ZyeLF5OXT
vdgoQbcbwHhCART+QweSoAK72Tc13wcD/g5U7o658aK5E3MjxA6u1XIUJBLJHOKP
UkkoQh93ADSd5Qs+c+lBv5l5WShkBqR42YlCsbq7XPRQTRVZNhIx+1axtlkWIcKt
HOL01rkjRrQfSyKFzWmTsIqFsUqLRDvHUDb6t2cy6VQxOrZT/91VTzMwJkS8jxsx
eNKxOsHPFCEOBDXqoT9gay27fyetGG5aYR1LoKTAsualAZ6yFnclXnREkUQcsBh1
nV2DtkzTM2uQHSMLw4fWwuIrL6AfKuGPHqRzfLSyLfGeYZkR4jAaDILPHd1k3cwB
LIOUWj94V5sqLWUauMsM+sc6UoyA577dFC742OVMg3iyQ3MwKgzwYzcXZgSijK8M
VjjwEJ9t3fwET0mwluZhAz/Mhv5Xx2j45htC0sWJuJsvKEWHljyyqzIdTWyPJ372
R4kk4XbLosvG7He4/iBirUeJCwbUc+3GrsmpnS+mu/2sI7tUHp7UBDXWuAcLJ7dj
wHKcmdD714GQ9TeQo+jvCeC+NZJsbhgg4N8xqvfvV8szHKTojeRi24yOaQkPPQKy
QNH4SaFms/Epwptuo9s4yvAu8Z29s3oFqzDI4NB2caddceQKyUvRDMSS1oxU2fuE
ksADqrSgH3LqXskhkag946jYqMqz+H595V19i2k6AD9Rof3QCnYZ+Zi9y8R65M0c
Y6BXtiAzkr7vDMsXb2APGMWg3rT5RZU4zXhJ+xSLAfT26rD5oZXhkvh76PqEb4GN
tXriZkUy5407GgKjZDrNOfT/7HP4O3Q44lOJ1wEg8H5mA/2T4f//x39nZAy1K7Y+
ih21sn2nod7yGaVdAUZ0lVTbD82wYzn6x3cGvoPkxPbS+NHypQ+6zUPCeOvpEIit
6AEqqrB9oUV89UzhE/t8hpdcbfZNPAT1h5m8jQLr99iIKydiXPlefWnhm+9QdCOp
FIBwcf4TEBwJZvkVg4aLzIG4B+CNdMtmwan947IT/3VonbcQS+Ad7Wt2mVwnf5N0
pmhaQZr/zBZPmApb+Gt57gDJrwU7tFMridE/6j4kgFKuqvwioqFCVzzTbkGzkjdU
oH+7jfOrwwemvjxcyEbd6P1WoeWlUOafH3mRwvExPtRfltAsv7/Q4YvAzrEG5QME
FX58qDEaAM3goOo3qOAIpdd1kNtj97ShezohxgHCyui+vdNxyazyRYSlyf4tmspl
jhnTgtdBUYH0Se8MI4/OksfIf4TAzeya6AT3gr2bn+JKv+2MtPJqLalZr1P6tU2U
mDQHkE19YproZfRhuQ6D+DQt7vkdgbWLVoFdMjbuZe+eKIY521Hrd/tZ2UpolaV+
8VS1TvYVC6BPHTp3w5iRs393lpJXtlaf6KMNFZcvs3vC8qgZFtGRpR999rZma6pG
UuTF1zAJb0FisepcfA05RUVlP2mFoeaKdEf189/TVq+xAxxxl9CGMKMlkrF93Rqz
6gjL9UnTP8yO0cXMRKqNZfvTykIPAIZkfOnoeCCmU3371SUCHs9DmfX0wjPfDB7+
wgde7fRSLTNLcwFTJt1uXAxtCF9tYCpmX+ffk8hm/3FbQlAkWw0sUpjTUGzLJWEL
S5ZezfErLA4ilNAmehXpTL95nz8/RNdwRlvU5dGPtQSsRjLneX/RVtZaahm+wTNv
uxnW8p+V8LpUCiTHdcvgY9CY2RFtfat0U+6GcHBksYdnLHt7S+0yzTiCypZibd+o
ZYs3pUqvBqqx0GSQp8vIttWTFo8iDCte2XfRFo8sj/944MBQaKdGwHAuQaHVS328
qrmduUwr1/EglbfSBobzOhvohkFeRbwPqWqMejiSywtZcAPICdQ5HIcj7qJz5Nmy
EYGMk2P/9r/6/TkoUVPyrx0eoOBRuOFRGnI2eEz4ayU6qqJB5PPjFnBJA4Q/d6OR
lsHxCuNcj4RQdLfGwNfbYJW14nYhtzr4ijBiNT+E4YuMujhmGsOQilWoXBidjJqW
0Zj6J1VjHgichsMOuKxfLJXoJph8y/zbkd1+Psl56FVCPIDEU7DgWs4EpKC7/rWZ
96s5u5JZACb4jwfi0zBLWcYRWtX6Zw+Wwbtr9w68N5LyBWzgCV9aQ3Dl27YCzX6u
Vpy041nCl0QE8hXUi7jLovjz0aVmB93gxjgrmqGunUuU8Q3WqSjzu2V2jZCfHVDW
pcU2kT0PTdxUEgY+/lpLDJ5Ehu9FpRtArRheqZrZWW/fLe66OM8D/yBYrpXyKji1
Fj1WxvBQwHJxKMn3qyD0Vv3m5+CFNggK0vCEJDggBVai8rB6TH8/ng8sEQcsBO9z
NYtR0UZpX2EUR8/Lk8bmPVWORAKwyig6sPChBM6roB/Arh9eS664Es2ri8WLhP70
AeMd+ViyDx8L/PdCm4sKEzdhPoVAv1TvsXEhskzsqIMZ1oEvdDa5Qniuk69sUDzQ
QG/6NJPmnT2PUo/NkMdBht632KT8S6aX7ZwtdM4GcrspVXk58x61WuEdeYPaql9k
WAIAAiAqSEwNQ3DYTO3AkKWy6LsloJIRsdGJjgBImXMztDPYlAige3x3NHPAIubw
cNTK6KvSMOrzPFa0G6pxzObvsDhcHY0q2ePMbQHrKor4d3sfwvO+C2qGRIZfVSLL
ir8/z3O5GDJkCBrZkSky5jPbFm+hSE92gPvcXQ8zCP9V7giTKnjOo6yyR8fqOPGJ
6KIR2Q2XNOyjVlMRN0rZ+iXZjXYxRCXJcrN3XJ4Je/ShNwRllmI4n1d1TQSEFYVQ
hjuYFk2uCp5u0ALkl/pRB3iC03JJIUTIDyQTgk8iyUI9hheKcDDNe4qxzFnOhO13
5AzT3JPCYMtseiI5qICaKjOXlG6ODHheTycW668ZsV5Jodc9cd0H0NprExbJUaBo
MvyB92uoun6XEuUqQpZE695ZgzgbGKuO+1VSSq3yV+vF6SVG6CV3KPRfNpyFC4X2
3rynipOQszofRU44EcIs8Ox4XHP6cdqttfOdVKeS/1BEcg9htaqRJtMkLBjrI3N5
P14C53iFoy//21iTcCGIlrZe1HhCRpi1BX0COJdo6C+zBUly/V7763mSA7BXbXbq
+MHakw8OycF9YjhGHB8d3ic13xAPyfWAwoq6Sw1dYkxxeNF2s/OVHxgZMCKtXD2p
6fvoVCHylhfSFIHJyo3uhgzr+NlP2oXcYvIVZgeRSo0xPyi+ahbBAM4kbb1dFm7m
993VZUWB/keeKWO4CyKMKB8s6PgpFkwylWlVTjakg805BIEXr57Xd3KB8Tdsq8cs
2jKQNMY28SvoR+ttZl3OJ7Nsv+cWPf3y/o7YH8JGYYeFoIOFaQvW2GvULD9orztW
4/i+KefztTu84dmctD8sQuoSfVlrUMsa7mKcPkCRG3eKgavp/CHC+8mGaD2+ZJZk
QQ5kQJn6bN+sKGSQdQ6IN0easIN4M3wEQqQSE3zG1J3MA2jMgZ5PefYOCXIilMul
m1ppt1YzGiPj9ddKadhPNhpOpY6ESd8GpkEP9PzFxtBTq6kwsi3y6rkjRauhSuun
ek7H34ceiM0EKakYn6W5N7aqO1xycKewbmjlQuceWQ1Mgc4apsdKyqFBBQyyOQ4b
wZqEnsq0R0DE5DNmcCncMNad7EA+O5XAnkj4uKgJm5s2z95noMPMggQfviNo0+vs
FrZf3vqVxna23x7fpgNkaozIj6t/J/UinhQhsvkriGjKGW4d03gmgIjYG2IyAVYK
WoktBeOSXgcGUZzJh96Q47ScjRt0/iiMELL3YIleQDTHCrCOtRChhbuNury06OFt
7iYRO/FMit7F4RPrHjei34OQ9v3hwWdGvtyR1xz2V/5H7HXBByij7PqJvQlktAFa
fHL8QYSKtIbkxWpxc3lyxLyugALhHR4W7Xo32O/sH7u7XzAbZyFIZLznmK1gyDTI
hpTY3rP91fzSsnD09b7PAZH2KLNJ11w+YI7XsC0hS/A1fhPCQy2OKdBU0TWOCaQc
CgjbRDYCnJtHMAjhhl5MUtS4p961CAtok037boZpuFp948ucReyGwA0FiObNFlGV
YOOTtGiwAiNauRAeQ1pWTjkOhBIJiNPCtKOZDC7M0Lctx4yTh/w56MRa3NalXssE
kJnFAMPDvaItB69fJ3kUnAwSj8Wvlg74+9UBrwxABTMuNvRSYKbJBBRMSCS9jmRS
csT3pWw/x5pBjgfCyEph3btKHlnCQYg9Ad7s75ZG23StTEOWTuBlBLJi0O9NP1Jh
vc6l6qwGRewcmDY2k/JDWW/pbDqoUfthVB+V6mnpfWU/uAGQFNGzIeBx5wJ0h/kl
EsjxzTKJKRvJKI+2YMtU8ITWn1NnuSr1q/2FLoYxBydCC6Hsw1hFBDnwwK2UfBa5
o9flttchmPwrUmROdS8uP+Qq861m1UQkZ30dN6JYR9OMhd0mukLBJyDweCVkJW/J
n5MYGlf/JD4u4qsz+lgF8rad24p+vxuWJ5rY+uGxdJavtlZKmJKxOpMvZHm+Sp+T
9zgDCnhxUbB+xvFX4/OCUpMgNcHoSO9TltRGAcG7TL+lUVIF/X2VMgFvYNgpMkCW
Fk498N+14uHIrkSBwTnaKFc8qsvLx98X8jP13gLvQ23juP8iTqKVgI0xKj/ruOxe
PkZ3aXT1T8Xl5wjlGCrIfm9zIKEqTub7mpNheZ6jVTSzAREjQckVdx49oIP4Cuwb
+cCUooqd5lQLOaiOcphJP5FpDS8emqRSPhPngXoshKMt5OUF2VDy7n1qtTjpLkNm
ufDxetjKH1BfgA3vOIQaPBEm0/sBtfu+28sRmqnFTXUakNm7l+D6PX0qzU/LOoLE
Nu15Q+Gs2TBaVtMWqWqmtjsdrTXUstKrCgzdyJycpOfJvJRgLibm9OwGRR/rg0WL
GpydR+9oeLh8uHfNnsxcgtVMoTiIgP0H8YNSpttX2g/1wtsNORQHdY+J5YNo/A/d
E0Dsz++2UtbYWlAufEl7GMCgZ8KauQ8e95mEYSfLYY7TbAYcaSlfQBstA7QCNF8K
MHJR6lMayNcdN4htiPTkINGT5crVoDDkdDI8fBi8ttZ5qtC1a4Qs+uFbX0O8FhRN
9QPGfrVU4QryMgieVd+tdkHzTIB3a2ymsaLiLbxX3OIrqnhxTehZdcN6H0DOL5Dg
wXqAKWs6sViWW/7ipe493jaVe88fuH2cwO3lctV9TW76Qjk3DNBkyQzeSNvKfiJ5
NtlCWeMenrO4Be3DINtemVy5qTwfxhatJ9rDX0EsoKZ4v8JJraFA0NZJ1WXL6u3N
F9Pk0c2of2ti0YRtsJzMvl2N35vMza4iIjcYcgFMGjF2yjKKXzcFOIW1L9BqfbbY
NCuRR2J3RlEAn2wBRTJmRB4MMlqGXU7JbaRximtBasqGX63AUjCNTWnIM10t3D7q
SdNf5tPSPvjWaB/BuK8+gzjKzBqmZpT6FH/+4NSL1pkyqgLn4+F/Lt+f5Apsceaf
yWpGH1m8vsi+FglkosvaxO1ToixlVAr7fl5bZQm+kYmDtWIVhbQ5Tf0aI3f8dCaP
mPI9pvIrwk/zHnaiNz30cZswC5pUlm/k6IK9TJnu4tgLX6Gx8QWXmLBMc3EP4ydK
JT5MtzAdnlt/9akxY2chfmIElhgyIzem8guqPIOSf8gnkj/a6rU56ymix1R2K1R6
j4OW4zubjUnystHXH7XMTQuT17kVU0wihmZ5ss1/sjSsUffKdpYKNFBOZQc0n3F/
+2Ha16X/s9yiBapCudKNt1zN4t8bGaNwXa7AVviGbeY9Y4NQEXjNpT8PBumj8v1s
4lQFB5X9Fik7xltnFYTVjCZBZbuvDGsXSVeiogHpsfzjj2GFIA/uKgPcG+EdelNb
rx+jbZbc3pTb3qt9zGoveIAualU7fNLRnQeqfI89Xm4FGdCgI2/LmhRWb00fNITf
QWdSUOrob4E06io6HYl3xfpV8n5noHa/3LzT3xDMWh+41u3FYy363bbvJ7vxzuYE
x1CuGuxbKol9qoxP+ax/N+uUstFPUt+u0WrZrMzO1pGmiT1wzNR512VIORW7pTQr
04vNieVrg2SDmhy1r4kf3k+ezY4YX/0sc8bifkDUzYhbO/YeIf9KDCV2JHN6TdbS
2MDDKiV1BD6s5JQUmOgpk2xXPqGE5ASnu/MaAAs5UeKlbaBxiNxB2VspEfW5UApB
dhQ1hgxAkirJqiMmyLW6k+o2dPe52DNkCBRL4CBV/qJrACbJnLPEQ+b7r8eVNdft
0P7HMCV+zsF1Nvx+qOTP09cmnkUy6IrPRvEH7eWRS6ETZ5z0muiJ3qJGLf4W+f7L
W1vEERevanvyK1+qtXOILuwPNNvtZHj/8dgd3po62wa4DeaSzYPAq7G3+0Cc/FQD
bvQzcJk5aLInQZuKmjTmh+WuSRteZdGA8s9QfC4Cz+5tKcK+o7udUOC5FUHwQMnC
QBj0//1T3pzCVpfmXRYGv2ex1BwkMEhHS1+5OSfMlFXSzBX+G1saEgidI0XhOvt6
w0bDltwgBBMPdiGR3IOCn/Dc5lLov3PDd1x5XvE2k8LoHqRxuNaKzk6cGeSLIDie
rhuk7awLWuwAh5/3stPth4aZ7xH6yUtccNxr7hd0+tfZFB+L8d9jOHMvCZkBVH3X
WLOhjKZjI1CBvgiC52RQVADZexTYSXJTp29K2ogSxQCFktSPZ0brVkeZVgLI5+AL
98858NBMURYei4HbYMUMHda/NatpI0SgSdGL9COS/EilwhPzVWE5qhgLCySW1j3x
2NaOI3z9UU/44QUIg+ykQWrs4svQret9vStvH7XTDb0wsPLTH9iNq/thCcIytVs9
WA9l2B07nT4JwuNpf7VnDZg7iuZQ1AxX4TCsF1g3VF4tYFDfyEjfRiSAG++smMY9
CUX83iHJlY77OEQRpOTK3TALFl5NEIadwgNlK6goNTCMW3mYbEjy5Q551ss+8620
QncjqMqJR/y6EiXVe7iOXsB2HMp2JOopLUpTYIgrRkqlzjAqKXcMGvgGbx6GgfCR
+cQUVU1sgPpPML8n5q3G7hRot5LZO0S3kcVrv1cwkMH2fB3M4p654738y4IXh2oD
2UwguiwRhHmlBo68UXGAFOaEJP5RLU5nxO9q6shaTStF9x9uVicDH4jFFRFgm5IO
RuPWKTmSVZQsQGYXlatVUuHgoUFyOlteSCLiJbldOk4x/5qEIdHOYJCr3i9lMHSY
8rgLdXOJhvW+ZmdePPBxndmUtjHo4X76k0sEGds2fCNvLQRhStuvyk0vhn7j2MdN
VyMyaSs3Or/7zLrXBTPKmtqk+j9PyfCcOL4BxskEx1Z4XfSm26NUa38yWO2wESz3
0NZtxC46kkyuWb4ECnuNb/OwBKSzevq52MsrITX7cJGsYa3rlp7okZgnIabepKBa
wjxw2+Pv1/xfv1Pks0Jz9d1/XlWBRMGvDZtCkXE3+4niDzqHj5rGcxfYU56+ZWSR
SsBP3G8/WgAmWFK66GHze8d59G1Gq/n7APgKZ3Ts8+UUYBZQyAKrJOHC2rYBqaaC
mRMgykfUsNwXiSQzlBvdf3VNczuKaAZljcd2IEVoagYh9GRW6ZluN0RhwMwEABJQ
DIQ2iv8xe0RSVtYPoLAoN7pIZm1e8P3aTwrjDC6PaAFp01PGSVQF+LZu5RcuN3sO
7iK0uxQz05M4rTLDvkb2+thvzdGMD+vSe3PklYSrJhh/9Yfhhkr0C2rXCkxVk87B
Fd/ZVRSy+g7ClNO5ab2VMNUNOkM5a1EEn5F6eiuGVlj+Mq/U6AfDNi/NQtVF3Xqv
3rZMKGTmSP6s+KzV3syJm08mh/sHmC17z7JPXBEbk0IEvi0Ib8Rc1W5PTS62gEx1
6JHPHUqLPiYJg5pBfqnZ4e6XDVEB+hs9RW33KBGHv0STSyGmikIdtD97c3wtmfKc
5LT7TLAAJfXC/ZDLPcmOkAuvm+4+vCchU3+8FCkZeGSzVp7z30Ab4ZYe6ZkeOg8k
nxXedIDxwyrWxF9TZ3P0Q1CFccS9LWIfEz4OqSOg+cjwfHWN60gOFPRfWM24Ozjs
FE99VVykKepiYstgV/pOKe8FcSBoLNnu+Qm8qAKa+IP8SjeqyfLFBr96fHNfRJ21
C1/XpsoKuGlmLiA1oDuRImMfdp8LXU336azBKM6zdEXEcFMkeXN4pzzXgpT2L3E9
VMIHUsfI6m8dLnKHFpIueSGk+GVCTluCIZcmv1CmmCFq5cPm9a0m3y4RFBF9BUTi
8K03Qj9wKaRCXcHDmcyBjEO7kMR9HxJQc3twq/qEdjDglhF06EFgcjZNaeu45q2e
pUDnKnGvcVrt7m873UWUmVpW1ol3CuUtbGXqFKt5tOlA/mXIwieUWN1SGMERkzw6
WTI46pxKbZU09rHw8KwwcwajoBdXcm0HxLa3bSgSxFJ2FWwfFaVaxEdHld0UH6l0
BwUh1A/jJhmvx+hN0A3oNVDi4mZSaJoEAyUM8woaE7dGkOGZX+kHa25HMteMkkGe
HsdH68gvPLeQHL1gIKKk/IDyPTaGAfeHz67HSGR7Eeg8a4wMLpRb0rZznE5EGdaW
3LLGT4/tFV1xwxHIrVKwUbkOOfZOMt2r1tzzEmt+EcmwfHuLAjFh5nCU7cg8rZNw
X+ywzYx/REty3Z5GAL7HipergHMUiUVejYEOjlzVRDAgkWqXoRbKXwBYk74zCEPf
LS49tWxsud73gibvjgN3lBcE38QqCQutz+Pi6RMXJzy481Jebw7ZjVklDcFXZsYP
16038pDZuhmP8Ebdb8aByo9bURqyioVt9P5l9v9/opze5R8foFyR/4/g+fcNNM5Y
9s/3xXQ7iLLy0+guzxh2PhOetGb4GvIy+7PBhMWueBYpeBIY1Vdq0/aE+LsHdOHF
fhBz/VK+1VzPYaiTGGY6u1r91ifPOYLq50sRt3/4WjSAfUzSU9nNLxZgLdzud7qQ
/1w4GGU6bpdLxGJUDVZYSdmGtxK2JYYoJ5/A8TFm8SUAthpNe6GR7TiyQkkhh897
0yMD8zzoAaJARXY+pXW4+su/5vNEOSKsempAA0YY73qjmoW1scHI4lVaNRdc/x8h
tRW9lZA5ycy3oi922ho5voBVHW9qnIWwJPxWSPS203LMrvJ9GvGnVdzk45y7d64U
d4/mn1GTDzZ9KjOxX7n6651sI3lX1a59+DA6CIYNmnDqtviR4CdK/hbWVZ9rRivQ
7s5DNv9hAUZrV8ga5PT0rNqiHl7IN4MWwn1SRACXOHDHEmLDZu8DRd1TIzdDYe3F
6nFQqx98PsLwCLcheyAIC8okH/qB2+58LieCcw1A/VSdEHCFmyzVUX8cBOYXw5ct
+5NaxwApH8fR2xXfiwolStsk2YZjWF5yb+aQDwNmjBHz8E6XkojAWNAj/XNZZgvg
Ydklu0lwrvorBwN1A5g8eKhgylnqOSmAEahr+Cklahv302jL3y0e6cYFH/vev7WD
9Anzjyy4uzPWFKdw9Jzy08ZoZwh+7jy6xcPoOnlkw7C4Pd3O6MaLGYgz0UATUjBo
o12gl4gSfTDttf5Kogb/MogFdP/ki3gPO0IzHlqW93RJexwuIsio5zF+QcJCx3G+
EyoaByArDiFdaKum94wtk6/KPMYe12odi7p+kQWCngvdYwQvA0/V4hGTYT6wCnfh
oKmysxuB+AHebcOhH2/tPsEFNTyD2iJtPAw9RpEbHUEPiyimxpsxSIMycrcrsVFH
9oz66rZfdpONvQXKM1uG5VJCzjjgjn6osV8lO1nPaSzbNUBT0iu7FDgMbAlnaN1M
kRe8PLgKVtpdjMZvZbUVRPINvyG8Ov+LbrZGDDIWEJuOPHz8AZLBDbzk69Wird18
VqamKoY2orcB5yM4EbEd76xPC0FnASB6RDZLKokoqE5DiBuo0YJSEsqag9V1+iQx
u6X9Z+BSkCkTDM2FMfFcBwpGLf+cMIOVZLaGFaXF4NIoMN3W27LUvLZRWFoFnqJ4
T6QdBd889InmWtvjacgM28P/zgO+w1iAWsSzAuKpdQBNG9rYmEn/KE5yDgHovglM
XoinjXIsltxTQEedIeZpFvPLKzIJtyVSEUKnzAYXJWdOEFzoI/H5u7qNNdNA7n7/
z2Pc8ZBHjsupzWb5apIVLXMINsfYKcCOqwpR3Bc4XrJ5X4XvpQKyiwJD3FUc+bQL
ICLFUcASKUjjiIN6C5zGn4bDBC3/BIejM6T11XeC/ank++mMnRIkZ2n7eAPfANuA
U+6KOJKTFuM/CsDXgL6UVG2aoxT7oIcfkH6i//MEVLe2umzI5szk1bH1ACkq65j9
/oGXf4zeRHjEsnjnRYOSZgVNSd0H4XdtTzLPDrfTs/5+yOy1+F69aEWu0MQn+EPm
qpw0ePR2HrTC+smDlO3UERWigVKoBJ4AyPUh/3ammFE7XY8duLLizNq5Gzb7xiC1
3tQVWSOWHtFF9ea4AZhZ/kJ+aSetGMG82jY/3IiFM1XJlGYqPKST8Z9Nf6gbMdhq
hZ/1wsEvo9gpw5cmIhgm4rUfvk2DlZzWoNbve/5xBTMqv2VpzQw//Z1XiWH56T+u
/pnaHG+fQyBFSmB1MMG6JX5sKhPE0dg9TTNrhln1i4igtbKVpeOZtpgfT8S9Kuh/
wjqaet5mfcoenUk+oKzrLAKUtaK+utSXhJaqXJV9RIkGLoiaGOaHesPf7lECkcub
Jnv5dTXwRMc+/3JIvExX7PBIWcrdV2cK5+GyDkn+/ojcUHFMHc9AOkFn2dVBBDs4
LNGOQnGmuw7jKMY+IyFYWI4RNuBelKxhP4LzmEtFBXvybuLX/ZnS5ZUcJ7JvnCw1
fvRDw9mt+c+31HiZ2vyVi2EddjscwqtErJNWLAHF7RS5YLdGumU5mJUHEmFWxIic
27b5iqrlgbbilLcAG5R7R/9McU4KBAeFN2T0EPbm2/5MrGbk0efboEp5qKhXx0jC
j+cGKcXdJPU2VE6c72W537Zv4YYrfEbMNmLW5ey3Bfl9izGf2SEnubtFEsK1ibzn
DoNDBRqj/22CT/mUuaPH50Hm9R1bgOWkYJQbEJW2DspJR4M4I5OHfd3hS0v7ylWw
2t0YSx5YD8l1w+3bo3dj3GBqRVGREBneXJTqCTfmiD5CHmiBv8oJ74/jZWUD9CVW
ReqZoX9B+E9c4fDon94R+AVprev+fzmuBPVh+SuLOWEniFVAWP+hWWRF6nPIruJF
6L67kMdfsBoLQkgsY3SfEVU8XQ3uggJfhPZSgpqWc9DySmcVBaigrE1wQFQ3OtWj
LVGKJdBLigy6JTut08wJmMCui2Zvg5LlFS4OatBjtOdb1ghctBtTApJrvK6qx0Cz
2o99/KQIsF4us/JdeFk4T+K5Y/sndtPbVlU1LdBO9OWr+7zDeQWjpeD1UxALJ+oI
cevfPdvYkWXAo/qB9OOR9/xnuVk4sTClHMDSBR0/haIBvCpPtAz6p5wrLuDFnLS+
mBPLv1Ev7HB6hndoiQXwnAifDuzFZMfHOIOSfdQCzopBa6LDyBhHC2H0tp36d741
MJfnSC8NyXNB5L8hvveEZMYvXnzQvjidVLIIYhEnXGlfS1byiq6ziGuJO93mjGDN
6f12CdMSBiOXP7emd5XiFYp7abUnFhQejOENxoyMc9tyeCopoLsQsgzWJSWBF63t
OgncNr+6+eSTmogYFi7IdHQpfmfHmY4nn1rsRoyjDxfcStGAbZYMiidM2X00oz/3
hUfPohEZGGbErmrBgM1wYsBYKYeAGdhhcFCmp1qaMS5iMOTPgEAyzQgSadGjwopq
E0l8FclTkCRV4u06THmVeiraF4qW1bs8uK5j+RHUPioj8zSrB2RfURn7Q0jbALSg
YwsbOrI9ZarWskDAdEfYICOT9CxtfKDdYFA6ZqOWzp7PW0hA2R7mG5nuKuBxAr0a
FPO6ZEVz97rt/uDDhK/4Wz2TH0AhiYJe9+5jw9IS0LjAAKQd8X3Sn5yz2J02TyID
tqEbXQ72a90B1sAmd+bXw5jibODjkiQOW2KL9J4oj1qe2HE6oEq1e3z3lzEaxqqX
QrNNjqpZPB2Q/hEMNlkPY4EQ9Lj14E0GxrVaT9rEc0Us/R4MyCJxE+ZYbXUFmGS2
7ylx72o3ji6CYJx5BWsffrnBZe4u8kLH091361Hxk1mA4HZl4z4IpEzB08tOD4bo
khJpMl9/uWPLV5g4/JXhiRcMPpdOxfIfR+12isClzeI3O7wy8VJs2/+3v26qA25R
nUJc8q7o+4qLyit5b8Vqnjnp6wdoBjSV8ol0u24r0dxwQAZpMKqY+u9JtsY11Fdf
LfXpd01C2LYVIz2isGt13LOfK5ioP1vcUkhfqo7KuMb15DzpSH5ZFQGRuyW/YzqQ
5MkLC7HvQ1HXmvvFh0AHz0I1Kh0o7Ynv+QadvMY7/TioOzBSlkp/ZQA91sJC2LOY
PlapMYw6UdkfZDnKst5b8nzWpapoZBRRkhhHnH3rCvSrg7Imo1yUCrz66uMEg8Bf
iegHJ7pr4EAExy91CVFqyVibmVWHuYmA+++UAnUObtc7knRNpgGyva8rMLdJenBH
hJ4d640HKAQhIYhl/84CTyrPIYhoi9kpa+xR6/ilbXVrh08htlxjg43t251CasJ8
D8AFXkMYgVJFB7sIdUr20vkDZ+uqn7BCGzkiz5i/d/N+2ot7jUvpqHC5doZmGnvl
Q7lxR1FDvbTP6SOcycTSMSDPks04oNwZdZFeyQUgmJU+CtmuLZWQWBmlTcUqOt2k
0RZj+UiGIABYwxnVmGz6bWgm6IcfsMQ3xi1eSnVfYTJNQ2wUaPv8nh+ZPcO17Jok
7RE6teNEwZJrVmtWb5PWuMGUxLwGPyk9thQE6km8zNAYZWLfFDP9xO1C6Vn7FWV+
auwzUrFOHdLQw2RQdLqNaho5BOVw3nfM6Q4c91ZQcAV7wMQqDepSLHwsUV/hIF3N
gOEYo96gz6WrHv8/AxUZ/faO3fydTLjBiVUU2XcKU3RnVzm2F1W2geSrpS8Sgzrr
jogrokYqDNJxhopaj2fJe5atVWSXThvWawk9bqzyEVtavMRvOTtzebxsbH6dn9GZ
Kgjr9PnnNPFgX9fIxuVFisHeO71NlYh1cJbXC0d4ZMhHa6uC5NOhUa1DLPr8IM/b
ePUf5+GRFLoJQ1ZA53oGjC2Mm4yuuzIyptEONGyfv0h+Imd6t4A+z6NOcMRRwKWM
dg1LBEm+42MW3Kig5F0ypLBdVqP4+lSusNSRJH/bYtILhjOPkTR3TPCuAvjd8Htl
eXqxBQAv9zpI5KrjIV352zqH05ked5YrRS3QAVJcOweSRf/l/+2xTZTq2jfjKvmB
n3BmGqhXHVAqgkPYB9F12eL/djz/dJI4XFff4R2Ruzf4eK89pXhRqNECiyGLThdq
s/gTk+cCd8ZxYvgzrCa26uIcNuZSz7RL+cPRxkVZfAKFEn5IJtz9XCbe4aiJ43Yb
gPZvJDUmHLTNATaUp73CCyc+PH0GndXRKxsv8H+Ciqz1ZKkB0lIrc3xlUADiOMco
fK4Z0CYkUbN7o4J1rIkbCDBXuHA6Pl36Ke82skkW/drm5sy2iIsH1DMGT4Vefybr
XW9L9/7ZxbhawmPXZLeaJ8UVSDM1XNFaiJ+IIDWVtoWe+/3TZE8Gf4sydURc0qby
7aECTfrDwf7J5zX7v9rYAfo7OX7h/APSs0sOVetq2rAlFI2o6dcxeVAa6Eweu3mB
/RNhjvL6UlqmbaoqDm9WAbCkKdArY8KYm8p51vEk8abVOHf8bQlATIcUJNVdx96p
eDad9n+kTSAH7e3l0+IFoTPOaropwadx9kw8Yu7vmwYXk+ThHCmWSXLVhbX0Wz+V
DsGDJv6ZzrvQNstLDOBa7T68nE6U9J6zkbEKIUAF742GQZrI26ne6fFu2Ag5Stqt
D22C+u8VtcLeOB0HYZmdM6+iPLrsRr8VzHgvWHkNpE/iwd7voiEjQdp0ltlxpLah
dAxG+zKVKrjGR0JsBRvxF9UFQyHOlR7ghRAjLAD4FaPZqR1ggEG278923+fol8+h
cnzJiZz4V8wIn/sWNMgSZ15waRVEdz+q5IrqJnYcuYU73ok0Q+Z5M15fM2H1Zbxt
uFlli3+3vIA8vA1gURBr8vWZyLLE6wbL6KnPFGR2Ct3H3I4yQ1XdQT+kH6pOg+98
h0rtEJycfhIU2pu2AC3++5a8NZb49JgVPZIemmwvDy/3HPcwPeNLcnB5fPbUzGDY
94FBhv+6+OR2lxWiEpaoN76ECwme5MQ8yxhfMUcfvdgewHrYlWKUYtXOIcmf38sb
h0MsZJ2cRFoGELoxTAOsyqSxCPD4R0xqNhn/nk5ZO9Wy3y/ORXv0s/COXcI/jCA7
OzZR5EhotCXQ9Qp158B3f2FIw6YU6HdM9AR6tOD0Yo4fV3iifS+7E8wuDnU2mXNw
sM6vW5b31TVvnuLZB8Pppcx4OnhnyxxnlSvg2FOxJvbFZp8RlP6IOvVsJqjDMSLD
6kr2UgP2hW7VWZZdFYc2vNumVYX6btXDJkTRV1PNLAU644p49EKoRwKrr/ys7JzZ
ewLhx41v0UzJF8jKxmkDiDpBfPJNg1rJGT5ZbZbg1gsIAztvAQF2Y+L9aGJwiDbV
MdVOhHGzj6fNNH7F5mflBHObxIGUSTT8hXnX5Gg7TmCMmnecpZOtsd+yyz2Nz2yb
AjnK8TbvQJ5k19RV2/Weq9aU/tou6qIRqm0iict9FJGERK9+HT0jD+dpqSlVpep8
EGS3tcs/n6Ok/aF323UhSbW+i4DYkD6JCjXoAK+0yrFJayVayNvH12n7FcSTECke
tJ+/P5uOonVuj31/gs3kPTKxoh2plr1t9ijM0zUyeirqxufWeUwm4fnVk/1CpSyZ
c1hnxIiO3ycMj3JS7Wgek34cdhcOQb6EwnCG4K0gr6RopxvOEPo70yEBb3K8jpdS
jHc3JkG6MrJAyKJeSTAuSk+zYZ1LArJsvKvout8V9TGggXweKdvXNRsKQHqJ+W/b
Orh+oGjWB/os1Gclzr6LIC45j3np+R0zJE3STc4VKEnsT4PGXwjHMxj/8PvUaHlG
rdxsTj6oX/NMzxxetfmH1Jn+H8HPPLLoOuEKD+Ob1U7RoqevA1p9tQbm4sojM8hj
PaGXrO0rMTIFiCq1cuWfmSOFnpEicbmjNtOEckCoTDGNKpADJo0wVR+eBdLVKSmc
Q4fRrG+XtKYw05ciczv2KDso43Xgcl0HtfNfSxu5hOkCWAD+N9cYmXXPcT9hhMVz
jHxOhZVFC9rSHzNtAdXqwakW92wPhoYZz+7wLQvdTlhV4LTOL/JrCUTYHQsp0VQ2
+wF225MbgqA5X0mm9CZR37iOE585mVoI3Iop7hESi0P9Za7UqRYQ/I0qoCnAVlTk
Z1mvAtcUw5UCXJDGk3OkXledRCW7eh/S5Q5j+wbgXBFc/vdc2IC+mM9Dlg4aPX57
xzL/XdNi+3cYGNe/sx43N/u99bPqRqTVVyArsdvRRPdME7seDSaApkZlSiafqe06
1lO7cSuDaIjI2V41bDCkRJ+Y37ad2DVIEDR8RYg3rgiZtUih5GWlvsJ8XfHn4bv/
CUjQs1DYKwFZmUPL4Aq+dPJR5LBWfAt3Yv5hqwXbLFJmroK5dRh899NbbmGrVdp4
ONnZkDsyOF2worD9L8JqE4Mk8NWRf9eLWcfnDMN7WXJGrymVeGwTl5U9jwVwDc4B
7dgpFVwyDpZmYBevZYU9ARsu1xMVdjxfhUqs5VYc+R72f+ykTJZI6etrj1v/uV/a
tZDXy9/dlETKMCzWX0YGIxSOfa5vOM7Oc83CvAFIWXpNVqKGPjW1nI53xIwVA+re
/Suxq3ycM/DWhxqJtKWxL5hCP9GbD+znjZALPypzAtFmLwZcPB3JAcI46QtNZdoO
fkYpei6M+D0V72Uj/fIYftUkB+EpsGgZ7TklLVf3Etdr16+S14JAU0HUxunN0bVN
qga/tZdXNGECH0XYHdmofRTxujMBZjXPU7XCYazWyP+AqqiboHFnzBYyrKY0wwC5
KHrgO0iz17jt05j4h8VpCrh1ipwJzpQDB6jbUrK/z/NAX5VA9AQZzupYBdt0XgcK
OEecXNslZBy0gDuJDNnbkxoica+iyjiJFNs6hLSUMlvWVwAsOVK5nOm1h5u3AodH
d2aQbuVeEM7LB9kexG9ePLzRD6nuPL06ihhE2tZKZRWUQQxZqOxgqax9XFkkr4If
4U62As7yKj+t4yJcSfJZCw+u3UuwUbSGhH3OsvOhSqX128q1HzyANoKuXWwU1u6I
fcDjFPO8ZZJGkwTObGY9g/5SLoLo56MV/fMTlLNS1dr/3w3k0Fb8p3Tc+KfVttNt
iPqJeZXI8GJi6tFqoK48zZsE2PG287kNLfu7l9zGfRy3AsxHyYy9VoEg5IAV1izg
Jp6+kjVbFEDHXGXu+qaZ3pBJ3/eTm5Ex7GGjwPuPQtKbaGtvKn4wRoc+AxtPt9xp
K5NmnNV68sJY50IY9pNdGGbGFxM2teJAd0gOOyUKcTBLn59OATNPKTKD4UVAHciB
tasUESpxTUrlCYEK0miE5j83A76kSOio7OG4PtyfVX7Lx4E7Ue4Pb9WAtxjpXBXa
3V94M3vTBtXhxKahnYqEXO1R2alkc/rD5YFeIFCd8hivIfJui+NMIYkaui0/9ugS
RRJo6SzW4XhyTmPSvxOCLuQWpILE+kaj2QX3JcQT8Zu0VWq3KbTFJBgMX2CRjtal
27tUIAXWKjTk1kx+nYcO5Wgrprzy7dsBzLnntgWQbuaZr7lGx0Nco0rmt7EhHCsq
XPxYimcd8o8jnZuls/XKsQnfKYXUKsjzPDe/BTe01NLPG4xoe8kYhHNVC2+ShIL2
UPRWi/dwWSyqMho77/L6i35Awqgp1Uha4lND8amHGAILtfwtnzosqkw4AkrT28yr
xsEVPOIR8t4GskL68PVzddWk++kIxxyni8JyIDz+mVJufIOUjTdkgUmnm1/RBbQD
ErMWzXBjsOh1cRV/nWvTB8Yw/V3Rjqa9CJTajCvlj4uMo47rkDbis1slUjDc9ipo
c7Rcq4UVYt6l7w+ogSEKXESP1IoV28K/N6Azza/u3MUEhwlAtmzY6hYLDSpwdSKR
kHkOh/Pw4TPwfCJypv/RvISkaBJeLR/5p9WYIXL6zSuak7AUFb+4OPvtk0RmFSkc
DuU4UX8+KjBWAaGTKh7hRWRWk3QEJyQPtVJXmGJVoSmooe2JBymohiaKEG2Z2CKK
2wyQWgxZSGw0+H8Cf6tioZV/8SSYwT0DlO2pXoICrONsU+x73RFhsBgkaDhIypmt
W+22SFv4mJXWUnb4Upbkd+HsGlo+z8n1trXzVIDjhF+la+7brb0L2q9a5zMmscTZ
b4AtN2EZWTxaehH1bHvAtLFMrl6E4eZ0r/6eIB4UAnLiIRvC9vM3I6hWSabwLF+5
fOxrInLF9HLl4SoQyTjukpytDR8LT9KPbL73xOb+iRksPhgRrfrXYOu7cRPk1xRb
yDalUzyjerdtlvEInqT5z5Wsap8ZgKGDEpXXq4Iij3d816ljI2KtIuqFhqrt/grR
x8VUdl+7A1Ti/k6KtCUc2oLOAy5fhHniIiei3DW0Hk3v67X5QScnv/5vQ8EmVSsK
CRbcpL4o4sjUileIpI8OiNoLiT9GBsFbILNaV5U/B2IY32tCfZPidwBuYMqb3x3p
dkfI+jNMfrPBGhhJdGd+NHI/hgItUp3aVG58jzP9cyFcLuuVP5BCd1mYKDhJAiic
pw9OY64QbXAmSOhPbszDQAqJILd9sFzggxXxWAW6CAiOuX72N/an8dcarMUociAi
kLSmilFen1F7g7tLhSuV2wOp/oN4WpkgFuvj0UXdUyqZnJijL27yZwIzYJnpjXE6
wknQcocQL0OR27r4L6d7spv3Kzi69ck10KE6aeAMpSCTj2yKrZc2WQvtWeQVn77i
EQF3DxSdMuGJv8gJTt7wPUzjeVQBeosRiVCkZoViem3IX9uPOe3kTLSYAETxG7ih
cyCC4MOv+f7YOdoSUkqBMQFm3MmIK1J757JvIzfSqYNbZxIMHT/VnBJzuBM3vfYE
mStSwMwsksO8gkwGVcKmjAkQ8hQVDrbhbAt4I3AGp51PseHDdYU+GtrTOGxIQwCA
TbT+Smjik4APORFEfQskbxKCKmGrM8b4oSDHShSmuN5r3d0xsefkGRrYocgomYnH
wZpZqL1g1d3uW0WT+u7Pvlm73qBGDigP/JrNCXyIh+jknvPwadQWlCVkq9YQb/ez
DUMbbHyPolnlUacf3+aaosv3Af0isrU+/iM3yAQN99MJOaRw7a7Uhe6S78YhDi7x
SdheEQ7kMEt6+speko9xfFEb2nRREhQqZAPpFGlqwjGFAbgjMWBXOwker7jWwqor
sneV5HXBqs2Pw+QCsBXwIfA5QR/faLzwL9DTI+/ROgk05G+2aEYKdwk8vaqZmeDF
4r48xCl5cL63jBrhJRKQYiN72ReBccLXCjRzoK0moEva71PZUGvt3NPdlS6j3sp5
WRj1K9mHFRt8HhSYDvTymzkL2fO5aapWen61vf+BV1unD0AIpohdNtYzYnnI/CKk
cvJCX2CwyTQHAop7wCp0LECe2ZOPhe7AuvvEnOnR53z4lSIVvCSg2WtRPYVGARC/
fmmg9LNvScBtP65V8elkJ7fNixghoySux265fVODZt9FSSWcEfzyPJnW+Ve/GVCs
d/2eDp9ucUcMg/kevE70NdCr71VArhSgP1sA9CwvR7SQGUDYZwMfGv2QcAOTbBwJ
1vyPQeMYAvnxRUlg5N99u6AHBpX21n49MIu9n/+KGoB48qR6gVX26GABIaMrNRdW
3RxRPppMBxqph+hVnsNw+GKPHwIPs5okMBP/S6PNAuVvXarltvYBaUHEona697SF
Ona3xPzVXSG5wpxBRCusMrouGUpE7ich3xImANwcO61Jqq5WxTd5MUJ7UNJSRupB
yDXdgTazU6gWEsHMsOZYULLncbmSkURhkVA9GCLDoO/0o33wsNZetA+XYQOxKOSj
B92dyz1inrrz69uLWd1V8GjXRivmzfnKN1G2hnnjKwpI2mPyJIF4ns2H7+D8M52q
B/1mHFE3LNGsW5MZ6tAF+HbwJmLOb7kHGKRSFQNwaZfs1hKiAGGfrOtsCNG5czJe
dALOhcKMZxy4U1HOox9Y6rJhRwoOhg8o0N8kwIsCldjO6wpx3HT2gat9RYZtdVti
OLLgMIwLo4YeV2EG0yQUPl5iPOrrSQS5iZoLSLNf6OoAv3Iq+RRKtysiodoB54rH
Vz7hYcA7FsDwgrZsgpMh9WujVFeOlYY1n5mknGiWX5MUNzG//fvSm8/Aw/a8Nhz2
/4TZeqDgczCLXiCGpPiu6IvEd8J3nfYl01fhRactFTz1gDeUKJ+3Qm1HAn56KxBm
m35W9PYgVcdtF03dio9taDS9x28WIxn60HeNY2QM/3m/LtCqDKUF+XJAxGPwP2js
5czMtIUU0GYbJmgPkyWIvzClAyqf/TuQDGfdv7U0Q92+BQo0FWQeJ7UAaW2VJ3PG
srLlvysGB//nurTaVyxT1gtbqaa4Q8A5p87Nfd6ycXnjv+tkw78KzbP+Qu3siLLO
WcjrDyaryOmBPMbwnmHLSGggdpWa81Z+dxItPG/9niPIa9QxzFPTSzPtBcD6kwlV
Aw36EjSu+9PXfYTHaP6ygoee4au1gk6RQpSCU8vNcH61PWwm8KZuhS90EiHuoNaE
euxxRr2ePiZsol1M+QwaqtE/nkf7wxaygzjTqfq2+mGt0mZzY18A72GjciGYeT5r
h0/o9L6ASvfhXGNd7AfcwCIis1N1/e3bwX2UkTnI1Sg7FC0FJHkPHJGwGFqwqYYc
esgWANYyoHdWYwgOddzHCC80/1bTlF0ewn59IzOoqIczI1o4qvyDI131rFpDbjvf
jUqQqyorpvc2c1XukV5vUvxqJO/NZlfOVyjNKH/iRLSxV+lzUBJXaPN3FURPLTQV
H9arhSXVNcEiH2YLH8LeDDMdKHZQwRlKSzCEP1DCIR2RhIj53oIff5hlhHVg8nfm
3qgTyKGtUZ3CwWpm9+GDCSPQsEy0oclAi+K59x/HX3dNzRR5R8COw+71ZPgRsBDW
P6/7Q/Wrb9ltdo3wSbw9YZSNlxyrQkd6QeVkOorDfqNoVDnCymoFfWRzEDoADqKJ
KP9KfQ7Met/MBCDb/c+8RAi5BdbON5uL3Qn0BXOQr+kdcsF/rcA6lOh1PltaV6do
DV9/zr2uInTAphOArDVbEQO8AnLcGkEeppghDBk2ANqt7NyzkWx/74xi8mfMwouk
cSN+yxQgSl8iFgv4cQcl0l6LRVq9Zi2PP+SU37m/tKcG/KelOgjpiSYmOaka/0dx
KHEu/EtVqSzSGTC+0t6Rfsl5orf8u764qLwIXYv1u5sZ5CSR1iVrpiMNAgbW13X6
qaYLI9nG/jSFvIl2k96p463rUDMJ+4FPyYZYoue6w9dDd+ueCNYTuOjYIPEMs46c
JK5/w+0z6BEyjrCociE7q/84cwowMWMSyMRS93J1K3zVOdGgbQl1p553xC+L2R2e
wSjNpAO8pW5lyocNYqgYvvTaywgl5wn3n4HxDWFRa936OFV2GHs1keYbuhrQA/Hr
p0uwYd3UK5eLRpKZgY8U0EuAC4c+/67BWx694mXZpIpOFZYwhtCbObKpgG68YY8q
t42q6xcEShueh2x/j9DkKII6qySbNXynrKVvOYuZAMqjdnIYfQMbzPbiDIu1FpfE
moFcDlv74Z04VxRh4pTfl0qLDwYAjXzy135uP8cpSxng13r5k1asW9tpuFYthY+5
t1K205p7EgcOOGlBxJTC/zpLnczWNox/9RSB+U87RUK9MJNDaZ7tzwFIKiOEiCzA
QIhTi2mqwol2/C4uW1ZaU0bLdqYM4fAhcwNqXBxwfm87kCZJIBNLTiBddBbdPSC/
teb2PSLfSWRaMRlzwvIwLeHAyhHAueSzvPO7x1NKIcc5/WEMldoGntaKnMY2R/sv
NdOdp21l8JFhncIY+dawhen0B03IbvSl9Znnt89UX+frXr23eI9k8STeG+IDrVru
`protect end_protected