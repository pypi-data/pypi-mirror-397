`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQMy0Nic0oPYTT1PeBRgvHfEXUqe5ezCWTP7/1Lc6Tdzk
shkulhf6pwVuIJD9PYzoYEWdnbtKTlCicQJUlo43ALyWUd+3GN31NIGEY3Ok37lw
Z75t1Wb/XSUR6Ix1ZSshdUUzm+VVMUTVeROkeMCPBsSeqcqV6mduoPgbtE9O0sMz
JSkwl7PLVAJEXxx/32F2N2UcELoOg1BuIJxRGgyACP+lW2xZ54xsLAee7PfHDamF
oKugNayaTVzYw/mYURtnS2iV06ZZEyN+yYMxQJAevBYv7fJtW4b/hsIr4hZ2FCAn
pZlHhU810Kjhp+aMeJN7sh1CJeUFn4iXZp1FxDdCatYBZO3eUJ1PtCnSrfcjs45V
e/W2ur0qczU1tDN6+EZJ+Hnr1+d6Wip7bgmDGM/HIWSibnUrIFgDSFF8cfrWfK81
IDw7L7YF0W7qfrF85cuNfJo6eYWhu9jxni4ruyy/8vNNWOclVc8GxDmAbkGKsT8w
eUcizBKXD1N8UwOw16IizOGDu8slclHHshtt7LdO0U4sdlYflrV+rKE0eQNa7dHn
qcjrPEHXiq3TgXYFdu8udwiYgBwpGsqYbYOKUNhxL686h8/2BK8bgUkeWXjsyrql
mkspcX8SNFkf3UKg0QuqOw4t5eoJgPjNUaac+ZjTWjJis+NdSZA8cQzno7Tvcmwy
nr0btSrtGNga7Rxm8/ILSgCLXfJ/Vpi/7YlT11Xw9ibD7Sxk2mXZwnQdvySvEi6n
jm3W70/Hjhq2syyCdKCcVaHhyNRqZZwEAFcIMlYvpT83visAbjuEqCCxmCiZ+ytT
KwZ+VzTQgIiwlIQYcAkQUZjoDaZrJiUlBqTFXuwBlk/7SlodnHKAqec+94v6ynRg
uI+mz3m9bwpepK9qqJnVFNrhJgAKXnWO6GdjiPAZC+//dvu0q2Gn/Ru8ngfDLp9Y
uw2jSnkZ9V01Ev1G43lw0YcmURTyu9D1PfxUtemM49kMFUIL07tguek4XXaY44hJ
ONwGNgowm4QlgK/ruHAR79ZMlbKFH6EyS0hC1Dh6lusDJH8iPpW0NEo6EzN81rPN
e2sOVKSg22/6tU87TzpvCotS2pn/UgHSuZDOlBpDkLTYbVuSwqWbJa1LhJdbLlBy
f0ppQlateZgkSVoG9R4qEL/IqJNeu3OD52AgbKlKT2/fQNKB1vsUlrwN19co9+XH
6c+oVCIR2WadcXnNGKbUOJx9kmyhapYAyhXzY2LMsd7ALO+v7/cdPuDHQsP3/6GN
T06/JOXjdQHsErkxAo4eocN1/9PQR6WRPwTRuaATfFSpcx4uVQEvqoZdcE1KFflI
jdu+vecNxuoG4cpRR+V4hJOVylIhO/5ZnDMAisRvfDvjbNrltGDEq0kIvPp3mjEX
Ys2O/bRauIutB/CZWFOmPTMeE1pIVNfEmdZaQ05A+6UHXc6ChYVw+t4fJh3riNDu
Vpmsm+6LsUg+AOrQGww26Q4wauVWb0ZTchmAC6AHNM/bxMN0wLjNJR791FTGyD1T
HOWnv5RKUTjWbsgs7be46Mpq1vjAfA6JrpPudIA7fmu5ojDBqHLfgw/ecq2mlbkN
JkKBQwjbOd4bcXx2nsfzthrslh0BvuDxD1uQtpgzqLZp9pF28sR+L2oPMPljgePp
ltT9QNJMn49OM9MRtryt+Rf6Iz7/dns6YFd8oCZAN/ovaosDgc59XXMvi3u3ump1
A+jl1Qd3YKOvMM1F9DZ4eXJsMWC8OSKC9TDb2hlUtkpA3ZMyaCysSiByx9p5Rtqy
SUSqwFs+fey0tccdb8ZtIIXHumfPNuWH08efOfqTi3KecxtJjlQ2+/CMECVXt5mH
be4hlhS7Io5gHRC/bOIJin58YyntTFP3BFfh6TaUraCduTIh0alFBVfQeP5qyG/v
/GF33sufHctxLPF6aWiK3G85La73hP0Q55nC+H8+XnCD/i7P72XiYC7EbEAgrh7P
7GDi5GoSqMtUPcpqKwhqvYp42qEngZybSL6xd0Mtu5yczpylX1aO/N2E0+NbZTH8
mDxrgPr0qTQQig9yV/jDnglTohqenxoNWAOvaA95h7ZBd8dWCQhicvUl1D2nzbme
9AeX6f0HHZXD5HLIeWjWo8ROqBAVAyhLXCHvlKmEMcud9tv0pw9VvtlJrpH9nYam
tcFCVN5tQ8WIAk3sd6nHownqE5CCTDKeWrMIeQHq9u24iCZHg9wbefX34DTDyjrw
ctZJJhKHGI4issYd8MNrM+nOIT1rI3w72twjZoDJMU1k4AL5iogytX5rIACQHdv8
btl89DblGWEExYm/eZT2ubbVbUYzLBNrH7EBs7hC5+1aH3tafRKOjfNfr4Au7kDQ
ERGHmml5jjnNr/Yl58GbSIfcwb4DkucGoSKk9q4IfZH/wpGCL0l/mEqsKX0qEyEG
i/pkKL4Te0uLMWzg9tNXSSvc+m3pkQqQ4tiTnXmVeJyYNJgx8A4hWFM8RFJuIHQF
jmklaDg6dCiE1oaXVgwvuVt/euvuF8ApZo8qcznq2LKjPCJcnv+HM2vFYm4UbcIT
Hz4Xt6/I967fmCo7GTZrHHIorSQiMh6yvYTzDRzJzqaCLnyUxyGL0Y8wQ7AVUbEu
lRc3hXdnn1t50qEESiYCFxd/bJDqkVJ7/e0hdUZnrqShZckogZkmUfCbgdC8M8q0
bNhQ94idwPmYBK/kSTOmOJC+QtLIgzvcRuEeuoP5aHHQ5/jOA0m+q0KTMXgVuHeX
xaO6C3rEs/fADBoECBca9DwzxiQ2glAyglp1XF3YAEYg4IPIdBDoQlhop9EiFTUr
0fOwE/GE8AqxnjKg/Wc4ZY6BLwKxOfi2PQvMU5nj5xYGgY7uARa+GpdJOutGe2fZ
YKpuutH66SPErcaN8tQI7Q5X4pKz/cYfqi0eVW0OR+lweExSBRzGZIumIi5yUHYq
25+txeIGFwi2L41ymJr4mZs9DsFytof5LqKgUOOthjfYbOjiB6ZGvT7HIBDw5tqA
mSLt7eQ4RCBxq1u3WFj/lSE8lCN16fr3VCavTJtwl/VJq7cLtsLIosBZv4z7F6Jp
X6zyLAZkZXlk+G++o0JWX5t+rRSOyFcOm8Zc6+GgeNyDC3JrOmRLZNW8rrLetg5R
5t/uCUOHjgu4/zGwHIPrh7M+wbYbVz+Sl3//cAdhc7TSlKRd4qwBPJILuXjl8S8y
1VQYghXO5wM6cHpVn+Gf+H4qQCZxgMDRTNGGDLXHv5ZIy9ncMKkmBMDne8TmoZcv
s93JlWM5LYO1E/JYuodaHxY8tQTcvzK67yyIwzz63EMPstWuwCddFefbd5JZlxvG
G2vswfoYEL6+o2SWY3DZOC9hbcBXAgTwwmRUbINOvPi9Bei9XpoRwWIakO1cCvRI
isXmIG8Qik0Macdm2uwjXdfXyr30d6HOSWuTOAoyAZ94oiZ7fAcD40OzlwmEuHQl
mUTOQqwmFRs4BWOjJ1rWfDqtHnCEEKQoxabdoXOHth6R8/k2b/a7sMnTWt9mfLFo
3Su6R/o3F3/G6yvzKcHn1HXjsVNG/IB6MCw1zoBMME8wSXo7qUOcmnrS+HMJxGk+
GNgovvnzq45Cr4uj8roowx8E4W70k9uDg3aPHyCYLlaMBQezhs2RI1bPP3MpbU3G
BlrHmGN1+ToW8lRDV3tPhx3JhtYyLVBrLVuXoEsEp/z8EUxpsswvkN358GVyK/6f
SdoY7SttYz/5gDgtOUGMsmOUKp54s9HFqn4aqtKXpTBHjb+0RaFbUMQgB7pY2ABm
8IgSsmBf750hMRlIV7ypfafWSC7FAoJq+cZ31CtHjQ1NmqvROYCI1jr3VomGAyRr
vdmF/pGJKiPacbbeyGWsRU4hx1+KUAgJoD0h6Q7i4hmj79EQ1zYQcyBCbwujQmx4
qLHh1olPwjc22BbjWzN4E2wSvMs0mCA8iYGB7ykY6x9ryUTSPrXo5iuxhePoj0ZG
QfnbAmFk+zKTYbPrI1EtSTb9C9+CyOBQSqlGel3AKrcGlI6DlI5DtxzFwixdwl2C
gRYcJwkTPGaJeLl0dpa/lC/YndEl2FIDPAgG4fHxpv7UOW7fKNsDE//rkMRvszPM
zbsNRbLvJBLJkKSY1v+/yuFGDNIVLPyzYEydO6AFyuUQdfNT631rqJZN7M/3+6mr
hDCZ9Fw8FQqG8D28MStBnsxjIh4sMcD0DZ4auu0PsC9L0NNZ+38y3fQMvwYtokce
SnA/c/gsOUaOey5Dkv1fVj3pMQr8QViajKzFwryfAvI6p0drC1UhbDoCSa6ObVRL
vdukQ7B6NqqeM7q3xKGsMHHacfzTAvwktbhpA2jli4ncXi3BGQ16sfSW4JoX/C0k
ag1RKJ+fA0kVYAgPynF/mXvXc8D8n9BEUdcrdWNqOoPafiKnvaBTggh8tkx+O14i
D+J/lpkmEFi09g8qX+seP22/Cdpbqi7fpOxZsEZQg9a5GLCTgz8FvJAvnF9MfWNl
A8kdcPcTga7MTdoFgDVLmGlPRt/bzVM0qLVE3JRE/kmBtw+jHKUO+zue7eM6bYMM
OUEcK34dYFlyK2zXMPqh2vxfM8KmUDPRfDo0YGObojaHSok1n54UIp684tpuiH50
Rxr9UwR35KNzHb/6ZBuXwdq6Cfly2w+3fshM/7biHDcqWy9vp3FlWqWlRnSpsQac
HOQBGxd76OdWwf61Cu2oetfuLx7I0yyzqtwXBqEsWNmYlKI0SWnlrD0KJaPhEAvh
i5VMSiQRnJ07nL8SX9eZm/RutrmwSgGWe3v7JJ1R96nsHpQxpyk30hOt0spRlNZW
wCf9UTL5SNZtw6otqE30z0fAld6FhvYbK3pdWCVYixStx1LTbnr6UjHpHunQngJ3
IwC8zDX5sMHTqIvxniB9NevHL1OyUdncL3mQLZNVIqgtwpzEgSQJupocI6s2UkIf
gHZHmTS4YT0kw27IlyBfJpZ42lzQkftzrzlD+r1R9t9JMF2Lbz0WZtpP9KsxLikH
prSl/9dLC3N7KyhEgCD2a0JOZFRarcN6kdCoFNkeZsEkZ1iId+tiKi4a8RJeILNJ
Kge9gWFWtNxryMDTNIkx7LTRFEqE/8m7q+1+9fNloER/OulublHY/9DRoE88nvxJ
J1xA8PMW8EZcTszA6v6N1X/Xs76TPTcqbp837aJP9WTYXMChKZ+wnHV37VWRWkhJ
i9on0ofevCLY/izmXwTwcM4c3MHf49HflHzb4qew+2YCUTatrA3mH3QxqwH7goUI
r6QpLOnHIFXB/9uLI7gL3kwR33IsE+lBdDPrSGRWWAjGhLKHHKkh9ymBxACBwH0h
hvDKb2U1sd8O+h5XwjKdkDKboGhMqcdGeATBdstTsJ5Zdh0XvUZ3mL/CO6jEAH8x
fb0bCnrohWpp8ETU50FjAuDWvJVMxhIBpIIbOv/1YHj42W7tcddY+ZcmbDPECooT
rbyB/qEqwHtqDv8r3H6sN9WMr6ulvJtDV7ByPBE5F91D98Fe99LpH/5sWydFJy0B
Lg263wPBrDxmS+wb4dNRq8XjkpznHw3hVJaUm64d4Jsh99gpSQf9jMKCkCUSn0lZ
eeFH+3LpSeoykbendYEgjxelcdusjnzq26vTvx/XlF2sEMHe2T6/j2Ney2ArAIBI
hHo75K+6dqDVinkE4BXcu46RRIVvWl3+oWKpCt+UeCmHbZrokPnSUAOPfKob33b2
zDRz3QkPeEnqF6aAbhZCObei+PT9SzR5o4Ne3jCQafrf9Uk7phPv8iHZ76mHWg8z
Lc6hxxygKQ/cKd0QERM5PN4rmyEJrdfyr3B/lTjVJxe7f19uxjp38TBStfBDaNIq
EjFPvLaS13v6mN/Yh0AWBKgBXB9vlVQxA8mhPAxVCkGN9GFarDqF2aiCky9T2iDu
OAh6ONDMlSY3PLTi81ioshZWrPp1O499obw5mP8mSSYMhJ5lTO+y5zmxEIXPnF4B
wiW+m7jUY2LGFHQPzOq5FeQWGlgl/Qp28591xtSttgM/tbHukkbsMsIxVJQNEj24
YjAC5Utn8F4j3BGvX35FDtnOnjukZflQFSXoERlb71E9TSJOEWoGE2AKyh40KM5x
bmRQ40s8Cel9hRcY+jLi7D4jikMmTTJm3cWApF7MLyB7/rgfE9DqKeiaBumuLWkg
Dctvi++LoYx3hJYGbincK7bfLYAo4zyj3cLwU1xurw+3nKWyJjbDlnsbY/jktiY9
IjV1Zdz6EYToqH0pc7E296b6DoLX/aPkVB56NvCBE1fPi884e1R3U3K4Sx1x4FDJ
Y+ng0EH2yT+lUxD6fhBX/O0gjb6GqSI+0j1zFZpgG7eR3Cswh/hWY7Nrh8Cfj6ye
sYZWujGYt+/bBo5oDoFlwkG6R7qfjWErLrJJT4I1jj/d8mzBOyTfB3NKXAZJ8JTS
k9XfRx2BKidRgcAdZZhkDi5bcPls4qKLB77i0VA9vY7IZjlYSePpE96SQNsM8G0Y
bjG51lctxAKA2om31hJwEFY5qGgmPQg2XmhW+wS9idbhh4XkpfD/1jGBAlqS+XuR
ZFnT04YgJLXJm8Kmoig0qFmwWxXsgB72b9ffOpZvXGK+sfhtgXuV+U9+98Bl7ax0
+ZBUV/BHOFFQRAIZ9SaJPMPt7lvjPIk+TswUp9WCm42D7eVuaQHz1O3+5FOjvSQk
DES9OY4nvjo49rx4blcMZMVfzog581ko5tru2U2K+gTaic0RY3AICAw343CMSli1
/QQzVEbZYnRfc4kT3wkVqXJyoimjsZHkTGLCtg2bg1DgEJvET+QOaBu3ge017Dsd
Tc2bRwJCUWwOj3nICeaM75/ZtiijfoP8+x1ZeOrBblGSZr1oB8P8QzITbxBaT5yx
KCszgEz+icX4Ly6AZMiW4QMXfklWqmQ1LJlfo3m/3VCzwY9cbTm5EUFnNcy3CoxP
nw4uVPjHWXh/ORm4xdi61NPRpLBjHYrOZZlVk1jHP3NkIGx0QX0WqKw6i5CJg4dB
fvQNnn2sWhkAbXouJ+ENvVQ66Yo5Sl17OhNNZN4tQTWlMxDjbHky4wrmCWIT3mGE
u7KuOG1LxfYGT1Z/9FZTJgAYC0JYreMHmDzCpylawKrBQvZOBHiWI2MJOFdRuOc5
jeGdcvuckpsB2sGCT7HdSa4YLRSeTzqQOOOGFKwEAgRvNoC046hwiGSqd/KXz16u
1GLYNzU5ahFaUeK6gNIOkv4d6Y/Wdr0nzQcCDqIYpXMvsbKWQTgDox2SiVNL6gOD
f3uwZpoofxjVfsQ1nylp+zE6AUoOmlbSuFUxZeP2iHFNvJ9zDz1Fe3v60AgdZbHB
wDxNi525LwFhYiDmcfZGc9p/TGKFk6wpgrXA6mNqkak3kBECR6j5jNzTqqEM9sBu
1Kf2XAXtSR0rtRVlLth34vPNrkOxLFsuotpu/KFNpo1wrEP8yhM6XRDS3eamY7He
/MVlRg1crsqty9gYO8i2x0SshVJqO8bDmFDoCKIR0pYfd3UtsV1tCHGIFBR3back
xzMzD4qhAsAhIsSXLL+N0qDjCcj0vPcvN/fOgoMVikjcamuZy9EfachbG5bRGiIX
e+I4TLWEc2/0ycckWMdTUou/qs5EN+jLbXVerlk/nlJV2b2BFhXQP1KiPBeua7co
vz5bJgrwe2V6XZofyt0DOVNtLc0e8BigGJ93Du56R0ZRtAlCaP87KRC+6omqjsu6
lHNo84mfFcPYdT991PVxgoT0Jvz5vJFt38NerRAOM46ryPKV2VEY6KTCc34S+CGh
h0nhQRi7cn+71JuZOlHw55Ec4bokqDeWNXpIAQELvPfpktOROnFjz9wgMId87gHx
Ls6QMMXGma5pkRbdJ7wQtkb/cIKfIGZaCicQsl2kY3wh/dwykiTj9FhFZmCMhd32
0cW0KILhXhkQRDv16QnMjWO271X3B3+9346Pr0wppV2gYh7JuwZ3ImZFil2RDGVL
BpEfmFlRQ+GCeDe9/E1JuAJrSdNGainGaEIQZ18ELFlPxjB4ZEO77osdeTS8VFUn
0Ozkqd6bY8VJmre/ouyMx7Z8KHqf3rlTf9P+oc5zXAH81z2orls6SYvNbsQxFyfn
vagzfYH5zgDbCPKpzHc3Es4J5pbVfnRp2ZM2G5duFbwM9MLdW171WU8pgO6zWzhd
pFyX7kvJSrmH972JllY4UrXCWHK8AKk/5X+1Zeyy5qZ0VEC8dfx7gvfx6MBGd++1
8h35fkndiRNVoodXJHxX7gaSzrqJfH9Z+jfVZS1fUzrOnPnBdfRKvsCaQPjZBbgw
j8xvrmLUav4UwkVDrCBsbUQP/kTt39+i/6aGTyWMfFeAIrdOIYw9Z1OCywVKH3vW
oWU1umw8b1tnjSo/Px5iEMdmHGSez8qxQRJ3lyvk3qEG2bis5m5CEpwbi4IVZ/gC
M9LtU8K9uoiJNpOvT1qSfzLSEdAESLizk4PkRK5QnITZIBN2Mcw0tT1IoFXpgdzf
p0cPPhRGJfNLjelVKRS2LF90H9P9o0xiz3pCgvlBATjRWv/rLVmSgss8TGusp87E
AnLdzbI8sfQjK/f+CCViTus1WJHG9i1R1wxlxjl1TttrQrP0UZ7W7KGjjN94AkDO
puFGf5uCmy9kjdX5r+VI7foHvbLdvlOJT0nYpcNO05qvODd1BZSfH22LzBd7i50v
SP6IdFRHgxSvsboXckKulDaZGFnIBEZwNGSvfuO5I16Uo/Oe2fDi+9yyMeJyV92U
jXT1sPD0jLaUHh44o+0kf66CNOjHwy67qeXfjXST2aZcIDbsy5rp3H8i/iDnHclS
XuYcRP23e/JBTXxsQWQfcaYON8pbWb8pTGKSSQoMrWdIDBwPf5pN7by9uZW0ONHu
RJsUY1fc/Ngv8cxFTeNGv3ePHMsoa1yMRmVeo7O2IzEq5c0LSGaOnAOZp/E8jZxC
1gjd1A0CE1UnyaFbXdTJAoaxOB0CROBvqfFI8D6zcinzj3+4KIua74ZNslNz9nSE
/cLpeGQB00CHD+nUzOnc5nawxBnO4zdwYPvhCeN6ytMHxwPBbTUq2hRFx+f75Y1+
+wxLN1xvCau+bx2YSjObpEvDPrDPlAk6XdwgHU2rG/DFfGCnWbGv9ESxMDXXeNHQ
O5tBFLvHvYNbfgxvvCSyR7AWEoM2GrKTdGM6D/wLBYDC2Np9SXL8cFsUJN8jadZh
jaelcN47jDwF5eCJziFFuYxDWdqjwyNXcIYY2cOh1mxwhn5Efh2wb7PjeiXTyswP
wwiyoGMSTHyws26NDy0jkgq9mvOk6oQ99cdFC4NILWs/6uH1/XuXW9uN2am+XVu5
uoAhV8Dvqsk8MZ768UsmkzObQ+VGaefk5gkcO8yySIwYUWxkmLQl+FtB4LYsPmWT
Tt+XNboSVTHD8/KZiZhhhFF2hs/xT4HJGqKXht0AqmTFU5hLe0yScRR3RhS6SuHF
LywnCpCVN2d7k+TAPYae+4QKWTQwcNcdX+6a6Qsjty0akZnw9c6oprnDJHBO4n3j
sKQoRNgHrA3ke4KS64+TvriIzekeTLYa/jhRAk43UM7DDoJso9vZNrIkGOg0iwC+
QvYvIq1xCgFTJVlcQaTgpApBRvcvE1t7T6zmU4862mj3L7Ga17Jn4Op5KsPJhNnr
y2jXMUFy1dOzPmNQITgrZs7XyovyWodxmeLtbO2/up3CUOfd8SDxAsip8/0ILmw+
ffHNVxufkBbS2qFB4cYAcr6RPrTcDgfU25m94Y3K8tauXRel7L0U1MTx+IP9o6o+
j6YfEvdt5h1VQXinKpOgrMh+xUXECtSeL0PTL1KjjUjV49itIMKjoy3v9Jq8joTd
5Wzz/slWJPbwKIk0b+QThAfBe7ydcyRkTE5dPB3BjYqvjd4Ta7S/QE7N/qv7UdAi
+P9qMvpuZKu9P3LXDEog7Zj74TOVZTQFgtS7Np8ROGqmSz+9DYyRIhQrp1YGML1r
44fPWo61lPANl0e9aLbcVG9S3VmiZnMb/HWCV3kltwExui3WkCFDUn1uwjyvEvR0
CLtVvtNsiSmCX751ItyaR1SYRvzSkkRpc8ZCGJCi3FDjYefGdBdEmbPsfM3SUzlg
Q4BOMdMv667MvvRS8hRIH9C3NueuJvWHDzfS94kXxBBfMIC7x3FHDo5ebnqqVsej
HW3gXcD0TJYsZvNzlkMAod2CryNdHzEobUyV8ZzK0w+96g6JntSrokOU/QXq7qKB
eReLZXe6dnrqdrZtuAxZ2j3839vtxE10oHthQ3lUR/qHfvEh7Z9V/cRb/JLT5ILU
b5blPmX6Av56RFQK3S93AeMkCWMHSvI13OlTs9AM8cgfABGXgkje907HedTsdlI8
4fvxjrSDVMn2kn2ydzCx1N1EuhjCJBfRaXfHQgenoQNahjR7ni/fNULApGj3BpIh
MerXKHDnCWpPCoq3tCdU19vX3j52oLAdZOMpgPH5drRZmvbrY1pP9rdQgKBXUfmU
zBrdm2L4KGWZwJ1BI49QfH3nwUfBZy0Zu1m9SnZCJP63JA4GQ2sdX1knHdYImsD+
Av281DgljXzi/D4pa9kvx/Jvy8CN7fyFhwiOD5lA/p8whPo4ZjlyGelMs659Vgku
pu2RztbmfUiAgDytlrAOVVOAHv5my4x1eExHnvLYAJ+dLRLEEFJ5W8aB7VaD0o4Q
ECH15SIzrtUucV+S3hI6NSOtw23aYlceApH01j+19m0XPUtvKIF3RyV6O67VZ/ZZ
MwazcuZq/0q6+vJyTD4abKOb5SrtPnd8V96qd3HC6e8eLqSrp8Uf6gp4qvHd17OI
iSjhKJGOvN1byQwGnP14XzsnXxqzpn922E7FF3olRkie2qw4mAGwuRo5o3QaBTky
qKfbHyECnjYXlxf89BSi/teAo+aGjpYzuExdl1t4Qts8Tp9WgIDde6ziB8siHV2q
YuvIPC1Qo0gPrX6HSqyVxzRWHwtMUd8hZBcWgpMPzdrbBh+QqUeLS3revYmS2qhe
da6ZMO3UH14pgk5ScPqk9MbNsNS3jueaQL2bnbhbgBz+dXjB/s9bUw3warloRd2Z
ouX+D62UiIM61mQUiqkAVXu4+A2WV7danYKA4iPqNSoHAdYS1nP5xgzOA3gyzRVp
+yoM3FSAimQfY9Lyx1m7lsu8m53VNiysrm064GOjrNp2QtH8PwazMH/cJ0Fk3ZDz
2TvcuwV1ehzDMHbweLQC1Ysqgj+H+2npFRsHEl69rQrZhtzF8Tnl30lu8Vbm+ttH
A7L53b6J1nzAeA2YFJrA8arX/OtRVPgUbre91pJulT3zsgq+ulPfNqUkHxkChOeu
ES+UQDYvFUFdXWTibcrIHm4Bv1YjVOwgp34dvMkFcRO634Oj7fhO5ebmm/wRHdVF
sTaBitB0NjvJxlT+A/xU1tvhMMxvnAFiuva8M3qj2ZjnP3QTwok6e2Be6I4BwA7g
R6ySm/DHvMvnqmVPlREgxuFzQ8HY01uuUWh4vL5u+pugWUgUzrWXlz4M1YvZq2Wx
G96oOuIEXZ42GNhaJ75B5Om6xhrK4e3ROhh8d9l2f70elzucBZ4XirqbKmwcloxW
8YloXQdB8/aL9/ZBWHy8a3yhH6u0CXt/8gVEns+N0rNsabaLxequA3jM+bg7NZze
jb5o5C39S6QhMF67/uMFEwx13zUq5I5bbUbH9KBFSeO0lho9LHpeJJMBfiOUi6ao
5iH62EF90YwD+uWPa0MM0uSyxdsrFfv5AGcd7VbArcABlYCL8VZk8CcNycj9MXFW
J0WDOD7dLd5AnSxMQ0q3HC59tZy6QBtnb/1XWbBeKjCBvgEIfDHBQGlj7JZNqgsy
4c2CldPtfjogH97x09e4aEpeFEgdVJDDhk8V8Gl3MCJawXYIBSwiGmCA2V1Ouypy
oZ6O8WfOo604LRrGsjuheJlLcq2mbDEZLCCLUp5hGCYIkirolzR1F3zrljA9RYfC
Of8z4U/PCi1E0b+E+NDbe9Y1zijW0XSQ4QSleeEJdn3+aPwn0debGDGsyR+k9UCq
HpS0pJoJARxsrYyNS4w84pwxW/XUGkf5QEfrw+wTmJDGtX6/7jnyAvt84AjnI+1n
jFpEKhHi9mRjmr3mt74p2NUVnX28SXpz9A/x/QkeljANpu7y+k4wFaoMCsqLLeHV
pICRZQW+gMLvFspUcx7Hk2Ib8WyRxtCHqljvhU0/nRswmvaHuRqPiLjdJ9z5eZIM
7Kd68uJw37lOOE3Yayo1wYHy8kIJhj4JxXXMuqSrolVsCFDCi2NipH3nfkGPwm60
izG6/h4Qz2KdmSitGbAdGsli38h2RdlDWWDIifNvE/dsFDqtk9PSIqWfsDswLz0Z
mfGVl4VrChYEkGp7W6E2vL9vksvjryNQQ8cEjBFDtMRuAnxBSxzNp56UViGXAIdF
pBCij3AlzogsUjPca1mWghsEhg/irA0NdnIJ32U/e40mJo/pl1npWr1wcKlDj9df
rz58X/RkaU4qfeZQg5ZkSFswMECKXAYnuwmoifBxE5tw7teIaUYKE6lYwL+pzGY5
dBttQw8WI79gpOeYdgMqsa8rYV49ALMdmoG98nGaEGogVeRTLxuZKkrKJPhFGYUF
gUk9ozG+GZTl3gFjEF3HsbuR2Gje4DadVgebnD/HMLFovueXYMuGD2sQxm6SOEe3
RKZ5RAG7IcP680q7m1hunhoT2cZvL6yupGCIUolEtbwqEc0pRdRCs9bKXNrn2ePC
+aSKE21y9IfMVeL4XFbK2G1h4Rm8i+WNsLHj3W80r/HMenfAl9AV2zkzHouqZAwc
wpEIbAtBfQYu0sv1G+pnCxaqVeC/1SYTuhTP+n1hIyLL+muTQjWYWbS6UdQmEoEe
q3BnxfjSxq7f1Ln6RdIf7bBN5OIJWxjPMqmnKL2sdhLRLNiCiyCVGWQOdyOhclvh
MUkAgGYjFS0XieWCk4++XrSVBCK8ZgQTIVHD/cN+xti5SBw5WDJlMKB/KzUMPgUm
j1gNHAk2R5bj6Zlsc86hgqDC5QVxHtyAdkJT6nYo0hyarpi5dQG4TRbwkB4RckVq
fwQpDeckpV3q3/U0KzKex9a5BUMejPyBtiWvQXwmUHxd7RAvLmm8p9wjBamhbXLF
jSuFdC4gSHRcNXTWxXDQXLKAsQb9x94am3SFSubCOEzgAQFo2CXOEjspmUTprNHp
vWip1s3upF6RdYXzT2B7dJjdArJVlP4RVA0TzHhMkb5kx81AZfxgDxDK7458UVEa
uVvoOGtbsJYhyTBKZD+XYmWUrHRVoqI9wzQBwgIrtD/D9Z0MS5YOGEPLoMXP9a7h
i2Z6fjpPbdMwJFjKjdIt0QvBnDGG0/nkuXjrCcAnt5PctHttTEKNLzJikeELQy7I
LUWJqqmKyDqSlyuk3BimABAo7Eb9CpmU864nu/HmxfxAge/4iInWudMfFW+jdsDb
tyT5mJeSqwclpVUO5A3tIu8tkc4vLVs4D6XYe6GCY20zwswreod0oMS/aEYyVXIN
cUadCEPcHhWqsSnbVuwPgKMBKCIkUL1NN/L5oYeMA3yVxMKJ3kbjROFph5r0f/we
1Bscl3FPe76E329JjVj2hWfQnp+2buwD+U++pU7Tsy3WJy1E3T6dqCAf7JHkkEBv
I3V7PO/PmAqWtUN6TlRvOriswgGPPJSihB0rG1Usi0PsrEAu/66VYvVwixFpDTUa
+8V35tdIYol2vHQnvhbIPDS2JWTJgwhVQUwKqhAwsRqp1Lma7DZctw0MNdkTRcGs
mzCeqCugOKjY8WP3yF4y9hRlA1g+qEjiroNPt0+d09ThP+reDKJvEpVEAJhV2k3V
8oxroDxycihcdlQvAY22akf7FE717ruG5S7WZFs8opsxxTx7/MK6q09xE+uSk9Ev
NaQJB6+y0ILm4rX+10fnJ06gKRhtZClV1botuMbdqObG+X1uOJujPZunE8RQKUFn
3y9SkYt6tt7yirT/ZycZM5XLSkgZ+ia9+yqDlpfCEmlJEyxxO1wemuz89i5SE6hc
qhMH+OIeWH+jCyPfA+4yxvLWZR35eZQBBBW6w12aRvjelXtZuOxW95TfBvCQl3qm
9T9o0AqW9tz1y0W7abeGAiC/grJEK5ZSH4YjpFWAXPPBhBaasLBGsPHU1LaWJbtu
qa6HnPWJ5Au5N2DjXhmM1aOZazsZ9MmBtwWoYHj1b9guC/6r67pxD0Cs7/xTNEtQ
TeeQTPEM354SUzYNENSV1XC+TmISm6LCvwPXn3xYyeee/xmg96KNWjV2/VEx+dn/
8sZIAaX1uUNX6bswMHLo/W+wgBNRaDpCh+yrldPq7rs4xs7sf673qePqwn6MViIX
RBS8T96nCFwffBMBOicavh/Q/VE00XpUiafw7EtXoYv2wYpleq/7b+YJPV+BYeYZ
rl95c0gEsNAOlE+x+Zs8tFkrlnuY7t4Vp/dVktPvC0fwBwHh70CNqkkjEj/OJCW3
cd14QaxNwgSM3Fsq4hQ52L9KdR/G0NaDL8D2k+x8BhK4YyrOjLZNXS0n3czPkBge
/Z9yXYRCgqJIZlu1Nk+SLqT19pV1CPQQfpfu+gQWkKsgPpZxLnJECGI/f/nyIkjC
SKcU40tYtNJHrIdJzxqjSjh5nrys3DVRJtIDKbPIOWW62uI9wss5nnom4IQJUDEp
L1HSUSPoLw/NFF/QPb2svPucABbR2pXwmxWzVV1VnGS/Cvqjj2cM4LsxdPq7RZKQ
1Kl2A3UdTA4euJF/LdaJge+HNo50+hmxrznrvIO/Ng5bjtylPVXqS3IkWXbzKQsI
bNtmnY+cCdl0Qqen7O/kmbeL4ZrOVHFlVdj5XdeHJxtGLlyAHkglOAAOFAwGzLpG
ADxRmObPn9LR06yrOWJIk/lz5KGqoU4CggMcKOIzbGbmnxE3TuHylQ3XK/d7N1fr
xB3aJO20jtTPlh7u5R9zSywh6X90nI9O3Y8du0oi+PBm14jKbdLLNSS6nvk/AegH
evMNxRf3x3ZAjN+rwZGACmCpc7fumjiMp70l035fmQB8GHg7CZ/lnYzWdVAw12Po
9hEkdp8iOEZxJhoTvM+awSFOQiNZH32sk/qVjzV1LptGCy7dM/GvdJGcWyXrhrkW
1eAB6AuPZuYg81vBW0pjAp98ZjQEIt/PRkUsqKHk/BX/E6Rar58S04RU9ty3fhP6
W9Tuwdyc/ZCcbidFLJDx28a3OrOWoBl5vurYeH63V2mMP550qVwbGyUY6gI6JLxl
wL/NrC13RCprhNNKLztQDAfMf8Q8mVDZakTANUDy2Pt9/gLFFanOk2ttx8mupudC
6t4+UP2jBCtC6iKJpc/4Q2M/wPD7sNHIVMcLM9+F4FGwl3y+D3NF+4VnbMv0jjC7
KXu1IdO1nDrf5C1YZmsFvtw8myQarHd8J4QHYrhfekkCQK8t5hkhLVtmQTKUK3oT
0DmnrnDI4+usEwOBATku0sdXjudBseP3s6drSVoRjkNfj09EOk2zEvJuLlOyf8iN
FEYcLem6owwTO60ey9DYAHAmgQjVP2/JIONd04rX7lqhbb7Wk06NJ2jomr1VNbWA
EmWtbRb1c1GvT5S1dPkbZryM0WQY1sNK0aU0p/R2xpBnOloefSvomcuVW/Fs2HOk
hvFuJmXYqoo9YsYtDNfsNXqA1Br6lFyOkYzijYU0nWXN101Qm9IwAKjpp+oLEgY4
Jkcg/CHlW+SPoBMqceB98sDH+yfNyvRN/Ikwatk9b6Yn2YmQiStRms22SKV7/dX8
N7Z3Oos/pNRdmDqrvwZ58xUS8FzXDmYE0k5MmlOUY558FOMmu67L4cJ5dUSYOvO5
PGE+izEcGl+gl2RWL25iXnuXa4RZ1IVUWDqdKQtqgXSd66guQZlGJGuAet1TQ9nP
yTy4E6N5TrP+fSQtGMByNuKELlBBg8D2HntgJZdkclyRbxU27hKiSSBtnz0LR40P
UWXl/kZF/UBh0M/pY7uF2aMU5bpYVD+ptMEuLHQH7IoZMWT1dFLrf88cCxQTzx3R
Y+jtzuIXob75J6bHhdhpYBunCyk7FiFDhlESieFwyJG6b8cjhGB3F7yiOuH5CJXu
dcMY3eJ9SCRYhsF6sy12GdiLy85s1aB2nOYTo+//+I1abX8NO3xNEIUpOhJjMvBO
fCq8cF2QdzfLVM2ZXGgJ2idEZdCa/C2+cuDLdpokpoMXwcQsWRh7JyjrQoG3tkAn
r8cjpYQ/EFiHP8n+vLf9M1WXfkeVag9PVs34jOlmUu9ZIE3dpx1dc4EfO2n4RaHw
scDSMWhtcKqyaNonM7HqMfP7ezso6oE+kIjL9VIkZVTLqf1iDfn0aJYgv2IJ6yRv
p0Hna88miX99ZtA5pnMyydDs06Eix/y9dCmURUhbmQ4MMC2A6L0ue+ezJVwZJN5m
1f+Az7Mlsp+exfKm/acDZZGztfHGlh1vHF2U/oYLkh0Wj5nAqu4avU1ZX9BYfqOz
yXZdDPBR/vd7BSBIM9hjFjcBm5K8TGA/Hk986vn+6qhuHEKO7yNvj+J2zynHwBTv
aled9daDzG2C9F6yORYGWhMQJ4n/IqoiqHEObSMjZxaSdlig97bxukfD9XPY6/07
76MxOk7rL5SxX+INtubc+lbxfCUDsK0NDCg8Mn8qYC2jzczWyhAaa7zRGaypWlBr
SLjbq/58xXbWBZxgnc7XyaX5ynZ+fjBEsmfA7/mw0NiwvEg+BpuMld4AGqNBf76t
JRkmCtlJ8zOw2gayCyt2C59y8bX4iBR2FoOE9y5SoqvoLG5Wc/Us5JErpAljoZ0Q
MkC6zIK10STJlR/DAHhTfnkxBYNJm7V4UJpjEayZhKma4WcfX+AnxWI2ID8a8Jzp
nySnOEt9K+tKOxFwrthjo2At2Otl2IMj9KtcX1NNqXeVLbXzWWQHzujao9ReLQf7
kQb8XE5Z5FxlSs6VZYunWBaVtAEUWbiTRW+wyBONe1Ib9NR4lVdofTpI/z5rfeW/
K7+2QN61cFqh7DI9zNvwNvACVqWf/4cv+cLBVi5C8hwapreU0IGX81VLgDcaXvZx
FQ7alRwh5aVYQ1XvdKTat6srQZHWd4+UTMLmqU3fbhwgMO8EpIqGA1zUmrikBEyY
mOkymxPiyhn51aXjzbLIFgOcWVa2gfOK8dpcg4l1huT72LpB5dG734nmliHhsplX
IkkUBMCbpsxNnvY1U1H+dpt+8d+46qXy/wcUHMo0PLRksZKGAPUuYDJ19oIjMT/w
BdaKuCR0QUqy8NKqAv9b1v/bI/SnS9qd1F5aTOzMgLFFLXVmoX669mFy7lqTSA6Q
tY6gz3QvaYIvyEGcrVyX6xpT29/uRbxhEqYf3/MtKEY3jq4n6ADaeG+xwlod4aFu
/twJBy9A59Q3J1qcOL1necpi45n25B76Mq1iTCNlNdMk+4NRtWI38iexpE6hTnUQ
R2uuv6BtLc1ULAqvUgQKBtkgfBzF6C62Sl8y6HItNxVY2Fk/d6W5WES/mOKGT1x3
p8/Uxj8u4kFaJesuO2jLSXzEFCanzMeIQcBKx/92LiRt+3rwJZk2qRluwHe6FIj7
IfwebCf/AMXrVgYzbcwdd9ZF/eSChkrebTH9PqGEVOsJwoc9v4tx/vWbauBtWCQY
b3F1997/jXG8uEX6RrYJ+etDbPwMk3b22mHjRfjgEzXr/e8vWjr6BDXfm9PjHPU7
QUKdLQHT8NoHsFQyJnAOZ5jEjKYxzKxzJ/A5WVZcW+PfjtF+NCAMkTonBP2q7A7a
uA+v10RR64r5lcnZdvpsYMA3OYDiq7c5Y6JqrZEa1t1uxvOAS8I+2VuULP4xp4OG
YZHoxWoHnexSeGPMYA7WvBjWWLUGJYyxq3wB+ImrduaO//vTDHcoXO6dZfL6mygi
5HkQUaKCaLJ5UfEsvrpH86W47CVVjFTUWWhj7XIJJUPmoHe73K8T8qZR8pwusJ7d
WG/3JG3u1KFHBRr9/sSi+1Q8GQWgdAnPXgVjJMcm9vPaO6/+ci6dfHFz0Rg//Gze
W7Wst7L0S7Pe+Au0VHCMNvOLqfYimSsr3crIxoFCFT4Rx8HDliNznPXBlOLxqnNZ
I64wn6Nmtcv+N8LYOCwm3FTY28Q2wUlK4oKvCC77zlQVi7qLVOjv0XhqTHqXWfeP
1XXawqBlFOyMveY310vIZpiQmBL4BkdFDrQCofIFQy0LahD1TeDxllQOMSskN2uq
JRQoy2iOc/H5OdiOEBbw7k2Mo9hkhtQyCTLiqOP1g/rKWdmyWYwAsk6gD8ms3x63
s6pAU4uT9kjOL/I4yF4v6heYU2sGhLqCL3WHhEVm2Ty/J/PfbP6rJMd9COocx4K9
Phn9Nl/EuT09XkCu6sR7dnlyC9+7e8vZxzFhXKxou2xdNL0+O80Kt6Va/C/1bq7A
qsci8bV+7aNGYUfUb3Ahkmy3vX578BocCYelwCbUBsGBAUjxwCYidj34CYba2OPI
Utiar+yyAesBxw0rimu5E/ce+5oBeJzc6BmV7xAcdZB6FZCN3w5taqrIkVIJb/hM
Uvb/2+JwPOGT6jjsRxfhSNvdOxMWT1wN9bSXxYEs+PB+GMgP6dFAyGc7N21+rANI
3IdZlVqA0ywNwt8gDHlELV8RrF93TAmZSWGZc0bbexWn0kaDa6qUhBkRAMgq53R/
p1lXg5Iy0PEwJXRGVdldz0BPzmC66hufnif0xtUyRR1hfX/fGcG8y/2x1m7o3PJz
7GVByK8C6UOFeBNCK681q81VSuHs6hTR6JCJOsjEng3C3zfOpwPKbQx9MlbTesEY
D6id6S3I84M67UPRIBBxjNHxMomwNW4o6y/YUWks6nMuohuzPpi8twnuxIVjoUAF
TuJO7EXPvROpFvPDAcRcWm93l8aYVWhn5n31/p31ZyI16InknVNtpMyyI3of5Y2U
fR2E4usMh4CQxGLd/nx9/gVhQ/j3fAb0D5NAcWsHB2pPzdQSLBy++6/9L7l235pi
d50QTkwEMtrT06en0clyXwP2AcxEfgmtbLAnacpylmCNBb5TxGeO0tqZvTTDs2UL
G9h2KtkBoSslBOZ03V1HDdkemVGLGWi9Gudtbj51WJsm2u9FqoWLYGz1R8e5ZD+W
SDGaLS/qKCwefBiFxhYi81ppwjm883LATnZiVMY3FgjJhx43yTLL39wT4wSIh3Ee
W8grZS+kAznx+6IQ+InC79e/hUKpGFgb/0YEIJJaYVnIJmS95HtVwo+6pPsAU12E
LKGaK6/BIS6mxUCu11/wSy1QIGhMLwdJS7IUr4bg/Mq4ndiiBoN1QHoPZ6TdD1fc
PEoVtctM6fF0wt+sX4OaSdgLrTBP7VA9oUqknuoqqbyjhvtPCiw4On6FgQ50YkV9
xEwPh+qsckpb/VxJZIL418/ehkLUDbHleeYFtXRWJDZ5ViOkaeYdVMBt/Fafz7/7
VZsYmMqHcOlg50kD/0qjsQ==
`protect end_protected