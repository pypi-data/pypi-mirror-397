`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
Hm0rc5KfjNwPmEU/4qyz3X5GLDpFoQY/CHbAFPd7KKaTg9BwlZoohH4KzvFKmLaO
xM2rsphB6j489gjQ/YpbNJe2qpMHv0pf2zdLMvloPSrgTh1ik2Wnw+aKtRhKYnSV
fhcdKptIdlxDvuOZ2BiebWx3BplyxGnlkzexcDW9sV2259MOQKw7LYUekTzp2xiR
5tAa2LItepAcAQdq95NMO+wtoPPVKZ+hMyOfo5K0RxCwRun1Y/wqR6ASBSjT1Tje
hijaZHkkJ6k6YjqWlJ+XJxPwWq8gzTWqtRH+ynGZ0oR6EmBfAKf1jIU1jU5bvepN
nmPRYFKlojvKgJM2Ws0hjW9ulH1KQziStmqzx33rgZRFPeu+lEk5ndKSYQxW7Rjc
VaCwOXqJaHRM6+W6DmTVTUJP8V5lf7qkJgNPpBO5GDGSmAfiTHf9h44bxtKtNd1j
EDrOqypbMeTTz8bj7tQ4+PcYsb5sAjcETJrlh7blfBBYJsPhpJomxiztjs7oTfFX
eke4E4XVKXBdyR0ZMif74UnVXtO+qu4pYArCmI1n3IDU2/xowROjJVFZbR+7poMI
diDPAAlBxOJjpEj+rEzmVZ3YEaWbUqXykRpiXv8+5tBG0YSNNJe/yuj4Aer1Ovjh
62XlAKEcMOk4Q1ihxjShOKFuk2FqcxJWWH3+mpmHMYeA2bPqFyz01RS1trM/syXi
4DevGVbWwzAhX8Wdmj8tdwuJeMxoJ3iy1VGsdFuyR1Q2gs/df4olKE8ROFwv35nz
f1Ad3Mrr8uyvO/7xLcbYIrOTTwwqwwckdbyMOBswIfUYZHayCGxIrFzZv+kDssRk
9tpKZ3i7GrzxG9HdiacoioVnKR24rPtiC+nGVTpxCWiyPSL4f0u+DdwNEgc4/0ud
zjRfzRg2hLcCpAWTvMNzcevHwNpUHHdNawayImfw684VmHBwy3rZONOzuEXVrTNy
1s/CfXnv8aw3MHpAdECb5bUku1vE8Fgl2KfTfZ6VTDsROQYlUGa2tBAsu7qGmiMl
SGmNX65OceHi5Wl6O4imjinbQKE0K1/dUQ5bkuLtX0LlFrkYP7wVrcPVPaa6R6rK
h/iFQqTy0SAJKVLEdAYQXTG1bL2R9B5aRcPfgsXeLy6qa7iYszFalsCY13gYyAWr
FYI9h3U0xv6ermjRk4NLgVLzRWk4Voy4+NSuaKoutDnEqmNi7vHuuvGIrjWryuiV
rQDU6ehDfXXHZe8tfMEw79V/CnDXy3ft/OFZfWVGWq+aj7v8IgpcclGs/cYKszgP
DcYg4v/jiAfQboZSL5gzrvG5FwEknVPeF94KmIoA3iI6URhZIMFhX41As6icSb1s
hVug0iDwdqxu9biTYfcwdAW2be+5XpAEUEXtXMRhEAxvWnfRP9F5vIgdGDwY4VzA
sRo92l3CDtW6DToSrhIjvIovUtSL2o95HWgbGicQiZti6aRoXrhwEgf8JUSgKGic
Cbs9Im7tGZC7qOk7hSgfxDuF9D956kZkcLaxOsTGAo/CdNzF8V1rCso+cDXvHcDt
3M/mkw4xtQdOHJoAblTwxq59zYAT/88CgvUfn5uppxjB2Ckb4rrUtilkRDcwUHWk
GdIkMwJ/H3PfYPjQrU2uJUttQzBWtzRSogrd4gibNhpL3Og7Va8GAJohuyBWQAI3
UCCRnEWJz5xbiUz8M54RHkUFVZKoi5SjbCUsG7FcolmpJ5XoJNJFnEnEXJvKQCRX
6LMGCPc0qFxgI7s4FkmQQ1U9FpE+MsuFN4fWgygwIJQ74BS5xte7252EHHK8uslq
71/infsNtI9nwSHsE6g9A0+e3r7lJuTCc8XKPeHy9yK4iuJLyY5WVOU+UmoendW+
UR+LQ7wp6hR/RGMkSebYDeSZcd/j7JQcqk3N/G2pNxjPH8CWcZqiObFBkrgTpyrm
jy0ZNWzbwLQpYjBVjNdmFcuVoEUH1vYO1wz5tZxfFKnf4rSCJadOC1CcDchFEPv7
ty1AkdL2821Ip9rtKXv/oamLl6Lj3puEn2idL6IjSM08Wop79AV0WTbwXEgUTR6o
a2aGKG4URksY6w0O99ansRbILMIg/ZeQeWK/WHPA+YbzuTjTU1894NVDL5zAsEK1
dev4yO5bNe1YLHMx9w7utCk+1A5xZXIzYrBLXMQwg/wWcWA7EhwdYswbZFeNJwW3
KW0zySYQ3NPvKMzl7LorR911lIkuuNVQSES65bmPCSgljGcn96YFZoSUDXvl8Msx
Q0iWKEcwnDwLY2UAkimNdQXm+YEq3uS95N26vQ2bnpG9/mMkfsIoHA4cl1/t/Hbz
aSovuMAFAvwwugLtfgt1cclY/SiwYPlBosidE8AaCuCaUt471wQiBBvxJpWqLwt/
OPnr4CSPG69IiNyKBspVV1mbg0KxFBASoDQGzxi+gGpYx7Gxnror/286kbLFk2tz
BPLRKe7ndVW/HT6C3vj/LX4Q4UCRYg/j224a94XFG3+eDMXFYsQ8YY6bCkdkiQNn
mE5zx3ZC4oztIWPcQ2QBlZDZsD2K8objzugEisu46YDMIFXUQQ5Ws5+XEqvyIUds
`protect end_protected