`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH6eYGTY8O3gkWfaoxhCs5Pqjt/CefBVmM5Wd1BJohl7+
2trCmC+8IZbsERcZukLN3IDyXu1z1Ivao01ddSIDc4TWqoEC0oCC1Ic71R8Yio0j
aTONC004HjHzGJa0Xbpsqj6Iy7MfVUUHnVHRS8MOvLJO/4r8MShk8SZSCNReeLIZ
eHhcGiZxi91sPPYPaVHGshhH3vNAt//tgv/0i8h5ixgloTtTKFdpL6c3HzNfRCUN
1tOU7fgAKtB55MtAaTDxDT/hopBhChJnPbx07D0qsLKmLm9s9TcsVMrW/QzaJg0v
d/MyNYkvIKQBqX0ixRaKXKZM1ZM00vkF59yxBpZ+4HtrpWBRP3ZiYcxAjEgeF9yq
RMwN5qlgbLVrfV1gasbNOu6Hc+0ociRTz2claKjO6unFgTqGeJ9yKou7VdyJFwFd
YCfkgG7WcFtIW7uWxv0NgrMUokFVlRDtQxOUoUCZDjceEpTKvyLwfLaK0fVrGfrZ
fBTn6GSfqeZ6Opsp2FWUtiVKrnjtelznuho3KmTmw71eBL4+wlyrOYOjfY5NcKxQ
PJkaDjwIL70UVoiDjlGHmTWNh3kG8LHP8yf8WHPGPt0PDOZU4ONpYx/LAE1wsy5J
+HJ4zyIREthb4OSTgp/97eVyZtzMpNOvv40GzIromTCCnEedw70CZ9oICnDW0ZX8
m0muJBNKY0vEuhOC7mabQ7UPievQkFrSrw0mafWs1DfhBf+WranQHp5Or/7dpyj5
uWrtKKfvcJJr853Ylv73W6Rfz6H1+ESwQivUoH/Rq/HILrl0wartmLU2UdEArS0D
L/DgmEcBBxvxZzDyP1x2pGEGW3IjX039Ht+WE76XxgKxnuCwTyx8f4jtRPX9YlR/
jhcmyDhdiFhUECGsK+yJKMKXRMaE/nTlO8/YOise2NYBoUJ/+yJ/M39SVEv1ie8y
MBCMLSnCXJBzIZNaddagZTeAwexkjPz+VjZz1BYgTTXKlNDuvA3x4Q8fzzPy/k4M
6DjmDHs05/ujN9qemRCUFs2VWvoHH1hzSo+J6Lv+ali1J+Uphz0rYqORNlALnrgD
WaFPeFF549uIrGbB/ww9vHCET4lAhNHFB8EnYoXgE9LHagkZY8ikmlg42HiRxV4N
Oo9VJIgylC5sD5JrMgDfO3zhDeHbOIlH08ZU5t0nMjXCGlB6kiPN3JTeBHeksLUH
SoTbpTiSM1WML1wrNrsdF1tiqOpM32t8S5lWadriodqZpOTmJ08zsqL+JxCRKxpd
yCw4DhnLftVUtEXubIH48oopcJ2vP45r5S873Ii27bV/plbn42cbxqk72lbkbAvv
aq9Sa1jYzxZTfyFxoBYDevSUjjVilwIQbGbGP+QOLoP3bCuc1Jq3qgzBVM2qPK5V
LB5LS1EfMkc6xTh00qDkSdJN3EUUMPjg51PjhT79DiPaJJwvHWfEi+tyeQ16gssJ
HddHhcoHjajD5zLlEAOKr98Aet/TNNsbrixLXi++x8azm6LeqvENVeQyw8AevILy
Z7T5r5uishj4MH4ggdXZcfVk6IRU5YXudH2GYK6Ug1cJNhXjJanuqCR0LKD3h7Bg
cG2iw/V7u8Dt9TxbHCiv6C+NNIJdM6N++i75aXWtUG6llUemMe3VC8IGtvnfmXvW
ZAB5VgTLVyQNlGg8yzYvYgRQ6RULAmjxzu8cOa2uJ1iNXOJy++suHGvLVRVc9VLa
eYEvmDFIXUH0flwjvT7HO/H0t2V8+yKih5BsafGtCh/E6FDHqqDLq0xtQph1Wmtv
6XkQnB8i101UwIOaU0iBVogAmBet4x8adYJ8LRCNbREzKLaOA9891pwuHSkFYETq
YNBkVSduaPx9pxPeekLOvZ5v9V51+MZeXmfYBUCrb6EIwQCFSD+87TWy7+il0wXy
MKPau/gIJ9v26RkJYzAq2rysk0+Gn3SgKoOwTi8hWUo/jOjgNVL7GudmflGwdHkH
UNctstA+Mb7CR1p/b/7O4ddvbUZe/kbyZPgsOcKxreAcRnykaawna3Lhl6uQuRDD
DjagCC0YkoCSW1qyP7dOU6ytKPY0YRxjTebQkV8o6CipcjZW4IYSnswzJwIU/24c
8ERJiqNBkEbm33nMZj/uGX4TXNmFxPoOjm0dlAJRTzfukcQUPQPPaf8Gbrneyhta
C7tiJKd3tY0BrUV26fLIQuNHVfp3mkEp3XDbLDVmor7g+Nf5P5wMPa7mJQ8umQXJ
DAJJgwBHQ0PKfDfT31MQFn0TrS+mZa+PrMS2JBDv6tYkLvgnbeMvrm908ayhDgcb
zzz+Tl4FOKBuVp/2afm266LcGkNy9lFPd5DL/0unsPJkicFHqmFLUzwi7Ff1zHqS
o945/ovWzC8THpRFTkDRiK5v362XKlrofaivZzDo9P0ssba77tRMxsn8nGWW4izo
yQ/ZWWBVd/ixPGr8muYlIhH6kLrXwYrrWjqDZjQr/Df+5D58DKtUvMyze8Lqtc4Q
OAsX0uA/G9xCcdK5g1Qyt3Pt0Ucvs4rt9FfWR5x8iKsvZHUvcLCIylX5HOxx/sNw
Q/yqmOErilrICyJZZ/8KDXXxiJc2TwAIO7sJMWY5xet+4bOXH1LAa39sH86IJhre
o1NQnlWiR7mMvcM5F0lS2+GdF4PWZH3ERgWKT7DDbLjS8bGQO9Z6uzVTTg8Mu3l7
XB36NaGGkw2p8mVKLsNlsUQirwaelC4hb8eDWqiFW8GqhoHD5ieL9GYv/QWfOQm3
PHtToPy+lF/L7gszb/eY/+I0MFGEGeyKKvHoPhxRXfbalmO70rz5EmRx60SmVNZb
jD3FrEyxtNHNZgnY6E3sfeMW9BvwBnlzIXVtQHo7sWmO0y2R/0SukaeC9IqLa54D
qHNcjwQvt5bzrRmO3kcmhJLInaqGHo92kG3Vdwte54gHjPEtCitUI/dXSVL94PyA
69iBTEQx6OZXWRCl9UQTp1dqA/EgLlzPbeLpUoe6sZqtJ92KTzeGjLSqy/VFZkjY
EcomdukrUFw7r9wHBybtFRJkb0MZBJBH0D421U1ocJ64+tzREyMt6i67uZBFBqRJ
ZGVc5c01ENoUv55hjBaqZFdE5sBpO5/c4cDM7o20Ey9RYHl++pSWORnBqxn12aeJ
FMiA8emZGOP+tKwSRq+sTregJxC+nnjUhpFA60fZgLMURckTy2j2/jHIpR5Wc1BO
APURls7m8xMzqvUqaFGtYOGXJdKblXsRh0dkslXgl63OC++uiDIpnJZOCp3Az9Jm
CGpwE0wq62UfjhdoNnN1kl1/wkjEVFUZ7AEdytlwUf2xR8V2YcXoU+0SHpey4HV5
M/G2mmXPY2ktWxEB+7PQnlElR/s34PVY605ggO4HQ/jSh6vWoAADcPMdogPqYDKc
3ngyawzhPlGd999ZUyKMV9rzJjInnCcEhavohBlyQpJCFSUzlagL9tuRNFDtJUqj
9V4y8QsC09BIaojvMi8A0SV4RdcVjneDclDTmNfX8YGFkJYedw/Ewe1iHANZIdx3
xJxD29AyCCHFJfjaUuJkJqxc1OgJW3DNL0Z7LGk+Ou9dOHqxaZW5ngquix25LqBu
x50Thk2XbZzCpcPiwfxd1lRa9vyU7gLGf1kxh7L2dkqpUZTGofPowdt3xRdGwkh8
DBWqgWsN5kV5X/IwrX8I9Bp3uvEbl6pJ6nEX5QDaYQcZVGTUCtiXtX9wGWqUgJcD
ruUDm5m/Vab7jitvw9BvZF7RncuUIeFoqL8pryo0oYYMIBx4zPGQSPjnvOVFSkqM
WuQ6MaWe9VdKMV6cSBhMXGtK9A8JcAIA097UrNkQww/PtRjzdAKR8CnALNGVGa5K
7QsKtVQBGYn3Wp11VCVkCQkdLKFd6qmvtK1JiEJ6f9QYGECzwZmgcHZAHQMxm1aa
xTWDgqVyGrK+WGty1K8lEqeV3WygBgHVmR1p2sfmKmQGWThuHnbdJobdOScz5o35
i4jjvfjyiujLwOMuuoK0EOzht2Ddsd1BuSiOdu+UNPWzq60FlJ5KMk9MdDVYKSHc
ycMG82HH2jwrKEoM1mYVSPuKVVTCpX3YX7QVhPF06X+0hbTr+LDXp8MLTcWgJIy+
7jGlYWekEsLMlJBMyb3E2mGOj6znWcf9zBs8xB1ED7kV4uJNgLrfGSmCDylka2aI
uuUD3i1OXgW8zWOiHkLKFMs+PqXPrtR3+gCRFrEu5Lj9S6PTL8L5yhns0zxtiepQ
T+agrhQ0Hup0yhu5STLLxn7oDnkIc2loAbv9oPGO5s/a0ja2wpuYlhpfBL74nklz
bbHLbRbbH45JkwuDb6qWFeAJ6lSvcmX5rY+lgzLppa2WSOtmeIp4MUaZZ0dwBZJ0
JQ3ILlLsQVqkbzGM2Tbgxyesttveh7mAhlDca+NGkoxAjNpSEDOr9RR6ALzAWWES
z0F1AhgQ1dJgBTDuRENzPnLKJbrKmVEOtilP5Xn8kPoqjr0dWuXuxOpugyPYzBkG
NZLlwE5fNjEjV1g75agy3Ac8I5O9rao6sj5I8OLBqR7FncPMl9JVq6hlC2eN1GXq
DnOh0jIiAGvfq1qMIuW2Iig8vHCLsa0yeOpXgp28AHL9c9y0RgevwsGbLL7uR+dU
0jL+56pb2FNgIG2g0vTsee+YYJV2nEuu2b/tTgW5CUAiOgtRAbE4M/ZkvnlyZLk3
OJxJCNfvjWwk2BXsfKVn0iTatPME88LC/pYTs8/fE1m1vm/IbYOhIuiqfn2F9YTI
SKg3EDjEklJDrx4YEAW378FT8L4kv2uCo3+/i/95w6kxzqdSHl4U84bOcu5eNHGt
0VfUYA5o0d1rh/bKhSGdlnquYIFiZMlrSIiZIz59O2az7CmJ+PzelLafz5vuMp7B
B6b2CV1zEnY8PK/6dYWXKknJybC1nRWcqLP0C/WYs11e3QS6cq+McjA4wMSwDxRD
NqragQzjp5Qbq1xckBctRQOntqYFOWmol3hVHjX58ZKU22EzyNJKyCNqoz9HnYom
PUBnvRt3EJR5lQT364DyW2yGyA2pDoOfW/umL+Ux5hG30sYwifRVUx8zRESfppJg
wO2Z2zF/1zC1az/vNaw5gZFozzn4iC7tw1ospXns9hVGa5gsZr7BwEs5S14ATzp+
Kgf+gYjUWAC/SRd/sGuqQ2nQC9/nZF3llvlqK3UC3AqoCSxN0KIO9yP3kpQoJJnh
oXr3GOou8lqan6pNDO+GrSbvLrZ/ME4UfGR7qbor2ZCBCTA7OXcVY74SIzSgmN1J
AM0+P/g/oz1yQ4K85WPwq52pE7nSfCKKis/nk9b4bCvzGoCbC5v7IiSRLxrgI1Jm
lSZiQR1txxy8NZlRioyGjqGDzTytfDTV9jZSWzFEPE9Gjh5U6l8VlPNhE08Ax4sg
U2kC/pvA58P3h3ctNzuwar8yqjMNK/ndp4kw5/4oWAFWOPTb8HKey7Nn/KStQl4m
CrcZ2Pcl/LnbSyFZMwb6d54mbYlwh+R5bZnRkXpvv2Qvd82J9VcL2YhvzgKpmlGU
AbivZqlnVyfuO2Bn1pmJI9zNDxoLkvO34XH12N1n1eSekYP8Lg9IqzTqoXRHDDJU
+erStVi1HJhpHYWB+wNX90KZ4FAiZqgRL1PX7vJhAEOqWZAOC/jtWs91sGmubv5O
`protect end_protected