`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH+OeLAzg7TC7xTfxyU4d9Liu/pG6DUtIN0rYSPBaZo7C
3RftLiLv3lnj/KPw2lJhkfn8DFW+J8k8sVVl+K0S5potGTt5b4c/hjHEzXCfqpnL
hv4OI3z3eNkJv/n8GQDwGbo/Jk/oQLXAb+/ugWEYZM7ipeoAfQ9GkuPsOFgCtbKJ
kiS+9beOPo0HM4SnLjHVNn6pBCr5wllijcTKGBQSKc0dfpLyvkBfaAM/GbqrPniM
/Xp6WgG/iDOin9BuAdIHUV5jMY26YcnTgaSBKF6RSgfhLeLImDefTv/2f6jwptH2
WbVd3W+WxJRlk+ONTjABK5TPSUyfOlX4wui1Bct8XdNOBsf1cC66PCS69wZ8ysdk
mP2SiWSMvlNEdFV+yjS0eFL9dBJue5ZWNN2BL7isnJSXhql7YKjplrhn8yhX62mQ
8NiIf9amt9ZYEwPsrkcOlxR4jZLBrXBZDBQk0D9zRr6xpPJvjtGav/TH6wvii7OC
03GS5Ivy6ciAqmm651H2SkvhL15/SzYxo20tsrKqNYWRdVHeWqJmjRtlVWjViiHe
JCKGHM1CW4KrxtppfOgqpgw42ZawtfTyDk5kB+tu+Wz+cI4WHs1oeMGmniFY83td
zHnQCZCXuCMJh0Nj2oh7HTLdZ75RlYcypgtQfDMF28vJxyn1F7Xpxos5p49r3t3s
jIitLreNP/zXGtD1Px9luHRoXEj/da9gW1UUyOUVqf0m3Zv4wkE/X3etPxz4KLvV
0HvLgboT7+igSlrp5MuNp9UAstN6J9F8oIZpL9rwBDPkD/ZbSjqkl0c8pxGzofKy
mzZGDBRKIdKN+QLV16OpR/HFIIupu/BcmD01WLLR0w5hlrubYqasazMKIp1AmfUp
lQtXzhjjHeT8uiJpzq7QT/jO0G1i+lS0XSyFxqUacFrf8NRfK52zyRe5j3x0Zpkx
TS9jMXkqBUYsEVgc12D4xOQo6cLcX2b/wYSzrtQBN0i3wGd7R+2VSPuxoaHw0gub
L572NRvBQ8atW7V+PLNUrJaCedeHsa9cCZZ3iEyMm/gMZ+CBJtBW48yrIIA3Y9Du
IboC+ju/iT6jd1Lbft42PcDNDNmdIn5juXDPW0rhBi2Ifuwzlro8KMFjP6LKdwEg
XZ+Hr4lTvjWqqzSRAi8j8tSojT942/Jd+uMdA05ZjgO3ytXSRbkOEDxgwdgy652+
amkmyPpwC6RgEj6iInQYfzdWTvk5DFo38EFeYt328+lhP2e/wKXOyYo9twFCq3PK
nTwmqJKUOBiJKz7r+j+D0LxxvixtbyUjTIOUOuXo82JM5SC7bX2kMAr9mIa2HYtd
KE7/LVBOGXlu72pIcThwytOhpfRg/09T/0XUeVD2IgFsIE3xaZ2kYv6ci5yeIFei
F8aK89CHYAE6j0fY4vsEwHS0JE4hJm65Cp+PFnhJk3EvP1oJ9H5ybKABPErBS5Kg
wOax2+e26Z9M+8S0jL07LhDau4tyK47OPPMwQb20DiJNm2IWk3ZQGKgWkSmOlCid
H4kPlaERQE6MxQlf86h8ACw3B6hHSZet0B0GWLjd5IB8/0EtJCYxe6PgqKFvJDlV
WvJ43olxdUsl7CFMSiLzUxmbq74MslDjlKxGwVu8MSuoPHpwXGZaw+saD22mbWbW
66o9Mj4gGQuKF2JkIza0Zkc9lkkjDqptbDNwATyCM/lOoKdmWrlV7EoARzob1m4a
iilm2M6OrifmV1FcapZs7oAiSLJEI21ulV7o/VF6nBKhI5e+I5u2weuMOHE3Sk3R
e/XH+LYl7VioMxNlMiMrbWh3moWE+NpsY5DAEY+W5ON6ll9g+PMf1ikpmgbox7XZ
FPVUihd1On3Ruv3ofOKxv/EPov6IhBMrp7Xj0pxVWy9Iw+DioamnrRO9RvjOhjp1
BHJzE32Rx8U4G30zJ7zFXHX+VnCTaIeFyP+UTJ2oeM20Qq/WtxfHzaZ8R8Y/ijQt
hBjdM0swGQpFib2HyAn8uDHIyk2wWt/OiPThAdQPi5GIQfAgJ2+q3JOAzl0lh07C
oJXCO4x67zWurhsOhWz2QyHkJ9IAS/sRA+w3/ZfAXSoxMJ5SrnkFKhf8S1Tugj9o
nqJYxewg3LEMlVs+Qtpn3OhX75dNVHazfp8QbTNNWvz2XwRRkD2WrYJyV+AhH1Wy
GqjAXC6l1kF4/3zKamS/ymU4jjWaL4rzxsKN50z2Wz2V37r/HiBdOZAU++jsT4a+
RmqVVE0mAnq6Bec3kkocNav/d11rb/5HNOURfShP3oSfh9NmK4oxzmhZFqgoriR5
Hllfgz84h2q2uy8Ph5v2Z+G2y+32O4GP3HIQtCcuomVdD3w+iO4II+aO+Gr/2VfK
9kXjeUjtMVylMU+k53kUbb0dU3p0Ia+UwDiO8Pe62B6KyfITPWgOoCK40zBtIRGK
D/cjvDK70mXVdIo8uLfpDgzh54IWg7mHAJ1h9aBH4bpLdHzUh5YmRoL3GRf7OqYH
OePSf7HsgS1vgLxfmYrCyXOMGQHiileYZJ5vIm14/x8nLPp65uuErkncHroVPbQH
xTgISvy8LElKt8QF9JTtz/r9LfzSNnVw7fOZzru/c/53xDmOXFPWEkRlVv1OrzoI
XkNhZhaiQPZUzwiuWr6NSqzXo9PHtqmlmLQs5yVGvdCge6ydDINJiPRS1OS98xqT
UwQltOAyjyFrjmmCUGjkd0Ymp8hlhabGLHqX7R9K9Q5kJZC8Valg5DLe2y70fGwq
l0prARkgUViP5dkbiTZ0tLa4G6+E3xXcpCbtwLG/3zHDmY64wmNW7guKzAvWsXwF
ek0IyWP1I8TuAaDmWnJXwNrrZnfFBJO1xL9fL8KZGFBA572NLmyxOcjEyLyA3xK2
3Chu71/uIyXOLwCkOht0Xafy3VS28FnST+gZo4/zuK7l1uDU6GRdsHTO1xlL1VGA
MDIjLUYioxIALvsuhYaUTmt1VKy8B8vXiIjdYVjMpg1MsltvK3d/hzgT7dJmPO8c
N8H7Ar3gr7VSj/T2S/qrK4Ud/pt5yG6DmsFg9iuxufPTzgn9Yw1/7yNW/NPQwNW6
IsfetO4AjpnjFeSGl1z+yQs/O/Su9i9AzIe16//3v9xqKCazx3QTjFbEmU7FdRdm
D/Xl3DwkqtNTaS8OnNA9oyD9cNPkkiQ4fwlan5nvO+I1Qvfhtf/MBRvc1zoy1kdv
FCF915fgBojZ0jxq4Oa4M/QcQngZOzhXzdhwlucZBiHGXkuwiGzdn0x0+8hVO3yZ
lGxZJP1PepgtQOkSjWY7YLcUWyeeDDaNHle6+KI/bOVolubsKv05JctoHjmfhpOS
Cus9lKp0AsppEuKi/3dnxPQOiAkGb+lxUHdGAM0kNAPWn5ZF0txAjYfzyXTP+zwi
NwtmhMeeeM1IAiNzvA2La1zHpJDJNzb4VpvEcL6xQknl7QVijNRrikJRVkIRhkYg
U+L/Ts/phLSYUKY7kgD/1OqC4sIwRM/r95eAGh78oULLna8Eo90ZWZnRsWF2LHg+
9YQXxvyG0mSzCPcPeH8hPCjCOzRBwR/nLhaPJOk+BynYipcR6uV/34Gmq+ycHfDt
N8ilRS0av6U/6zHqOwoxWlY+73XRdS+8t7mkj5LImgURfQh1tYZlYJlELjSmb12L
12QB/NWfVN1CRgtxbjdZLMZloB9gc5iBoz6TCqiF2XtRCITPngZ6+zzd3k5Rbt38
/ZmA8rRvoadvsexCUHdXiCd5iNRCnIAFy7rMFQdX/j+pYtYZI5kIEY53aJ6MTul7
fc4wjU/cwS7iE8kllpFotgg1lTcDPvjlS6gPYImlqA9eXuV8Vz1adRcA0NpHQ/pL
RwPeKS/5WRQAdENCmpKKukLIKvyIx54oFnWCKLvNZCHHDpBPIFgiQFjJwSK/j9fJ
VIeMdZAtweLZnCCSr6MHW/B1R2GhFRE4C8o7/t3xW12FbNaaIYUAKQwtfOG/hbIs
Spx0/oNBZUDAGhspsaHiBZQA6dnR5teRz+qvjLDmtIy9DUAwoNkCkweC+hDcdK1c
XNqRl+iwDRiP1+fQ9qDRzvpRt1C/q1XOlyRbqtl01uCTZkmrIhylNdqAIC7Bn9Dk
v0eSO+hls7rID/6tGxDT5MzhLvRkUZUCsiZhrsyAnNNeuIgdJ1CLhOL9Fj5sa1bd
aY2UAH7+r8wGzwbS3UQQ0tWISQt7XpneA+bO9cf2lyn2V2+U+hTxhR60RuIUkblI
tmaqNU/3YT2T6Ecyrpz83Zq793p5YqTsWY/rmU2QE5B3YmHFzcvqnXGJ73uXqtv3
QaCATX7QKJ717kTebXguW/5w3e8EXKG7FfB0d9nAo+MkV1H9d0fI0gqZE0oFWt3O
4fxedJqb6iNggUdaaszwL+wgrTO+n3OHup/9zqzKSHQpyC8RzY/2OquKzZr3Es/W
B/4iIehXJ6vvLuC7xPEyl8fOERNo82pvdTjLxL1+Kw733nu/utlidn6gpKeO8AjA
MEOCsM25mqaZ/O8T75h7TOKv+sVfa24FfZVKhAoun0fdnJHHsUIDGrGAimt+aa0u
BLY4Q6K+M0kEirLAKWxSRs3gXhk/qNNwIU2Ksg0757VxDQvC1q6qdRgNTh0qO32F
gB09s7wYHyMouE0k1OSYWfVA8mFRM2pvArChqSxGeyRqbiWEe9/uhKN45BdWIwlo
9l65XQ6AC7foXB2pCZwhORVLPqsmjrJ18r0qdaMpd5n+aj25pqla0qqzN42ziaZa
izOBMmYx/MXCuIlTQ0mKbYmpEC9ER9WGpS9NPnZtfhmkqPpDfsvnZtK7LDx24LjG
FBeLKb1iZ6odXAKdRrzB7tzLTwg+ZwUVpghLJQwo13TujMAYZeANuT1Wx/mHqHT9
HlzdoWCSv8VRYwi2raq3lvqTC/u/5bmR79NisoNsdK2uSnUT035uATAF6B4o4dEE
HilGWxJo3KM0749/JAvdhBVkfmwmxB61NxPSbXENeOcVPjACzP73BHns1Ym8mtsh
8w6Fke5NbzVVyPwjoN5hY79IgJX9ZnPxqay99YZ1MtB0XzEPLCa6X70L0lkntI8X
wvmEUJzO9AcWASYrs/kNZ9idN3pZnTr40zyA5bZfLOOwYCnU+jtfPqvqQ50X/mX9
9KAS8q9CadF6cWgDuvTAlY7Hjao9bk1y4+4QCmTpsebcfl+YThf/j5BHELPfDVU9
+CxxwBCwqU3hGHATzE++xOT1wq7+tqWHXNWguMPJFxAUmdMMsc94KQkN70x2W3F8
YDouoHFM7Yj2SXLkY2by/+NmTZ3z1DVtAoS0o7QoQjwMW/tAiuHg47wbqFJR0Ozm
0R8OP79MbXLRP9YItdvicLgY4dKqtaKuQBm8X2ez84zK6hX9ZyY9/+SkRVp8T0f6
1wp5CwUtHz01qrmps4lbVk8S8i+86T28ZnLZ5mYGjuqmDEIhsXRNjVhe8FKX9u0u
7NRaAq5E2QtTxCJeTiH+xQdk40/0utzkk7heKKF6svW9lwlovVqORXOsRA7CeNyp
+k4XXo/frXXpaUl3wdFl3PiLGSnJtLIicfSYTtkgxVI8ugiiW63t6Ex2n4fFm5cv
RbbnCsaT8MJn6H6eKoAjVvzPC0rLqjQfw3B3thtmAV8hzor0G0h5jd3l5cVBLHvT
0z+/fQADbM+2qQ4VyKiT1Pht2iETcrGB5QIqYsChNTQNkr/IeOKuGUVTAd+U8Gi8
w3683N49DMe9ZLd9Rmm3VNtwdrIkJj95cbqqjNwZqLSzGwCvb6iJi/HZG3K3rfPT
KNYqi8JGOFwEdn5XJfrrM6bUWaiOJrDAY4PS+UP6DaEBbqa8gMJRWw8uz7kVxLqR
xuyP0wH1T31Qpc3kQUTZ8f+9iPxChsHTvOAvDKG08V8YCLTblDBuF0Zg7pPj958z
E4dD6EOXhTujlVyzKT3StKId9veppRHFl1jKyNUfJcQMO8etFg18WDIAl+bkqYtU
J4vLchlTEmSfQCyD+WHfPpdmPSMd0MUR149QvSSaXvCwqUFJ3k/t9Kfv9axm1mt7
yzmsQ5CStm8UO6hSiwXQwNL46Q5b8QXzcm0xkbfx/JX5xzknv4Lp7GEC982UDs4X
f6E64jd8jSUMfY5M/BPHfYgQPR5BRFutyERSth2Kxn0zmbp2R3YKa8Y6qnKTYcR2
Vdjmsn/IqgW+t4WWBq1kZvYfVQ5n3pBW7ye0IKP42NvWtdblP0wQd7ZI849Lnc3M
dZm8n2pyGmWN29Eu5XQeFBpl1vNhGoKETcsw7d8bBGdzpwkaV8SFBrnsTtBeEtEU
DXk5Cd5djCq0HV2/IW5WLf8aCD+bC7GG0rYVeKqAUVVzNBdK2suTfDKVZoWdF+7a
+iXSuB8VWRVPLMUJChf2Dd11qy2S6lxvBN1r3CEF8nGFgXx229JfZXIquzLhI5b2
HfTDM9JJYNqqFRNa9R8SaisAbRQJkSKOcZfx91dOD+byJISvnc+GzsdfdJgywk5y
n0pWtHza5RV0LmLmEwFOkj4ebBBy50tWSAzggFu9HqYmVT/UDtoxxs9q5ETybObg
y11/0XHui180DGF4G24Qij1U15LgHU9mw4tsfj05nYoiVClxN4+oVGsETxZCTxsw
cZh5BTMbItYFPBnkDx/FNYd+fM0v2k7mpaTa2oA3pWH8zlKwS0E8JfU6033qykmn
w+FnoKlyJa1Jrd8RWkvGaq9Wj0FLhIJCAMSH8TpgOyczdnATHI0sMiGYUEWC+ID5
RM8Isu3u0HugkAWqdFm7yM5I2LQslv1KMVER+IkQEScZN7YK2XxSLSjk6YeYcSsu
EOKMTW54p9VLjL8Lj5uHQ7xPLMBy3EYZlQC2KBuTXCnx51dL4GTXgbFGkRftx9pi
hEZKy/oB8FnY+HvEG4DFB3paLR/x/MS45cZNhDuo+/KO41p7B/H22okxAHCSgfqp
GR36D66IJqG5r3bSiyK00L8w949sECclGAIbVXaZXrcy4L6znZ9B+u2NMM/qKjDA
P3V7S9YMa5JpWeqOa0/CaK0ySzCKqpYwpaRZkN4Kg/dUSX93omKH6P0ZAj4wkwJP
i/Vf89meupa4fwDoI2QSY7Je7hAaWFgtMqdC3EG7vi2t6W1lyL+1ggodYH+Zsbi9
+tvWkr5yTCGDcc5gqMTj190/JOc/AfUoaRze80wcRf6R3mpZYZ/CPZti+e7lNw75
OE/3bhYhIfxiiKyhbHcl2AUDjZQ2eWIqzRh//LV+rjY7Kr6HNNhEqToyVLdJLh9u
cCOm3M/OXcCpH1dllsN7XJVp421JjFK1YLvLJ8sl6OAN9VeaSGKUM5xhDYKanGOu
T0z4xggbA7dT4tc9R41wwAVay5ByoKERSGNIchky5lsfCrCnDrq8uYM5hsPaUHtl
2PB0D/DMctGOT+4UqvxqCY3QKt83mrZ0hX2OOtYvJS8eMFKLxHHuRub5Gbg5IxkW
8E+26xID8gLvnXKZGh5BoDOdShmKIRmBiDDEBZmSgjOZNUsdk7eaCTonS87FLyRu
Nx3SzOsMyVFmsJHffqkHe7uqnoefebZ0kAN1OX4dndel5Wo4Cr1AmkfjWnPs9YDX
bROni9B958MAihKIAlldlsCGgQZho7ltG/6VQB8Xem1dyyPyqmiyE3nhZrK//qV7
rdLsRUCJ16a09yG885X4IMmzHUcZ8WjnIHztMeyuNxPELvkHve+40lciS7Sc9Atd
XnXRP/M+Az/SiVsbJSyM3wPO8DZiJfbwOSZv6bQuBXvHGtHw/0udoy7lWghC6wnQ
qOqbhRSGAgK128XduWJPaHV4vmgElPBM6bCd91Nc7Hi5OfBuFATCzgASMS4KqXTX
7zkd3BZKhnVUTV/a/SIhR9aRwJZ7WjF3qdi6l/05RZGA/xlTDureEljg6EI+d88w
5poRTioFuUarLEyliPobxcrGFLapBaTskizupAuRh/sTj/tdbyTgGM7u1ra0FvDk
oZSwiKxh661370k951j3cc2niBPr8bCYTDm1lUHKaOoxMXl0orOKD9Ptseq5pvxK
GpsmLT/xQW4+UdLBxqhZNAq3My7mHKIqjHpWqL5LYNT1nU1ZunPdywNtElCaENOO
twoCoR6tAl6EHjJonjSrBBxRewQbNYsqBnNJ54+sgeEDNHtyxpU8CFgxsK05IY1U
0jWxnz2YHNtVjImary3FyteElZFPLQlBQvF2y0tZtn/ufTda6NsPBzJfeArrdP4K
cq/CK8lnVa4kLrk7XTpTfite9s6B1vTgBd2MjSmqbZMCU1o3GQZtIWXc+Yibpvjo
4ESWHIH21d25nhRH1kAE5tzqEWYPdf43+Zy2WZ7GzR7vbuL4sZrMkKmDYP8F01SJ
SuQbTP74TzIr2kJltx+X1zpIGOFBHni89K4ctfsxt4kK/kcGjgfhttfSoslUeGc+
GS0uB35DtskSY0CuqyT/cPy3xj5n/VJWiAlSJa3Y6thI/tsHcfeaN1awlT2dxsYy
HZlYZ88zwCSKrMVJLwdZdJ0Qc5zwvuPbUdVoM4QBtX6H9zcQXy7Q30EHpaMyM90J
RkPtO3KG64VkFkjpOB5tMA==
`protect end_protected