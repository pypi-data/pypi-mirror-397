`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
I5JJnrdmdIVaCewvA2Wm2iGhLZ8ObG59OCv9Xynwv3RJOb1vpsbem8lhT92Cy0kR
yi4SqGerZMTJn+d3KIjtbFZbHdyeaU080Qx4x//5awpoXD61pTaR+WDP3O7sgEac
zyJ00klSeWH/uMOax+oN8JLyt9DHveinTLNBDhMHQsTQbN5KmVzldekCZCUgy0P0
J1xJ7DAXhZJwrUMIxcVtVL+dSkHB1wFRKooPA20rnzNLHqhbZTEgRbnecL78t+Io
/KowS6nkLCJyYs3bZ+1vQYFtjUY6rGbM/cRqKEgxKgIPeJ/ZRYWD4woZtDZYReGO
caAL5swlZ1VFRHvzzITCTyxhaqeWeW3yCqvmCrDkHtRAqzB01J81wLleUMl0KvB1
5elWFyDUy3bLg49GfVJB+mvSZLj7GOcUQMlBC8uCFeb4HBsk2Cq7jycbBHFxLe96
cdQEekY3Az9a2hIc/kKJyqm6TrkCxpBzQwtnoPI/6vGiRo6FIfdOIrG2K1g+8p4T
HF65ZYoNEpbyaXplEYkmizw1GL8jwPwEO6geRysCVSSJROHdd3p/5FOP84JtXNeo
kSjeLNkeOKRkry2E94B9wfgdWE2cJT/NwKIXsx1tJ7yzQ/HoKqwO/75+X//M4VvJ
ouMDLJSzFiy7WoOC86h9oucM3WC0nyVMf2P9gARW0a1DV3lIZG14Oiy/6xyE17So
sS0Pw0Ihou23A/LGvKws2l05oOSqbIGdpVPj6/zX/TI0HnxvTSUAuTZL4hKFY5wX
6r+cA7zRfMO4g7sefI4bzkLWHiy9+pENGa0FK0qKxb4gxzvOG6zkPW0/Rjdc4/Ek
GE/JH+I8f1CYqtDzdKgJHKwgNKupz9GKFxmDJnRkr5RPL3KcMb9xXDr0knJejB+9
xZzeCBQOmHEK2/r/ML6x9DgRJ3i3/Qr6q091Kq+H2kw862W6uVzhdLb73NZfdvLz
CT0/oU7cEzeaOOyZf1QT3k1FkEm46VDHnS2P/pnBLgznn1JZTN8sgm6tbIfTMitL
ol+OycHrtgK1lZtHtLJlFBv6XnY077fWBFF8Nee0blansJMS7H2CSu4vPteDMx8J
ts2HvcNG74UA/8/lldz+7EJqPIDeOiSOw4DXbPSO+vn/3OG5coLDXHwL+31qu0sx
aauPg6lnV/4m81d9CeF3cLWouAwMx56nylseDcoMK29IXV7Q1RkRAZadgr5Ns/13
VnagaTe24o1i0OkaEgpZYoqTWMCG8LYkeV+a453jKh3qrILg5iHsk/Zl30O/Q3Kp
/Yi0Zbu2wDG5JmieRgXykQQb+nfaIuncp8t1Q7nHP2wvpRA6LiTJByBFbEsHN0dO
m6h5qKnwLkPuOTTox6fq/pg6zgR2w0EMYgIDQw2V6Rpkr1GDwRiVnIh3QzJ/By5j
z9RC9XacsmxsAhkWXul/R/P6w6Xt+CkAC9QKPVVtQ/RTrVlNv5lhSgArMo3bOOjj
ZJCHl1VCGR2Uc4vCulEsr4RJdEecLcKW+VMzIJGJAqcdfhw2eVFsPU0Z7VwKQqWz
nvyVSMXoG/xyibDengVEvx6eyaM7SDZrQ5QMZXxlJsK07RJQvA2p70rVHp9hVfW3
w3c6kLw9io8sFVxmNcLBSNf3PtTFj32S59LwFgCnVVoQjOuzPYpnLmmqekj0Pka2
ZAWCoMkfA5nDl/obseXanzHb6kx7IQfsOIYgznxapH8agouLfrOFSf00mlWuc1tt
avEwvGVsP0+K20JCk6G0n1t1TUqF1806CMtCU821/30KvEJ9hYWcxr0jPWrPtTKC
vNHy0wJX3w7lmRIvr2qmuM7wWBBPVxCWozFOkQXBNuuTYIBErwXU5gaJsgFOcV0B
2XL51in+deBeI1bFhSyhaBck6TSzu3I/6njglnVY/L0yfN9C9sPbd2PB7tX4+83K
qCNklZB7f2rjbKgXVeYfw0HEIrMT72/NBobvaemALN7smbVzXsENGDNfLOtGK0cq
S9tVgAU6t3y8F9xG8ULXssm3aATs1BacXnm8ZkBI2mUROCkkawxIzAUW2GRnHVbV
RqCBnbUQcIryyMBN5b6qrxUIqsW9gAXtEv1HnsvJh5r57zvzFa38reE/+IHfLm4U
qPOOUAHC6y9g2PGi6BUEAL/LGgrywXO+x/qvxzRFp16RckYj2t2mpxXa3Klfc9e7
7HsH0o3D4A5VFzIZqYfUXJOhqshrYn67HyiKJfAe6keSLyFnYRf4VWyMcjNjpbkd
SAextFUn4IAH4CwcQkhbgKYMcuaUuQKgIr/nl0FE/YEo6UHbG9VZYEQ7wg6mQIps
tNbNUAgQADDCao/ib9J+Q3FTMtNRi9cP94xntoOiRl76YdeqQsIJhV5BkWq59B5e
8GUJDU6TwNQ07xKLamij2b2Zu16VvMcNPOzV6RLOyU4X44CD7RYa9T2wZu10CS5C
HYkuevc5pcH13Y9hrF+jeVo/0VSDBQLCyqWPYRFdsUFTLh7ldkjUIuTEGheJMDCD
Y0GwW3jioYhhx7Fuf79lyUqJsTVhXL+Ye2RTu1kihQuwQp/VN1Q2FbHUa6m2nCkF
/LuqfdMszMBw7hl4hcRYChJnyvsIDzisRH+j9Ytr+EPecko+oBuhGyyvKT82Vrrk
vkqdVCCvgHL5xXoj3nqP1AQSU2qZ6RuO6W5W+yi2no8pmNdwybEKLUQLGR3rbWYC
ufMgoe59u8JpNsF96LlFT+sHLZPCoJ79W2zkQk8d3wefiAdDyKexhLl8bjGUtaJs
jC//i6Xx63UmQGHRaIh6CMyRWcUn4lie/Sv23O7A+PBzBBbetdxW1/7wb8wfK2JL
9oUiMdJ6GUfu4T8QzH5zBcNj20CjAbQriwGFx8NTwZQODIhd4dKiyZRTgnln3C4p
W5HYolqn5231a7uQd/JP610MaHrV0ByZYZOAsahbFiCW2Nngqb9HfNWvuuMzpwA+
i5QXjijHQY/0NepS2/lieI0iPr/O0Crei19bjMebwKSYnqZ0sjawlY3SWPVKKQly
JGQpdPZHJ3CTH77qJ6Kpwe3ntqIpeX42Mglb04WZCdmCPpDzcTrlK2GDO5kHVSmf
jI6JFBHl2j7rvGFRVXTclKq0m3OqJ7Vyu/eYATVUo9QpawzPUio37aDioMqAVlGh
sp0t6TOeBRwYkYDhxn0NyWAH0yJKYCrXZQae7D/XoKrM1VXE1a2qL104yyOBDm5d
2SfAvQBjeoLihHr67fXGXMKSG8a8tfiBOaIURaqohzcmIEvmUO8dvn08ScUZ2DH2
k9n0R8qXAEWeMuLqIyxF2oc3mxpxfudcxLbpvOyi9VCMDPcABoomvuvmDJhxN0gf
ZKyA8EIJFbbVIvOuNZY0LZJbGSOcMDfndcuZKagCVvcaUBA1uuwFqLztCzU10Ajc
Ou12SiZ40wMnnL7UIPLd0hd39t8PYSOXi+2urCsqGN+257EQt6RlplINZQaHQynY
J4w8yzW5g46+Rry4HTPN8JH8NNB1kCIoP8s0csID9Nz9VmKnnRbtyQtKUAJ6BH9Z
PozWWwJTPTN3GkkWnVmYl5Nb80l12h3TyewTSdXdShLUH/DBIoXp93XOpdNHeB/X
oxRKZ1L4DrZHZ8dsw3ORSSAeidZuzbGqudjbmnJP1rAEESoTnsC1Jc7iSNkrOyhP
IADfCN6eNtVEcogQCveY9YbUv/p7y2zZiZA4xQszN3e0/BTFY+FsmqfE030kTvgh
bRwncPLdTGCU6btzjaeVt+MDhMChNunzKF8Wvz1++lCpsZzIyRw0o1tk7bhSXYC1
F4D+jp/JxWwFjJWJjv+JenuI3YB6QOKY8Rk5Uyy7mO4sxsaXAcuAx72cwGkXPOh0
rSY6X/SFxcvBK6UQdx8DygByByXo7f2M93SUwyvKJwtDG4cXR2llD2zkkjnN3jk/
avtrbRXshgML8OF1OhRl4BI9UQq4iNcocjh+NP8ENVRjJY5rZQFTFq83wcyTMk3r
SsolwlKCa9x9ZbkoBkOPvdfZ2pwpM2pPaExpFKauzdHyZXFboABn5S5nkujVjevQ
xIDOANnne5N35XyTGh2Pb2nepYg9fXOiM7SvOFtt89RwAnA5FxAUzYQX6yCj1qsP
BdUnZLQ0X6zA1EuS5fwqf3Ttr8mPvzaea3cp+Ib85MMMqVKCv2LUP5HZDJ1pPPTi
P9q5Ots4S4cY46zbyUtLz3x5LODs3S5UcZIQ6rVdkWzUVYPKfxVl4trszNMv0Ek4
1XAIfZ/I1j9Wim6Q+9wuOMbups2X91iOr5s7ktDO+ToA2kmIvivdsplh9AFXOC0B
lrShpVDSWS+4U9l9qByFYFZX4L4nTzgzyU7DuijDAXa206+SvptybxLBgWT7EgLT
zcxfnA6X8afLxIWT0ISijhHQS0Lqz9O3QBFl+R5WEFIcauhoEOG8m8/0Pxn/CP6I
/s1UPGXQZHI1fzpsfCN8SO9F9l26DEkA7uD81Xv67RW4VFWHs+wWoCYhmW4U2R2X
GNJV7O2IUNxKmpqR46ruk8tufnV0euWexBFsa0oXvj2LkkeFrHemAeviZ0KsW5Ms
tc4vLe0Zp980Xxb6HmqSbatG+pVvQH7uIqno1AmX/2Nrw8MuASTD2ZG6vsTeas7K
LfPqKB6n2lKWZH9rvo1vVTHnP1nDARuVtkDnW+KzyWpMqflOIeGpqo3R0gzSZ5wa
Q6YK2YOihAD4NDVgarvlZIxPuHcds3xWD3jII477CGkCdOWB7MEsuiN+5zGKo63w
q3LtKLHGDaoIR8LBdZEuPKRdUJ+zx0we2nEnxv7z+TQUp3U0U0GfSYhcTzGCWwsq
1AWuFMAPsJ7Z2F4dDHng75Tpu9JQWesQLmmnZtJT0JWKlCU6jh1pH4/uMtmF9ZJE
omsXtLnONRwM4b2LeVer71Ql66VH7HZQiLWyctJVQ+BNOoL9u55CDtR3vhOd3GIm
0x1yg/12+5THziE7cr7ihrgO9IvDB8Z45t6rWfQAGIaYm0eS6C2Hsmwbg0pDUCHf
66xAAE1ato4N6fAVvNX9VXFTdgsQHuVpRdEO5ub8ASGglBXKvroHagDnKnFwrgnG
FXmkKHss5dknrEVrywLsQplFXGaJjoyAtP4VsbLuWuZ1ArqkvlhxEmp+2pSDrbUJ
FIQZ7eg008Dmpr3POtmS65m1xFLp5pZY7o00AsODuopc7m6r973PjI9B/Jq1CH6J
+87AOD7RWp/uVLVvvXMryO8zfXQRsYKId982gE/NN8Iz0pTwQKUmfGMVGouO0rme
7xPI3OdZeJrnvQrQPMc/FGSyc0V3i5HAH/kpV59aMUgUzOaKaS/QETOQWLrlvV7q
fyQ83MH/6SeXYNlJOBNNSJGtoDIHTHeM0LNKIG8hxzjyPpGc7ck41LnJNR/6efS0
ZSxtV4nF15B7PeietbYWXF25FK1hAjHX7BhQVeLyEATLXFWf0zDHjXeplIq7VPJJ
DWGxKdw9yDbk+PCjAgZV2Oh+T/HNQPY2I4mU2c+MAjPhyse3bJH4rvbvX6yP9/G2
hNipQk+kNAyUwrqTHt2f8IqgVbTZYuQlrRr66dpNxz3lPTkKVvi1ahymXisIrYQn
pCgCQoKZ0dO5WOVD/rxRK9/XQRa1kkbb1qo9ad1jb9JO6PkvV2JUi5NJgnXnkN8a
w/dyJedJ4GDUtLms5W7AoN83vwFFAPjiwlxdTjITE1M/Rg58MTAeQqjXGRNPbCgJ
eAHtUcsInNeIcjUsBFnWPMraP1AK60ekM2VIPKRRrmec0WtpllM9V6K6P4Figl7X
meazGRjJ4MNOBwwvWuzF6M7e6j8ngEcqJeZJl2eF5gTHaKuO1poS81nybNCJqtfh
iizIGy7HuL47Ev1Cj3a1vtVlTaaebE9S/a5V5UTcdt5XrMYeNmvcZsuVQNH3k5iA
CnfazZyFqvhTWz1xPpTtdHt7patRyMu4gEHt2UZtYuHrsEFn30wPNvtZJsmldJGn
63jEp3uMhnlXusumuKYsAw6QX2uJPAgyn3be55kP9HLYwPMvGuv9zkxc4QMjBNgs
GurBK/j/HkviLzPtRPPMIk0tdR81he3+pvrXYXMf727VCUPbt3yZDBcFYaGsNSnu
xBIvYPA7sQPGcT1eQi8PvmsoteJjSd/6dZxjGDNiHuZuLQB5ifzTcr9I32nahcvG
CGhF+j8+rQh+tGaTbUcJmNuG2qDjCQuRNX2816vqL7aFkLJFNVq1PbhiRqtOwH0c
oIoaAxEBzMBMp3D0GSNQkYWiMXeSfROb87FOVsCUs0TRwuQ6t7RnknmPK9vy8NW0
F2KEgToYhOSLutAg5E6WRUsYpxHeMbUilDN8yhDhJNTnI/sVjDI/HFs5zkfs+YLt
OBKiZ7a4CNdUP1aIglj0Acejq7hVoglrsQ+wSvKPrW6Semci9EiYcXd442ZM0FwG
1hq0581Qy7N5FmKT20/rEIjcR9wrgbQf31EbWcudx5gnJkDnYrADFfVDLtt+k0DZ
bE42vnRQLBBsibfReOLIEZ12nX9raqF8VNOlGbAjjnEzLRFX3AiyVPzDqK9VEAS8
zNzF84V0MNM5FF87Omx+Uh0F7vYVprCACbQof2u+P9j20Znlhrg1FUJ709p/I6cl
01hzhAKHyfeT0ta+pS/V9Jz6GIGSxOhh7DOOrBm/HuCxegPK89hO0TVriE1Qwh6/
OsJ1PAD6sHhUMEFXE637D22JNUduQ1a4Cy9CyMnPHer8X7ueHpgxW/ZXcLnKHoIV
ejgBKc4jZLpAN5wxvhT/hLb3qaMtGfGNZForIT0MKtddH+hKFKtjOtW2cqa+WAhG
PnFDdI6/gWfLUnxOlTu+Z5n6FksTM0TJLSMTeeNxmzRyPUpEI8moKAHPm8XgNMuE
dXjI/CXATcPQO6sEB3/2u8GAiLcBuoMoG0chNFuGPqSD13VGnfITgMMzS+LLoNkx
ID9ZFr26bhFudqoBmNMrZfcd78kMczYz24NAqjW9MeVABCJmuiJ900jGFKNpi359
+2+YMZDRagrakVZSPg+cewgzQx2eSxnF1Kt2gIPH6PYsGxkVmMvb6xvgJ513Hrfq
9yzMKIc/dgoYYX9GR2Bi/U6t9qvhjLRIqDKMTi6UaaEjOHDMlM33umL67VZXVhey
yAEZ63YlItkhgE3wEpR+gkXVgjllYH2oG/oZn4Y4XpPOc6AsOL4GGqYtKcVe2XBv
thsUVA2w4etOymvYboCIJwjIrn1Rvf3+BLVrcUiS/7Q3Ym4Ie3ricTflzHghGinM
CpjFDze+YsUzLEdBI9yxc5leVerUE5lDza93xOCTCrN7PFM+ga9xuQeiwgsobeCm
+4+gw+8LjpGYsKFJiX269QwlIU88vsRREr5ev1XcQiK7iXtPBG/AhmtVb0PKpweX
OCAxM9SaOl0iXx/UDOYM38nx51EDdSeuXu3cXcbW6VgWgbSPyriBTCzR2P+8o86m
QcPiwFOxj+RsYQyd6lTPGHaKc7c6p/llJgpD/PJWCQ6YkGXoUH2SRSKcnRwEFgt8
vJgSYRv58nIrksGv+12Qhy/+6NajUjKhrgIvMaOW+HKEDRo10tmZJepCPSH60F7L
pbGmEy3b3Kb1L4igKhTmuVnf4MLwU6TQLiiKGs8pvV5V7tAgsNBJsZBQHDZB+mHe
DrgDmXqX8g7BU86q4b5xmJ6Fdcpg/OmAuYxHuZWTsPV7MEK4Uz0frwXr1nXCWg72
U9OyvELRnfZ0wwBOAWQPjKg/WS1boeqGf4Lv3/LnoSBhpI7ipaN4MrtwRc8zZKCu
pfzHgegH2DZ1xA60nrwWcdYnVQZhu4TGJ85dnuUu1G50z8pZLg7JiF+mkEQ0oNcP
WNg6iMgVAMZKyeUVMVay0iyuaXtpwE7OhyR870qWuAgoheVHbXvHyEsbTTKGOOi7
+2YXvcsl4XaT7PL0CH8xLNDyeKOvcDcUqwYjuArc2lI769UR/hMh0fSvkKzCgaab
Bykj8jUgsF5Y1rOPFjBKZ4rKtC5MUcKfXiOHXa6Mel6UOdhko8IPGtJxW9TnfPy5
V3+nhW0Z1LTSaeJshl/9LK9S39hS98iRXbPSUC5Pi/MOPFPi050zMvZBFIA01UkU
NVo+Fk2MbNwURMwDXyE771mHhVv3EQFoUH32xM1iTkkFXpuCfgL6GBO04RJUt3Jn
8zYuh1/2tlyjk8Njhy7stx9JZxCptAjrM073Nl5VJET0D9gj2b9fG/2jRU+xx/M8
KMyD56WISVO3LcceMOeBUvBNvvxeBWAImQPaY7hUVM0SeKejLMhLf2eM2SxMgHSk
fdkxa8rM1BD0uAj+7PX6PsW70ZCHOddZfR7ZiZFtRbapFZQN557hT3ySG0KQ3U8t
matSGYyZOCJCeshWR9vOM4FZ9+qqxqNffnE2alHMDAhtjRYNAIxLlfPTr6VkF7kn
/W7GGEF3C4+YK8145zA1lXIlg+14bbGok50c6T0pAbPqIyQq9kNmNRy24/ZR08W2
NwdREJiO5wX6AtZd4zJVE7B6T9aGknIf015Kn2n/dXyK4V5dF4eB3fq752ThYG7A
eYz41xXNw0zjtRYcvKsf/oOG3GIcg1j7zXicaVvMFjD1fJjqON+fvHv3SY72NnWi
2fdV71OHJMOCNkr2RmUCjc4EPl4aU02wbVX0YiGFnpgT9d4O+o9SBSujxq74Xqfu
A2zbabL/qWCyOKn7sOuD9MXV5HBWJ3+pmQlu+0I+6m/kTxQDEnn+9w25JlIXnY4z
HLmI42TtuTVy/a+VSW2LOnaYwKcoWmpA3Q+L1NLy/LM=
`protect end_protected