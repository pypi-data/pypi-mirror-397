`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQMPUn8hJ5NkADzHaDE1+rduM28Kwh7fIX7p+IY5hPIlO
lgZBKcJz53aax+uDhrV6hxvMiGntSEi5HH+Pr2dU8G5K+ty1FjYBkBR4QdMw7/xm
abatbMIhuDysmmAyYOR82SYb6Kt9IE/CmhYkO9W3Q/KxUp4KpXBw0rq0pXfJx2KR
ZaxaOZpO9UWqQxNmMjxls1pElXEd5/5tTlSLiENn7tXzSm0rRPjJuWOJwzkg2Xue
VmolBpaohx38odf2N0m9RDv14I+krlAgOaoLt3BG1wkYynuJcS3mdICDd9ukNf9u
qbeOjfL69yOGyWcl3XSQts4xZv52a77d7WDdu/9Tm0Gr6iqG/g/HMa7oIf/X32T/
b8H6z3orSDHgE/MzLJkPESDLHEBnMr/Dj/sbg7M8zxJPoWnM/k19NYx8Eua5Bhb/
FJ5MNlIm+ZSv+t/3alWcPHQP4Y1yD2TXJks68IK2RPwoph0fheZAk0nAm+xZzskx
MwuwUOesgVgo5Pxhyb/xfD8PAbi/mROWZkpHV6KWkzO3Gz0nF+tiLhwBfLob+rYo
6k1VubLoIx8gMH6vN3UGzsCgmkodWRyoZyuvl/O5DZCrAkYCsLwfEY2eJ/5JpjmP
xYYxJ85wtJwK6+gdUiP94qDWneoGL6MzEfuFwhPx/6KDm+32kQuYTMPv6qI/zGai
HKWhWOep+KovaDhlG5bdt0eZxmLtdPsoRh/4FaIwUnPL0OE6gnRUOLT/iGbJPlcy
MCVPEV6dwG/EgSxzGotDDJZS8s2aPzQxjbVRoiX3zzgnyCHmZyQi+Op57bzebpVz
vn4/7T3tKPFXiK6VFLPSKL6ogBppFZ0WlC8AEUbFdRuDsUDKuTyP/r/JN7fVrAW/
uyR4awjuBAkOzI6in5+YvJLnGJYeUeMfm/CGe7WFpx+5yBa/2Tj2Xd/hOgjOx5bP
vzVHnn4ZsAV9HHSJAOHs+UEYC5tY2zbLLqSlbvHN7jayjIPM6g3SXshNYLb0sRTq
N6ZH7sKM/wr1eQLT1KNBQMrE0CnGzO9osH2blW2OR96/3SDpz6BKKKUYsE1aCzUI
h1Naef2uwzS7vedPtV9+sHWcFQJUTFlCJpQ4xQnhjEhFlpn5C5mEnBhENwMzS7ba
3M/mbVn9T4K2lzWlLK6/urLZ9PTiBz05rqI1DyGM61TS77O2fO8epT5Mk8Wqy1da
0YFq5Qke8zfePqZ0jBjhelCBcX5lo6fxLGlZREu6Yvk5oXnR9eyyWgXHe+dAJj7U
yfrxYUgtGiwtvCipDJ6Gh0M3YXcNfBad8eOQUkdvDFmfhBorl3RFyOc2/yivpmrB
ZBjrG5vxUt94wcoWNqL97jCMMoFRgvVA+TeU5ixnIGFd4tRUnC9jg88/lKPb0dHg
1u/vCgWoQecx2ZpyTMz3jo9oZnBYytoF2StKfBvd1//ZpQDPVo9XBU4aU4d6svmx
gFPztrsWIRyHjNH2lPdpzCdBKHVIgiTw/V4gd2YzFbKb35Bd0xtcTJxWcbtwxODj
l0g19ZkHh3+MRtjNJwfkgil2ETMq+hhUIY6VqGFEWojFwrEysT/HfoGauR8yNnno
vlWMPxw4OJlpSmwWyQeIkrgf6UwqAxQhbfn5ZFn8+QuAMEf7/MlNEF152RYMVvaI
bq7mttFuVldVhT2yyAFOaQDODqemwMIOi18PfMVfL6BEx/h/PuCXfEmiEFG+l8rk
3pfoGJmiTZ/JXDCfehGvnZuKLwQP3tpAZUB5BFvTQgsPsXy2N2wPH3kmtxnS/6BD
tH2in/bQtuFrXF8sYsQF+B10dkVretykGSJ+zFmjiItklZU+sPMeDow6g7gY9ZXg
Y5yw++oxFy3I+Fs6oTnFyQAvT2vqJ+Z4aPghhimN5m1CixQ0BgoCn76tgwOJfAeU
MF2oDiCGWPj5iTcjVpAgGs669SjL7K1iOWEJkOvSGUN8ZBfT2hhxpbhgh8TMUTZM
qshwZPTpwNfd8v0u51SQ+cVzCc0pjw6PmJFZG/yi7fnG8oaHm6iplFi0Dot/K7Zo
eapUcAe8qSxRCmjQh0PYaEkR4OA/pxF2okVQKRCfsONaqjNa8koY+Gw0abd+9HUO
m0yeYU0wT5SgQe/NQ6qcgZ8HfqX5wC3o2l9v3ZswFtyIe9puWqSBRTAKfF9j0bJf
+cvLIf1LuJTj0H8TgGcX/v9ws3CnxHxw7DffnwIgpmGna6MJiQCK5f07BqKul9kQ
r3L1HUJzJDJuNeILsHVYtN6bp5G/uAKi755WDzSZXCRXeheUNrMbnQag1RK9Jxwv
6NuyPi28/3fGcURr46bSjkHL8ypNoIsoh54ddiE7DIfd2k7qwpPd2FhM8jDY1dRx
KX5GEvqwgJkMPESaKOrhzZFYHhzWmOH4gsS9n4wwenqIR3qrgMhE2ssQ5WllzlLa
bpHSkxUJZUMUm4MQX8QFICxe+d13/cxE88f992QU26n7vLe98wxnvL7KjRvGGEjT
C+pyhz1Q6rqt8yuaUdOv1oAq/+Kp2faLW/tPiH6xEeWh36MDlN4SnJzKpq6Li757
s8phCfvL6kD9sqIwLWRImHqdXOHWobfuN1qH22QCROX6szX2EQmrVrR9m9OEwqKX
aLnEr0xH9734PSvg6QzS+wo208r4IHkPZjIZ4A7RY4EVL/SzttlNlo5o1HfPR+TJ
0+ea41g8lVQsdvYowEvLTaJQhMzoPe2Bl6Kp+8hoh3bqbJPajKfO3sOejKrVYQ+7
Jl0oPiKPxjYviIGfO5eCl2o+CiemM8JbyWKe/BdHd9/tSU4kpVDG1DRVy9OBB+KB
Dtkt0kP1w2tUcp9tD3EBdG7zIoTrjTmlWgC7hvbCbLOT/BDBrb4lamKNrDWWhBIA
pTmRGPbM4hjNCvZMF6/sOOJ3DQu/GTfGwc1eq79J/3n7ryuyxcj2/1hGM4qI10XI
eZunm4E56XM1fwlrl1XrcLV3W3pPBS36CWkMuBiD9Qr4uWu1jauNL+BkHwgsiOfX
CxQVc0jWbWmP7L2nD0b0CsaS+g6BZYmPMoVNI60q3MuoRX2p6/Gp+yI3OBsryYrl
1+ffYpJXjFYpH1TYL8U4vEXhkGMH2ofENz/TzOyUUS+EvLRFTDAXLANoJ26LrgRW
eLnsUt3LR9J4HBIDy/xrBn5QDb7huvkwIx1L0dVurLkv/z9ZPrRxbQkfDdJFrwUP
y78sHosvz7OmrGqIm6pAEuad61A405z3AslT1ZP28r9S8JXyVs/cy3L5UDDigUAY
XHmxpbQ13gKzMYQHSWttyW/EDhhKIZ1PGgpfLNcZSXUotXqNbIkALm3naJ7+H0fc
S0Z0z13s0qqlApHaev3P4Ji4Jtpv1ye4WknU4Yhb0MCHqvvAo5MGcJ7tXBfSoYan
WK3AoY+0qVM1MRbOLNmESYzyapl6eQoZFtnPB3lsMS68K8mC+P2sklPWykNrvv9D
O5QGJ3doJ62jqp4uNRi5pB9pu42bupMLKHw6rsM3OiYGiJY8EFIiYIe+umX6k462
gRPcpG/chSv47m3pbqmxzLF06xS9+0AW4RlVDCCscQcdw5z/Wc43zReU3vc7F5u6
HbkUUYfFER3Oisd31asop7aqeHtFBZ59zTHSzON6rROdA5xK/XRqRNp2lWZU5Dij
1N5ri1sjn1WqMtCYTqaXizGKLhmj2w0yJ9/dApR+7V0sdEgUELedNP+7G5DqnViu
Y3md/97bYz2s5/kVj0a8OfDlRJnvznOrBoDTzFds/0esR7rNVVQ22e1hH2UpJczW
2Ep/j/Kb6NYk/Y9p6zAwnkSb9JrWmstXHsGh+1W2z05Di08l5AeyL16PEfNvXcvJ
AV7ksPDT01iw8QtCL/ZAU9XfBY54juX5bAoCS22HQDqejorMEBbpNXlZFN744dOL
rz7ADYQplXU16NIqSlYccdN/Ssc3UNwJ9NQ7HEnCYpafkHODR++a4aYL+BMBNgXN
Oi9V3UvQrIX4LvOYPyJdx/1XcN3GO7R8pc4sU1oD3asTLk31G7V52bSFcsDjI0d/
PUpxMuPi9/Sn6pA/kp8QTh3ujGje/eLLKP85CyZluR4DoksvaiDmMBv8Qufsa6I1
gtynM+teAgIj7zUExiM0q80t4VlmegW8ObxcWEDzJxy38k9z08gr0DFwIvRYkQfS
HY9CwymrCzLPQuV6i4DFDNulChDagrDlrqvUDLDJI6OXLDGOsUqzt8IIpWZFapZ6
ipIHbdNixWLmNenmsT9objQUcRrmnj864mBm+YTfdUyFxGRrbqmojqRoOH5Cd3pA
JoDtUhRq0yEc2UklLUrPuTF9BYOqqBoE1Kf27CteROrU1ojRUqp5l0j3WjR6HI/0
IwREMZplQwxXdnmMAt+1140pAJdfRiV+syOX28bSmwdsp+LEOXq/g12gDLOmILGN
cWsFUCh3ZwTxJLkCc4BN9vQmTcMsQ1irkR3cnWpBTP4UP+9drmyEC8F3Pl9aXYi2
FZcx1dTna/JzWKdRkzHzU23D276rh79ajvQvKZQVb0TD3WHo28dEXjyfcKtCGxsv
JRaDRm43gLJjyYYQR/zOWUFKmbvrNPgCgnSO80ecL7Tc33wKgobbxUCQFroyDrtu
4og7mQ08vdrJDncL4e6jtL0UX5ySFDce3rA07UOSTyl5FOsr8YldZAOom2ysn0Vu
Wtf53YMnfix4luchOsX5tpwdVpOClLI5/7Pr4dhr8SAkgTq3z78pL6zlTDOz7R2s
eEFQS2qBgjH5ru1Xbe2D3PBhFO2B+KI5S8whsfP3uMZIoTUfgTyXbOMp7k7V9xBh
3rj6XInH86ytWQK3pUeTXNfQaXJn7t6emBoepNyYMpfWcMLU5VzJ1ErYkKfsqAOB
OPrV2oxgnj7CjbQncAj/0xJy4v6xe0UIQW2k7WbAl5KpSOZS3NdI5tDK4+63p54F
EamIypoZ28YUBJOLO/zZbjFtezWtroAVSjjc/325USs0fiddrizEiKTgj1NFKoRC
4c2XxMGFF/wsXVh1QbmKNBHKEhpp4gHIb2qPyat0zjakcsC5H6Euy9v7QLhvylA7
2WZPjF5s1LvY1SqCmRb38acxGYNHVxUrkFc/HjcB3mK6Pgk0psDbwTX/cnLkw1TO
161dAVverKRFe2h427BhjZGKzkRhd89Db2midbKFzN0TdHngmDFfT1wZEA2oPmz3
b7c6Hx+AgwNRthLHaZNtsPq8NXb+T7h+N45JIR0eBzk2IqoAi/KlOFwIxud3CDiG
ug++8TtP/pj4fv6VyLV3lJwhhoHy7Jesfveoc4JWCZBk1/NyyUhGcmO+nsp4k1Yf
uQszNNuIEhiiAXFW4XKuKUbrOVoGLaMxi/wo8ejOabb5q4KZ4HCpTnrazjcT+As0
POYYNgLbQwBuovwkURvC3XidM4ZLXoUmat9kS7JCHg+EQ9nNMQGvS7C3vDfS96Ss
sr6ynxCZArlY20WhNz4rhDH+optEi8JAJliXVwwE2zNFQ/026JYvjpeX6V16BB/Z
Ex9+3dwYvDxIKLvPggSqtSBjeGyF5TY4NoX4VdFnPk6bMVPxiNa/rJ0sor5cAgXA
GJzOr2Kp7PAWCARDUPo0YfV+gmz5J5yY0n9ND60QTl9FGJkneL7tnYKEzDvY9jLG
mEguNWuFjYup1wpTGkGlAC84J4FnYZD7duIhZ8vMdp07TLaYXLs7Tqkp+qRGy/WD
WrL63KgyiHGQLesD4KvD0xioztbA+0tus+lUOqQS7YCO4ALFqD5sZoJLid79WHZU
sLcuEzlVMd4fme4iqmICI5e9jOLoqGGIYW5xQLQf0dvyk402yIKJDAbtkpYySY/z
quyQs/gqjEyjYs3PHLcCWbbC+NTGPz1NJxTBncVVlP8lMQcPq+7iHdY/tbjb1Jz+
I3zQjJGkpay5LRxuVKo5MN2MgoH0j5eAnFb80hHOSDY/VgPbhYEaW8ZSZf96k4oq
fs/LRsslwiNjcCXTXwIN1y9l04ICJv1TW7DSrW2upnqUIz0XdFfdeZ/bw9N/fbQD
Idn+7Lt3G3T2Drp7VcP1csQV3Kx0nQ9Jwk97tFD120iw5TBCKOS4mOdEYrBjVHE9
5c5m7RCDjTZ1M/bShC1BBfUyPatr7oaE7biVHduejxLYV4JIZ0xPQOzsLhZVtg8m
dBcwyHaIoDxEHmQrFTyjIguWgvnhbmqF5m5kuv3Bk+1ULVlT4MbPJfjYx7E+JZXf
WYri8ht8MHob64/OygIAIr03dUyxw8g7cdv4FBeJNhglckcre4Tt8vgASEMQVCdF
T4pafOH1BKEbEIFTlVmIOndzC4aqytP4uER4tlMmf2j7iIRg6J1cLcuML0sEwdOD
6sctQBQefv+mjJ7TfKAd1e+GxPH9VVs5415UCIST6nwQo/sHlZZrZhhCzqvWtJ/H
t453pIcQ2QyAro63EvS6Zp1xgs7Y8bE9Q0IGubnk8yeMJsJowUX3U/+CAFl/vd6Q
QjHHzWclmXeIbQCr/tRiF2YZrf2+7E2xk0vBAKQ15ZmmbXGAOsuLrmFXTiGmSjs5
KQnMvU68JhSDrKgGGYCg3dsqVM3nEbFzOGr8dxpqiBeXquW+YcrYOgGVt6EeVydG
XtlsuNXp3WVxfpMkkbR1B2s3nwI2NcxSipsEqkGhsDMU1IHbxv/nXUMRndShRoW5
iDXP0Oaqj6p5v9oT+mK442TmUkL0vLUhz0i+Jn58ImRb+NWBsfY001PlN6G6m+9q
0ePrV7DEnC0Z9KQkkM8zd2hQVTnK3ogEhrH0T7IDbxGGJ7JyijAFIeA4IStmRFGL
g8xpcqK6zrJCPhlABfpl/T47joCdIHzID3HF+OJzpsthERn9pZgjiJfFUimIUjTu
neq3+AP+u+B5Sd0LuslNZUii2KtgKTCwCpmueQjbiGklBQ7D+2vqeImjiQ1EpWPw
J+OntrtvLVeNCbOxWSDmmA1LsqAJXb4MaJ83QoLqno3DfoGOJSsjR1CFH7KtL2f6
i1fYPoqC3B1f/aeWyC6OIWxLWfqsEVNWLddBGU+kpf455rhA0eCMTYl5P3Wgko18
kzHJGOdqfKHBPYblTAVhtSXXooowwhi6sqY1PVZzjKYQr+U482FgdZJzniUFA+pm
SSeHUh1dtbbg5zqTerRmd+3YKPy5VVgPIQvjx4wjTYnQGfRSpAhZxzDCPF8tQ4f1
SZXOdUgFvM+wkX3Z/tfqR99ZX2+4rJ6p6D4JdFi6fBpRXkmd9RgRRscNhKUXtv62
UiggIXW5PG+tVHqeVyC12JIgv2yIPzdfDLCjoVEZPlBpmzdk0yfBlxpg0k6qDXyV
ODKvMa1OA7WgxV7oMqNrKRZLbxIKzfRz6Aup70u6NOR4T4plJ/lfPFHyAwCcGCD/
K+fp8KCov8V2KG2/CtjYQBzUJhUF5pzQVAyQ8olHrlRf72Cy1sf69v3Kj3lg25Ah
cZW0RwtkL+3qwX7rmEeCvZ/XZ5sY9RAvm79iDJD/EU8XKKjD78b0/y+7Ca95IAlt
MeAj0XNdFfNxSCCEwBFtGxskir6hRnt4Nexp9/kxn+8Fg6yEIWlRv8dmKDQ9f/I3
t7CGfuELMFMDFcYekotHP5jxvQU+xYjpR23Z35at7/NzDtnhZ19HC6taWpwU8mOI
52WJ/VuHb0+baVhatccTwQjNCwp+cx+Yf8eB4lE86WADH/U9Dqqx4JnWj30lOrKj
nFujSzoFDwwh1/gHR+ts+TYcYfzGvCvXYT7mR9bDABAMPpNPi8Ixi5uxB5jsyv01
t6oaX31C9uwKwqaX3maGvFvD9VVucyhL6EdrMx7zh/wFqZaiQ49iI4HqjwHpP1LC
3g0qQ6yzpsWVzw6valAKgD9PTvF+joohb8LRKQZYDEpTFynQqEJ9Nwp5+mhsmCUj
cdhsK4QJLvP6TLn0n3yO0cL7WRK5PQ7trc1/3hdCLq7jvizgEG+uHcT7YI33E6Ag
fTrbPwSG/+dXMKssHxX1aDrPhQnXWQt/m6gvdpAcGW7uH11CbwAAkAmQCAm+e7fs
UOov+gJT35SNV5c+lUr4WpTpM52uFYLs02Dm/YSNtAqFLsqCA9+xqXB51AZ20gKS
UORw6mTk2AHPK8ejk3SkB8/83lspOdFOKJgyAknWoXpjGVb8KyBhWtttPAR2HF9J
AlRwtM+hyr3o9qSkMwaUKOwBbr/XwQw+3UJZCesZRHicVkA52eIc97nFIjhRcH/0
4n9/pQOAEU/ipxX8whfK2rd/7F5UVG21gkQWZlXn2oY=
`protect end_protected