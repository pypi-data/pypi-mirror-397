`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH0obzhlsarOKkTfjzL+TLLh69oyRPv+HNVSwPBFXGdQn
fwYajf63q1yJEK9eypMtfAZj6HxzVQ2rC5sZePeAz/cmQ/AMSxHKzvawwCA4q5z7
0oMNzudDi3wQhdf7tuEj0PJY/uaHaCCOOWrUN36JcZJ3UBzTjg4Uj3QThxATLeQy
gRgWYCPS2fGQfrJIPYvifcfcxum/ccZZGuu6PaZt+kqhbKofamBMLYP3JMHPO29h
G9I3gIzhUldkkE00IWh6zHJXP0Pggb5nERKnxnHWp6o6YpLDmxPNwS06Kk2X6Zp2
5mgQRENNTuimZJ73ITowyDE7LVD+wZuTDumrHW1KzxsQdCPjXJfCvY1slseE9b1x
crWD7g7tJIRw/sp3YixyNh9Aev4cDGIvB3HXOjl3I1L1fw0O1Fz6dAGuBX4ciXfy
mlGRDyJN55TfSg/fdFy60jMuBdXkbcPV8e+jzetsSkqJDC5St1a6HKLtRNw9XX2T
0r2MLvxJjqTx3rg8Pq2t/KVqwBZViNqaXfq+eOJurV0x/t0XSUt0noWdwKEyYEDX
UNd1D6txVClXhIcz/vFhjeppe9iNUqaY5ycQQdGHqTPKqlF6MIirQgU7xB98IraH
MVJ50q1qFTkO2eYtKzdJwlxhO9FuP7ie29RZ356ckDruVl2WcaLfHkZec1YeVVRu
A2AKM424jZ6u4AFT76/9xIK1MHGlgmJOkweH3l6gsekFTmQx5W+oic/VWKF/azXx
meItwOE9NCWSnX59qsqGjyu1j9eq9G8I/aX63LUrmqOZeZOkg7Ou6PY/mypC9oZz
fu0+3e8kxQl7df7PNvyXUwtL+Wfbg6RmtH2+JW/GBSlv8xIP6WHxVWV8KtkcbOJd
fWAFpER66xP/9+sJE8ddvRJUJTcLSlrbqg+CHJRVnPkbEbnxrMuZOkKBKZ0TzJiY
UB2wEAOJzse07YKc2DoAq2YtAXpo08AY8ixfwJTQVAfbkhJ00Je8lkIWwO4XxIQW
NI42kFtRDiGk9O6P3noh7jmMdl1tEoHFFIYEfJyUqv0EeLvRL7HgpMhd9jeOC1Da
rkDiJZo8+TKyuPNQiQYyDM0g56OYUwDUv5IwxHOcVoXURV1NNrIja5hIeI8L6q2g
pyVIAH9JCpFGB28kTgON+6fU6gyXSrB7LKME+7P8c/s/5cEq/MA6sbO2hHBp588C
sw1zKaa1t5zi9XkZ+pXQqw/gXKkcjy4wy3HM+HpA5WYoP+H7NpHPctuCA2owiwR8
ngduLtEndTmYIxP8Nb99FKDkIUIe2OQgFBjyIXvDdVPwsdfsH1em2EARYGvU/irY
p+hoe11+33+3p8ZtwDb61Mxg7XE6QxHmwUfxksouh0FkJyjQDiEXi4OxqUb3m/+X
fwzHgyEQ6h+JoHuw4LLKafhjBTQg6JhXiN00y6JJoaLnui3iA8q39/RP+9amzA+E
ixXO4YaSTBBzLB5TFjqIBcZkJyJuwYLoi5X2i+VmXRhQ1OtHpwyG1TzLPJhOI37g
ueh/AggYwYCOcoKpSYdhHjTJvZ1LBy4KIuco6+2X1NVYSYDqE+zyxGGQDNJNUTlo
FKqSBskctQ8Cn/wPvPMUmUclZJw262MYxuVvGZA5YHGjhjoYx/niv5z0Cv20D2wj
+R18HqIrt9h3QSzF3bmoFL+V2J2+oer3M8Uks0uBxKS/jlRB5NKBdSN8rMMuODDq
YBOhgm+7Fjv6NF4UFGDFMZ8V3ZoJJ9cYI2KpEu/MR0FKCCD6ZR3vDxW98TFEQp1A
qo6g9TISwkh5lmkKPyqdgxEltneL3HQW6Fv/UvpsP9KM2ypRDU4CENkfRDY6lERe
rPSBJJNWv7UHKf1K3MElZZnJe/bMBbCltsQ59v7pNTHd3VD0uprnKLadCTFz+1NK
DGaV6hP0ABt7ZlbstA8TUcTirZ5PrejqI2rLOgr7AJ32F7SBlaPb2nrZLT+MqRNC
V3RUkleY+Ffn8hc/E8em0cLkt6feG6W4pbEj+TCIwvYS+n87yJuzBL6MRFqsSbtM
WUZhg/6rcDd91qfNxV/5xrT2LVrQK7ZH7Hl6k3sE3okCPlsgbz7jw9dePddqs5q0
4rFQ74nmNCBynH5aHG1vDPbpT3mM16QDDgQEgBjpCiiGPe82qggLNQoBvGrH15iS
nPmrSu9BVV5XzQgLIGRfa1yAhnSuAvYey+EKt931XT/cizMLsL/2TjXSxTZGYKDe
GaB6uaYjQNYaMAT3M4FD3nJhD0fZ8blKTb7jSDSG1/1SMtjnSjHQCgqmksSK79Mz
HMkraGzMhUiuFLxxeO4O02H0x1s1HUXBRr3AMVW/CmYMUoGlIgRAh/obOL26S7/a
Oa0hKUDC8hCyh69S8fsmVL1IPRQxaxW/OIz3YkaRQmuwmtlnmfM9TjDNcGpgwb5G
TIqRErRDsjkffyrTD5BoUTh7KrxIkqm3HrD03hGuDUHEcoFdVAg9+QQQqn/FWGDY
R9U3vuc0sumMfijF8rT1Q+N9wgPNsXBOJn//xijjXIUOPs0ym54SZnOg6Gds3TdY
IVH0nlZL1xUzKL5d+LEXTQ8zQyksAeAn+s739Xkv/3InFDREDnSflKY4OA6VZP0t
KLfDkvbl3PtLd6f3uP2/LtuWLvsWKGD32yK0JXmQaQx2JZ/lv4TbRql/gyg/Tcor
JLcpxK3vK+Uh0VdJfKURwU6QC23eSieurfU6sMz/bx4ZPA02XWPa7dt0DAL8piZ+
KmqBRf4hbk22QsIjScqQE0tCvQR5B1vyReE4/L8YY+r7NmZFmPDKdkHnMaWLQrra
8C8BeLIm6sEU8Ep256wiB8i4XNnVryq8idSoorS8VqyDqNdGTkLD1ca2lccfVUJ1
+60f0DDGDAiWDrCHjF9gU/uzZspPxZ6SD7ABlMXwzr+qW829mERpIuun89OsPm7q
WUtZZ4m1Wawk8x7HuOYPxQHZWYn1KDUNwTy1l9CJXQhd0lXEj1Dr54EnXUfYkihh
zlJyABSFnUrizinG215tmZcpowu+O5UJJ/bVSz2cwjcSOcayBSq14UvZmPlsM4kF
Pp0BDAJWJUFQ2b8thskx15cSn80q5IKuzhHBXb/FWy8NcuBjzSb1/zljlUqQqcSg
Ggwf6j9GXN6dIQ4+xTrjZxAlmz97XM2Vkh610ZMzFzLvvACDvBB2vrKw71TXiD4G
LYyWJOmiSXHTtGw1dcxOOohx6TQ65h3nSYFZTLdJBzyA8F8pmqoTYJ6navPiey1N
G/AdrOArnWS3M7ePJhJ2ADSN6I6PblENgna8CbfMJKGxAUgXDFTkdRpN024yfNEq
wv8COFZymY8RzBdBpAMmhgX3DzTEO62hvFTqh2pdnTtDCUbmwDDSnwX2sRp8U3KN
QetJPQMDgjFUvJC+ExaU2R3be6ehtRK+FpLnignVzUhainFcBe6rOAbH9YbHMck8
/Xfy3JcSKYFLLfbPVbZp/36rdQSh0HUMg2NmbnVUyYjjMp/xkwTMwayje46/pMNr
gWzAZy6wgZwNP3l28IkXE0I94mqoo0X6cV+5eJSGYRy+qaTDuY3LvYGGwuSejS9l
TNEU749Xvzis/2AzM9A10FqG9icXG+Aq9Kq4IBANNK/RNC4QB+f8+gJ3UYmvpjFn
4Xdr1KTGKIri8AYRZFIKpBPEsTV9ZEHQ6RaBHBspycSiIJTKREckgO40ZpacBynI
F4gwhMHfs8eEsVbWDHjsVrMaBcXw5mNduExjhdtOGhNcWOv+g3SkNLzxTOiDeoeF
jTJP/Ck5VUws8VJl+aQ2WHIUrFYKG7wCBGUouh33I9dZNJExdnQgPthLm/OeqvpU
z36eZwoYET58Df29NduQYdEkLXem0fnh99NFvfJ5giJCCOS0RiKaO3fkHY19wsRz
mpjKvrDCgGkanJJuy6pLHwPF0uzDvl65BNzjOkhoaOTTR9M70q9MSWQe5nnC8RwJ
jCnzUSpw57D48fTFT97RrUYRbilWl69+bWBxPUyXtA2ZPxx/0cQpt+8MVe9UNi0N
41JFL49wgj8tNNAASWvH695ATGIGdWKwXuu3wtT7A64TmYUFDbIfylIQM2ozuoY+
tGBnwegVcwsP80GMi04W/nXR7w41GyZj6JEBZZbyOkPBl7ft+DxePvrX9DLNSgTu
RwU+Ev/qM3RRtamUBMPQsZ7NX44l0av+85m9bkekkz03o7vn1uRtabESVIwxzoeB
y/Ae1kDn53Btf8IgamJIa1VrEo0QkIrFdazBZfkfmA76+VYwM+blY+pmUxZz4YPo
tdhARv6FSWmqkRlkJjuq44F8mfHQ7kMh1vKFyZpt8ptJ+WO34Tkt8CyzPxTE9s6F
t2crnaD4/AZZblf7ygwMYhS5u/vaPNDP616/H1beePhpflmgK4hG3junObcnc1jg
G+vpXbPzz2gnyENgIcruxybRe5po8jBWhHIFLeqiGrUEhxLxpMq18y6t+Rj6gVGv
5x4IzBJACzOOwrl81Y64EKHZBgOSjKrtqRXGFnSYvrK/qufBd/scPGCNxeKoTF82
n/lYFfAHF71viA/SCWMMEZ1/0aN7K3DdKp9BQlVYo5+Q/GZEJ4Wn0kIgNaYpMHbn
XrANzlR+74G/OdZuHeGotrhCogSCyS4IJFpcXY6joFbespEI2hYIe8uxHnrSVJTT
3cyEmHQQ/ZG1ponX7yMZ09Z9yfmYZRNP9oTsNXRkbCRjLgJeFthWVPQhJyaRzcIi
zp5R6Aykp+76S3K+g0T1LrMlqAFh6OSnFwFrH+onRi10FQg2/r6nN5VJLihvpciT
S6JE9t/yFjnq0nd4Rqd5Pu3UjVWS4elFRvdhhGoQmv3WWmMhuQwShbcTdnVK4rL/
wzIM0rd7weepv+pfMfpZ0llglEbnV9NY3HWps3BXp1bTfhkMBYJUhsY+/t0dcXdE
eeSWQoDTsUrg1/ws+6tuFQlEDDm2y7YlEn2UPOc8SO0vu2WULOxuawNtNXF6Vb+o
h9tnNacp8K+R/bLqoujUH1Ys1gJCAMDdG3Z1Iw4Z3zpYQuxpNupUQ+xGLKlNIb5/
udrEo1WH9+K5X7CDNxtxqwQC4WHM7Z77b5Arq4nDNSv0Pp3//By3iqbrWDNdhnGB
ZDwTR4LufnHmSAOBarAER6uv4j9XWainBM4+oAzu1fe29QOMxviduYe7VjuXH35w
yr75MQwzoRZhCxWtwtD40zQwszhFlakfjfiFdfdpq4pDEXfLKAIK53vuDt+2B/qG
ZUxpdIF//p3bC+400c34qq3buEVoEDpVEZJA3DSCtMydskcr+/1XpdiAnyj/zfnH
EX+7WoCUrfgQIqGdh2Kej8+KdronlYH49kqamK7pnkQGb/ZcHGudng8eOrWOcCy1
wDL9mmZCYWJ2ucLC38acnSlF2O2o4EFpa5utwHd4Wk0j3WYHcs1UNHozJQohAFcc
SH+JnoE8QhFG2zoo2TSkeoroBsZa00jHLNguXn9uuRRarmG0UsheISIoHqKPEs90
fXABHTbJVWGJpNLCsXO7mjo851dcG8ZpsUtOUI7TnrDNcaEdOT4QWn5Jd6dC+7TB
/PDs3ByNvVu8JlsxS52kAgn1POf88QEOTMokZB3RpUhadKlZtUF/b3joTQj3Ml25
uahgQze10+XNndy2h5g2HrqCnsncDsRyl1e/G6VRslh+2oim3n4NDz2FIZNZ6J0Y
/n7r1hHPQ1ZCm3A3DEKHsuaWm1O/QvmZsjSekiGE/jq/2RAbrDCMlrmr1TaUi642
Orp/wlzLbpBhxSHa0tGbn2oJsHfepMaIUAP7sVqYSKYtFxtOUt77mEHoOFvgsaCp
0ZI+4rWdFoNhuKTx9Na9FRknAQpAHw040DXoNAuM5kgunHWDKtj5X7EUrPrQihYo
ekaX5U9aY3V8Yfp6IVBdbFpdViXeAm+eijAlvBxAZINae76I3FYMob/n7RApOoQo
CKJN6pYY/7SBHNCvv4A2lwesc1MkJu7Ma+X13HIIJEM7B1m7J36ppGqCdK+QRWqB
dmwl4D0qiUMC+FwcI/35XMnGrDy1X6VKcYEYj29Khj0zTTzgZ6gkSx2aI/Bzi7+g
gtcwz9OKagDNYIi/AwzaB+0yGdgwnrSGL0X4OqKz6CsvuRnZ1To2FzCkKKLFSHpU
TerEZ2j04o0SJd2ZZ8CyTzMPm+xHh9X+LqDuJiEL/n+9YLDLNAKOH3bTxX1Gu9b/
lPWos15q5ZXU6MHH/sSYUxEDEY7ofEHO9OgkXwHYGPsZi3Jz8u2nKqRdXK7YEHDK
ABV91G1dBJsAE6ztB3fZnOCXDHStVxmqZIYHhiz534K3IjglM/L5rKXf30a+YiQ3
6r2XyXqntDTSsZNffA/TZQaNM6vsCWLLGS8aXManBMQY6HKUe8oqGWBZnBv6CfuP
UX2eJtHXS5RhZbxkgaWDykEpOqSaUlHA5Bgy3C9RVUNE4f3RtQ43B36HYofg5AuM
sCikml5n4ZmFPfhUieQ9funQfzLgBNpx7COIuLf08LFoSsQxjYr2z1WvvJC9mwcQ
CLmFjYAQuozRyDmm43B7yTIEFfGhwM/FpSHBFHwmWXRJiWsBpd4D0/F5vbfb5WC8
BRS15GB9C7OzNQPBQ0GsVvT7kOnJi6uofyFzpwAtqyGmq6IOaOufzKbmNhd1auTP
8H74ZdfI3UfIzXOmz8hqhJ8WOG6t8k9LjrfPvo1zR9PGSnoue1o7Tk9bepBog7Fc
rDYibPYYCtC8Fomrr7RMdRqCUQZsCgeYk2bmXPMxabLIg29rjjtFM5p0VqSlF8GN
pnCMBJSPVr3Urg9E7eOw9rLBeG7SznNuuCmF4HTBm9ITqs7EOA57t45BM0z8J0jO
p7A0cGRBMmcP7q4GbnD99gm+UwD5IFp643+zMpax9HBBpb6Mf0MmyVT21Rd6hBqF
PSJwGEtgDkJ/yqpO/ecRrzWagux9v3X+PJjBr9T7p64SC1hO6qht4lwF7DccBAmK
xUg5m0nAY1x7ZFNLfypg11e3b5/WmxTPW8m/0ZeVHr8nhL62dNSyPHCRz4sohiuK
8KcpHYqKbxxOGUD/NkKwSG4KI/uT2gJJkImpfHxq1SrNkydvb7bdqLpbF9nP2V+Z
ofOYiBzCtRYRi11fR3wGK3058eX2Wb7KtFE4Q5/Mu8s1osVC2TETmj+PguHs3CBm
CmHHQNU/zlN9OiAXqn9jslUZvcvaVZE+zDFDUgriNkT3OFtB3slz7MhUk6aYV971
OTtzDqzbELGMBTLKwjVdmaF8JxOdRKFTWJ7Cqj6M6DpEjnD6XZoaMs+ejUwc1ea5
xCC6GmwE/cb2Ab3ilnxFAoZoPjixWFrq2j8bJ1vfpDnJ870GJEMCuppKEBxwNKlC
d9ZGsgJ5ERtRR00dJiE0wiDlsTZSogRZWWQQJBpmnup/iosbn8LJxL/baBcS478N
NgB3U6uzT/A8BBGSjf99RR2nKl6rWJtNHkuGnJiUkZzew85qn4bdPaRJ6WzSTxjR
wmFtVtI+9Hht82Q3TTwJ0oDq/7ykEwA8n1v8Vk28gTFrCB0pR/OjLdRqBl3gjrfs
wVVzuMp12HnaPAhge1A26zo7LhWqrdyxtB1Ed4/BUejckAzT7YZtXVtH3Ocfih35
n2HBTgCJ7OItQzkvSp6Aa4GFTzQVbYXRgoP3HhXIkZdouWuUwy6PH/Wb4W7wq1Na
T1k0JxZbpNA561HrJ29c/Rq/kPirQce9E8V4SJaabyFACmP5i8gN+Pf6NqRfGvcn
j1i4UMiVDLoiy8W3rIQRaJ7e/GSSwi3QFMj1U6yzge8EtyWhV9jDUZ/M03pGlaFl
1mLb7QEyBotcHIL5WSbcMG8dp/HdIYKbTNgx/SAe3XJtA/B8M9aKCNQqNkmD/8e0
51J7+l/Woa+cEeAKokMc9IAcSrLS46OHLi3IhzwS/jqg/O3gP3DXSflI2YBsaSZj
RiBIPdC+g+QqUnAc+SPv2jMXG/2XzpjSxPtv8Bpy4qmG4MWjnegQjSGyw0JOWXZA
OVFoYgXDb47VDuYkxMPvj0GqxcK3ryVHNxPWHvuMo4C4bbleSngdOe1AHpZbcJkw
brljAXH1ZtwdzArJ1IGlB9Hv7+ccnZ0XGwuEoP7CCqZWwJ8meCxWrRzg0vpRX7U2
PcasBbkucFEUNEpPx2gXQncteT+j87B0+BE5gjwwB0DVlBqDnP6nDiaV9AALAzfz
dizbATw8GJ9Fj5pozPvfzON998hbQ3D3tKJzV1iWCYMGUHM8TXJf3JPfy78n7r2N
olfiI5z3PiJqmCNlCWZlCJWJlIRVsml+C4VrHmTMl5sDBlIk67EQGdykhrf9F8W2
j/mMGK3EyfrhbmTXR2Lg3KC2knznQZTacdlNIxL2UlPH6Mngb7KzUIz/4vuFsq7B
0TBH5hsCnEzie7neN/pwZOgrEGcyqZYEYStdZ/SxB88WSvgh8D+O5+wk7ONmDh07
u6Tc7JEAsm9/we1LQ34F/caMwrsaU6lTSdYiZh5bGUk8hnNuegkONepbNSUoMJjo
E7JR9WLUbVtep4cW4h8DIw/B0XOI6pAn3azVwp47NICCoNNreMXar+/LwD5cwfrU
p1HpL7X4CjkIXWYae1RkO52xPZjJxm79t5e2py3QShYNVeeT9VRhw1Ia3JBHZQyL
/7UD5L0/5GI+FRrmQlkHb+uPNlRHAUwvJ3ANn0o3VImEwWMDIXIhEEVn3appXcmY
DvEVcJG1MxzAjQB/2ieTXEn5K9cf33LQ587zFhTtbbJONJcO1oW0w88sxpdzPDWQ
uhH68+ubWcGXIYS/MSWXqJOYWM/aRfSYH4Tq9a1Izy/GqhcxmddJ/eNbL1etSP3g
hFlD36i+DhW44kCliC9mVvLj/JyHdLrEXyiKFxh24OtNbZVJsNwt8U4yrwl9k55b
ruZiIHFCGV+2P30cmJtitNyFpru83xpUkGJD7vqx404mHS2W9KtQapvCTZh1dp1a
WhYQNPWv2Q+FmvDKQqnDQZViomn1BwLJURkMD/Fn32gThfZhJpNqyNGnvYwfXkNR
SCrUb86tb4SN+u4Cbh3PNcl+T9jEemtZKtHq09RFSj8t361fHbruee17ldaM0tks
qngNa+jc5+PGSsKAK0sP9fReZIijyDQTe4Ejjgd6q3V4fIaUQJXromjcmQWQXVYG
nFVl9OOR3VS0jqTxVFbbztG9V7Wqpc0NQk3k0sShQcwN66vsQbrLNQ0T/UBjWAj3
LXag1aO1Jr+Uk5VeXVGIxq86mJdHWGrBZAqaCSOflGY5/YTB70W36SxnW3sZlJWC
G87zE/bKmQ0+pr0YC2GFxNYD5H2e9S79jr5u2+8qs1RvRrqu6i8ShmFXBHwzop/C
WoQK1nd4r0TCcnqBSMr23BUv2cTFj6upi3CDiDVJqkofHKgaTxzrT8kPFnsY+O4c
Qu1B8lTUj8xIsrk/mAplZ+l5G/DOCvLvxRwAZbRG5kyaeDExScrWCzZ8bnJWsIWW
uYEEBrimvRI5NzvlSEgBIJn7XAkKrqQ8Nr1wKwcYO5JhImatdlNAx+t6tpY2PsS7
5cZ0D2QjXF9EojKZaVFnso/b5Y7uRtvmor/WcdKw06s3zkP/sorxW6KQ6Jj/oqBL
vATUz6T0HicvhOG13wmsjnTeIV4b4+aZNeICBK8djRCBKv4Br78ClwRpUrfzzZLh
h1cELdXeV5b8a37zMLJ8Ax+8AYyAjk5aNutIdGxw1K+iTw8OIlgURSMUwTVcapT5
d8zcH8ILKMp8/jYKCB9jFhMWEzHZTILrsipo702L27CqFn9bNnB5HBjXngPe7zmw
QCuIepzYdYcGqQte+TWrOrpAE9v1qKHXisOGpg48hBOjoAUh7nGxSiR1diyvwxgS
Cr7Tvvm0txH8iIjeAzL/3R8RgtsB+LOIahmXnEYwr0rVcwp16mrRwR7HmNb57btw
zIh3Igowdx+zXU7a5cnLStKLcylxcfvs+wIqXzUKRmJgJDa2cTrnoa3YCkeybw9Y
VW5nVcGbIzYevd/Tzq7RJLHgXBPjBsSC4uEIAue9drl2sK8LidYTE5AB9uO2gHSY
Q064LB+V0j1jgPahY7zJRWZ8DRfcoI99aAuVgYbny0LKJjhQ3aMRJSgGfEnXVd2i
MO6AvfwHkkgz+11uKamL7907ya7wqOdwBX4Ini5TfSCXTjwgWMi1/YsHZf73iAMg
XzS7DP2/U7zp6Hx7rZUAAZ3urVV7rOGcPJAPqMtL06pyLBOYVD45K6qzs2YJto9V
xBBxdWW3bTjFaCvvAvPJIig2e88WYU0anJu1xu0GkB1XQwZVaDf5HBdP7dMDEfGg
NNl+KYo9h71K8cSmkGr/30Tgc1RYbSam9SL0//Z34e69hfzo8FX2cr9Rto91ebpg
Ljb00wZtItttaSKoTA8N6Qvy3vk2z/b3HlsV8xg0B2zlQFATQFY+KU74ahagcNT7
6qOs7S8YcjDsDrs2+msXT38Qt8qvsKyOkyxKGjgsxpNcxnPNH6MeCQfZxuQMmGYo
li28WX4vLUjoKWkFSAAgUn4FsXhwowd+pGDOQda64Gkiz6yWunLtJdObvOVMiJZ2
mk1oU5BAmM8oNlEuRp2mzYeAKZJtFOAMsYf+wUB6s5qamY44LpVPqQvjOJRAtYHu
nPze+ETetcfsVV72FivuU6WiTvoYwcHUuzzYg5BcMH2dLNnfh9JkzWKTfTHX4HNj
2u4BWeDlwDSgxHC4f7OFs8zseD17+ftGpCT7J8qigFiCMfro0XB4Ft+kOmJ/df10
n6jOu5XzcL9sm7U2yXxxSHu6EoYJYjqhKg+tFI5sVaRwVOQ03Z4WAHcd5uQqASE8
SDNgbQHtvjqRIzF58XlqNA7xV/CvFjAZjbUgYLANq0hXnOS4Oj8b1qqPTMMzpJaM
PI3Iatl6ZTyI4yArd4xHt6rvkZ34HfSByoHza/COQNm+fgVvpsOxvfTTeMdKICb1
IURsH39PeoD9SBCTR/vzveknIJeYAsjKyWNMDfVuvcQpGEhCfKAFkdKf6aU+8Du/
ad4UL6JcVFi8DpeUUxa+4xxmTywngQAv2vFnJM8nN7oORHjZUWjH6SI2A7CDSYh5
dkTMjX9UrDiqoJJ3WmmjMAvwXqApfBGRHXlPTvmWs9T4LDZQHzqhEVCgTug/o7eI
vQ++EqbnSyN0yeA3dKNWpbuDtGv4E5y7D0XdAP/pnm3QDV2o960u3+0jp1x0pUNT
N7dk3MnVj4i3wEJExgvLHKdN92CvzkSF9lNUzTbnfaTdukino/Dql1IeRGhQxB1P
vGyslq+qoY6w9dbG7Oc9v47aWfjAIhpUhmxf/j44hqCw5RXXfyVrVKonjU5MAAL4
+tMMbKpIvw0xdPFeRqwaqDzgtqRPL/kztAxZMx1Jbn0SoB0tDx2LfrQLsnKnqMG5
YV1IqESDDsrdJkbF8JntmZSPF6BZxPlFn4rCQxcYAtkmu+B1KKsm+EIpOx2IYo1o
GqSP4D95thD5QAluDn3oc82rnKUJWrcHMCGWwbUARmH3a2aapx8eFZGpxQNxmsKY
UME1dcr7EubU2pWB7+w42cd8uuEbZYZzMIMOsh1HtYO4V+JrVbuuSMYLrNfA3O6u
/c5m+yEpEQfP82CWx32PcVFBM6IruxTQ2lSWjQnFRWr1RThYnKyKU6A3C/3k7QO4
zPP3sW6EjWxL5FGKVWLJKeYbhSdeYJBOVSSFQxpd0qTBJ7tnD4/G1AkqQdbcuooa
7CiLbPfEN+NaQtp/jlQdraGDyfZ0KSWyBNbdHiBc0hAtKHdFkIAWkb8IJeepocp3
VwMvGUw3SOVn4ESepuCrJpoNfTQt9vYk213aEhz+msISgY1QgpJmuQoNTAso2C2r
NgGnCSFR7I0GrslgsSYyO4n7Tx6g2wxXA+0PkHdzVRCOTYx0OMyrd3YFR6muf8NL
Dptz+B+n8aJ372t9oTwzzBHsz3AB1N2lYAys2EMiuGtT39bikUrAIbAe49Z4Xo5I
wBhkVAiBj2y+SV3hqeOF0yYdp3B7eQ0ApoEYZDBr0FNie98o5wcewu3Ak4EX1OPf
zwmpJ1oYvtVi6PBTWaR22rbUb+Ua+RuVBQiek+K4xKGQvIQXZQe8j0s/6wuYXy+L
eWqi5nhmb+zZL+zEAmOUjX/kcP0g6uzOU/HgJHHF92vYxk0/OkATSWkbfn0R/222
0v1Up6xxRZDIrZYBfO9yPGZyzBRUUb7uKCxCQ2NCZHHvpZDE7+HM8PiHTGdebaX4
NuhKiESwkk4jc8qHyRVQI+tF11rwVM2e7XuF1RVlH20BgGAAZswSCW27OfGfw7EF
tearqtI5e6ub5XJb8BDA4lny+WNEL7GD+ag0vQ5KMQyA4ZaRAXpbGZZ0GxQnjiiH
yhVxA6eDzBuCbwhl/P9iQzzJsmZv2XzSfR2obRTTfjnDiXiVLCv4y73uU3FNgtYt
4f9vvPBFpw1XMgIlGq5SumZC7prVvpZDO30VGknonGJkWQoEBK68q0FObVQ2kaR5
RWY5XCTkhMvXtaUdg+1Hy2ZJJd8JVQHjzmaV7SxQVsGCrNZH0DRZv/WGD8i/d3wj
kM8DJaxBODBr/oem1O5zDJOV9DCiwddslR/RGNI+SDUelaoxMdC9Cd8S8J68sbH2
gq5JDBuXnutzFbZE9o0yir90FjOnmzo8NhSStVVXwqAVOt/LOpg7d7Uux8QqiXW7
AXbt9jH46TIb/J3zlMEqJHWs8CLHIsCxuKp9hLUZR38UJg+67rBGFHsE6FEaJKaT
RYe07aHBe9ibK1bzyXqokQ+5sPcFUZUlF+YZOZzqvDReEbBBA3BlADqDeL6m+GqP
tUmkifqNj+pWFGye1dAmEUPhKMv/aBp4wCurpVCWNTH68ICLAOM8PIESejX+mAlr
fqcbrzXraPrzhuyD5UwXFexP2N9w1d5LelTdcAszrQ5S7aG/vte5H+g+y66+UHws
s1pZfCP7UtxUD1d6aJEA3nTVDDmp7+kjgRQHFh3Nx3HEEV5HlZBcIEaeqBSrfJwP
r3qlKAwXCrHdkwD3NjQy+l1G1grkE1Z+TEOUKT1AfAsruXWsWq1UCtTj4pKktf06
fcXxJdVLKgjd6L7MD+0dgKXOfW87WfjJLfm1AzG+r0uRbLHBCRle7IH6sBkRWzy8
/Rvr5jGtBrRekcrmSwd5waPrxcRjHX8pzQE6nh1YyFl8+Y18C5+dCQum/+vecGTF
lZ+Lgqrq/bTI6j3y+KLqpJsvU3AoIz05eV2F/idSVEDp56QrF3g5f9E7tj62vG3A
RDRvDGFp7Ykgzmdg/kotv4wMuiduM420mzBidQrmEEAosVCg1MhCBg4i9H3PpHX/
gWV48O9+c8pMxU9RKPSXwHBLF6emNBiJSoaqTjhXS9btnP44YGV3egx0CGSPnNeG
n6iyuQEfc64xsJzB1zdki2WW/voYCRDMbJkvU2WmI924k3OcQaQuzydm6nkFzk7s
k/f2p5P2prtDQlXsw6HIVthqj9qS4rv6ee0v6nHvQbPkleg2bSoLPxpV47K8/cMH
JTG7LVkptIBuAyILkj2/cowIddRdgbh2zK60+S7Vp83OQfXD9KtOIfTwdcXWwbQV
oggY8/Eu+N57T5itRa80ZFSI1uKXO3NX9YV+F05bCsa7JaBSvwuGi/cm0WVVi2yu
lXkoHOJwMJeakjSA9ly/gsrOKqPDzsiVZgGBshmOhTFZeOh9175o3zfVQyIywQHU
`protect end_protected