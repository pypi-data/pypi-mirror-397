`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzbgB/hX6+mh+pUJ6AzqD2vAu4bDKO/IptpVxjMX6EuSt
fWW11I5e9ZVu1+jfMWGWtQgH1IK4uVp6aCa5RJV4eeZcG1UoaQUimI9vLyX/2qWO
ki9RH3lxTXF77rt24TcuOmszJLIwLS6fjDM7iSHRM82GHFp6qiaXhB52WLEjXKwc
9TAU6MOxqx5CLjQu0rVxkLhguO44uKWW9NnxhunIdLpzrcOKkxInH71adAWauRfZ
1//lQ6Y2eaT388HYcJnzU7tjrbF+yrON5dMOQ761RFaauD/JCiggIm1IQ6XQpKI9
LMc8/DckI2dej28/UL0kNxyyabYSpDKrDxOsBrimsuas0+ZNPT5HO69t0vL1xkaA
UViJkuv9WrMYh7wtt29ArySN4j9kWVBEzZaak2ihfuyLNONjLbtJKA9iJrpFeoR1
n47mbYPf5/V8PdTADp9WgEwiijS/NVGn9AWaSlUWnu3tgGyTFyRNiTi3Rh0OUlAa
DprDvoYeVRxfQcjXLHsYjHHJK59sp+rut+OViiNcYxKYT70RXVqqJt1hL9Fg1fKk
/YvKi0siVIjykxn0Q0MyQC5XV3V9blG92hqy5XqtWa6H1mtK3cXAHN6nEiaq41Q7
CUB5FEGlH3HinKF/5ntfxmFMGXH9VZnj3idstJ/y6BJxC1OZTS4654+lyvfjjdpQ
fjcJ9pbMZSdyueGZJlavJwz94B0jU5zK3WwnwDFEQVqzmTshqraUfy4IE9I26/na
wqKmTf86RwYayk5J4D9LyCfhWy5/6xUmxW3IX5nL6oVB1aIUzKdIStJgQTyG2G5c
WELy1nTb+QOWKFHw/wUwGRavYN/fB5dXKtnvWmdf+uIDufq8CMm+iU6+LKJ0Orvc
qs6fNibVK0x7HsDcVMkV9Tg32IGXLWLjtEl3aAZhVHDl1YUSP8cy5obJmekSlvaz
/OobRa52UAi8xz9AdcCScpwV/Ga07QdWLar4Kl7yBJYsbyXlVSDjcNmWUiciUnKK
0XYKBNQBeGiCCz6pHs9UoDIuECvjYV96ExN2QmZv9aLBrfQH28xtWEfwa3g2ArvK
akaZMiGg5CEOuM5nMGxiryKpdBx98ek4naQ6HxgyrKLn6VxgDQZyLkbuRwrMXTFc
ZTL9VsaVd/KDs+Uo3nw/1hBpNKWocL3O3dsGS1bGsNq92Lo3HMOtVbspAW72+ALX
g/ZCUczXwrxKDAl72cOhEwqbuBhgBjQqBK7wJK+7LHgBJkXuDOQJ5wmaP6WCzWjF
J6fLXrOzr1QwOfElhLL8+VpLMaB3OWYFPYxUkZlcahhyDqy2MeZJIgn//cabLRVe
YHmmahlL8lPWycrZkKlh64ITS1xtw/UnH05XKCy/33NTAnRIHMOiF5r6sIR9kv8K
EH1BR4LMbb2hByHFcvY+g2k/4LWYNpqFTQgnL1U+69r+tLxaMFs4WS4R6CO10Bj3
yHUjCvCZMx2DzE/7YAhYzF+kOJg1rXSdZoG8WP3DBdGpgve+usz40NOTpavpL/y2
wPe1CLrRKAZfb5ZoE4DuBVyOD/fSixFtK4sYIVbSWaSyV/5vCLVjG/Txkcnejczy
O4Tu05qkgWR/hp18YaqEpZcPxgcqOxX1jmKtsDpwXgL+pa5h6RC6P+CVc+d1r/rb
JiorrJvaWOxj2UBINpSvyu9CdnkE4gv98pLt12W/vtC7TNUZdfEdFIEsUvl9KQeJ
6CCyJ1tYJ+PAfcqxn8KQFh4vpkbuSWyhbFQur8kjidaoJdvYUw61CeMcT5UWuY3U
JlBwFNY3+9ufJsqN22jDXCdyQ2cyjYut/ZM8P6sGUfRxmBZE3lYDuyv0MzYN9D48
soMpAQ0DX1v3tVJu2ET1iiuB0hvolBueWovkja97S5/2Ek6lZ8qV2KMG78XmmYtZ
4tlsbOnCaR/M6Hf2ZqMYYMeNIpb5qNGsT9ETAHR2It5hs6fsDe43iRFKekn2Dll8
9licNq4QbB4NmsHb1JSlS85M2RnoJoroWyCZCVpk4bGk12/ECAeOerNntHxLsbnE
IupcQtaSPKjjkHXKDiZu60ZLRi4i1LLuuGmgVa5jhZvrChoHzruMEX7V5jz2uh6b
okCx50hCEt5JMac34WijRX5j0NVyZ5Wd/z2UHfXg08y9tWBdxFfOzzD5yTjOdZzY
XECwuH1nh8M2u2wcuRKu7UHRkauBZfToWcdSB3O4gOahRVwftkI9YOBqom1cjPCh
Z0tYv/0xxQXs7JKxbHj/nJeJxxuZviJIkCbknYxeBBySX81+VZKcZGlTI2oP21xz
2rLkf4qyQ662+73M8eV3jWSfKe0nO4UPLprnuyXmboKhEj+S8EGqu3yyNVHH6BWl
RtN+BxlK5Aej1vBD5exvi+Id8/Vs8anupnV65wcwSS48inTBxfX5P0m+bwgJ9jrX
r5X0oCBfyRgL3tCn/x4+RGY/6Lw8ybf1T//Co92kB3wzhf+AIfg5KOBipRrUkIQ0
HY1fLD73O0xvM0N+ZPWRDXFzWXi4KPHQqDhOQvSkLF//mMCpwHWdmv3t8HdYVihY
8UrrF/fPDMF2e4E/Sj8rgxEB7SjBrPhrGrjdQBrDxBhVvRgDP1DGibiaJ0uMqnyT
5k+H9fl/NHFmGnqG7+Zfu/SpOpbHRdVXXFJ8AuYsw6DSJm1gnNrsbl7RxmznZl9L
+mRy3aPg5sfAWH89jIDL61m0jSd6HMxoyuigs1p4b5PPOGup/qNwH6ecSOGf8gi5
mOLHJ9M3Gc+IBvijoZDeYywey1hoy2j+lkVNua8Kr5ebG+BRSaotroQ882aOlgH9
dQOF//0yLPU4On4SLwMel2ZHohB6iY8zYywUG+Wnv4q+5zD7pidRIHcmYo7HnWy0
hNLRuDR9Rrf8P7HiREKwewFtTSgGDlor3L2pnkQVfbg9MwMxznDKiYOwlPLIKn6N
RcYe+iGMlii3UajoCa5RYjHdgh7s6oiGcN+y5jujeoVILMO2SZDSjmH4Mizo1IhV
BBEdsUHf0fv+kNRlAHC62KbYVooGa2eTeJxBHPEh8z2/fDZgxC7KTk5qoOWmZfDG
h0sSIF1M/2nN8HoKOFszF+w1G47VtvTALcLFPWzWZnCJ5O2LGdS/TmXr56gLlxdj
KCHu+OfCSIu+Kzk2Cr+4NuH2HJDC9El6uSOzpeD84TTvamygWnt5WISU37HdfmZ9
C1npAGCWNroA+YuvrYwgKXIZ4yt9J4YiRAnzOZEj3BBEtrVRx6PfiwPzj/s8Dn9L
WPvRQdtdwCshl20XPaFz5ddIYh0AZlS7NcnOklunyc+ZiiuN5tOKexPY8/G5NmTQ
z7H6bbAZoYbKpwbrJF8IPPmWVcCDUu7UlCcF5Oc8k86qnuiA9gEbEsBMRZh9irbj
eyJIy5F2ABsTI6ebsKp2VktLUiZgQrO9V3Mt0ai5LRKUv5ssJggflWggFiwrXbhG
p0Pxuv9asPkPbdLI3ox2cZOkjtV8EUKL0Uh+Xk49SKaNMunimts0LSJf02uT0yGI
8evGn7alz/hYuMGS+ofxr9o/Vvaodps9B4ABZaFANegp5Z0rqwTKqDAy0X7MxEW7
AkaAGNzHRWs0B7WdJT/9pyp6JduTnlxL5fNaJub7tb/xZV+Y7zR+g/CnvXz+F8JL
xRLMHDhmIfGdbeYBuDtwsB5jb2Zvp54dChdEZWJ0IlbYWQFdZolJGUpbx7CbPAqI
IBxYYRWMph+S8HRWb6r9KbRyVIkbG+QXGelA+PciTtzbPFj5kpk3k+VrqKF6ExOq
4IKFQGCH/SF9JZ2YoeIYqNcfVlX2aJxtMqxR6h5wYqSsEa6FctW9cHokK7GRPmwE
Q1wWVYCGtn1hZTya8hr50D0XoP+hrc6LY3mxkZkRcUUnKzAOs/QpCY3v7s7fwQYa
OfpukuRv9l30Tsrwo3CJs8rBoh2qjJ9FT61t6iwVRqA/dupCJ2LXlG490KKRO5aY
h6M7LpOM1klTz0rYIuPwlPXYZfgjJQYxuje6t1pJPzYqkJTVuTR4kSgcYzMGZjbS
iAsyEMWI8qgj9KI5eGANDXa33IGXc6TCK5bbexZJn5JplUMR5nIIrsPxGoRl3ofl
gaVwZUsJ7Uchs8o9upulRdiu8ZHgUvRTBZVimF48bxzS0bnGvsIdG1PBeUMJKXDB
LJwBQbw1OXedvroFTDL0PvHn9qzCzly9MPURJFsxM/0KmjCfDezEY+FEgg6bLvsD
Nf7WnOTnkTek7YiPkh9G558aDocBBnhbc0oWiNSX0K2yiH9/IcmHlxG8nSECpDwH
4nEW7kBjFnMi+PDT1SgcUglNmT+N8kyaFu1F07EaY8oiftgilMH2lEjBLsF5GEGl
QxTCspPNA2okRqLYf4yEgYkirGU+q+4JOP21NjcAFa1KEkeu06Rcze0dy4zKUMu0
CftKIPE/NqR52TJb6Xn0ZYOHxi856ebGFmgy1+vx0gehRF21D3SxIhkr6k+d5e7Q
LnE3NbBboihiZAKDeSYdULjlOyvUr5GaXiiXqabOeZzMGJpWOMaBJiy1PRmXp0HU
TVi4Z4kP9rmNgULtV1VO50jC0D9ujoWMR20/ajfWOjPGdrkk5SJMImZV6iJwHyJq
jJuqwlUBm4GZTUlf5WlJ6TQPaCO8HFKqkZtFlx7qYvRZJ3vKYTJWe3BV6lHEYfF1
C4bLL5bxRPY/gnuwnJ3WDnybuBijzVsFFMbEr3PGyl0C7CRnkMffaStprNaNZCUd
+im2aX0YiLKuTROoELECv8lXyJ/Mubsq/rBp8d+buSA/dNGsa/MPa5P7zzPm5PO2
zZxOcrXbm/DATZWEEmN9eycIdZ3EAfy3A9nRbCIP2E1g8PJS32FTfgQmwzYPGCjY
89tJBHqpJqOptFLUDpxeKwG0KcCEboxF12E1TKtvG3k0wixiS8qLz7J/pgJPMJOk
sJa/oDbZtyJ2ngJix84iePokTun0lCKlMzlFXaQRtv2jS2HpZ1BNnZZUZLdFs6IX
2Oy3WlfxS73x5qN6LYtGN4vkRvafsxijGcmyLNmvkUZfqUoG5loAozH9gfpKAW5a
Yap83HQDXXJwQtWaG0cb3cWRYTPLttuP6ytj0E6F5ubiCGUfzOYaJKxnwsbZa2Oi
guMukjnk/RgG/sEZXNlfH1T65JOfk9ocHy3TxAg0ZHLbXDwgGXWf9opVIEZbXPcS
e+h0TK58KADxqQeFFupu7cfKVhOTDG+j+oUolDv6mofOLHxYnbFnPAbKREQGqh3j
X4MWMKhkHs9EpkNqoxSttt1+qrwWpmgCPQHClgyBVCjs/s831939kzboV23inSi6
z7ovc241Pr6lhUqvH0/AwxePcTRakDA9RE8zwsEWtey33u6siBKjvnGtZH9kXyru
6fXeJXTr5N8p/relxg9EaY4sfr1RWpkRudEah6mmnD3niMD1UdHcQ062hcEC3cjL
UMggkP6mdfgkef1EhnXHO8AyOiZneJqw0mCPbi72FPtyMCu9XasrKA+zIXI3rj5r
UrXEPegK918KacJJz+/DSV0FeNH5SvMwdqZyBWfFRlCb42onQcUOitqv//TuMWPC
wmZhr6Y1J/ebHgtBK2MgfDum0qiAL5DO1x2VcqH+NjBf0onPS3TEtGKZ37nVsa8s
7rf1tK4ezE45xUikN41FhbWCYlAqR3j07bmbzGce+SzmpRfGrkPkacel2hzYGVsj
x+ICLkosCrz40I7HQhVmUNf0EHMzJqc+JfZ0+GYe6vbvq+DALLeE1aVFJFlPW/6G
YzHG6c4qr/ju3i+Zfg5Jf01wVrQ6On+vzioM/AJjf4s1hofV9pHgd2ZBnQoLTcYk
n3vTogXgeLfalivsTaw9tpXyhkig7j322Sv+KkTwWt9jnk3hJ0CyXZ1wfZAm4k/C
rq4ynwcOHNiPA+gWADpKNGfSJt1mKsObTm729rW1TsiqlcorpotjXSii7HeCZlSc
nqdjLOeow6mrDnvtcedSsqB7lXcqMZ7wZuXJIztc+iZsxDMbQnLG2zOX6o2fIHai
kwzixeE/fZk2FYZhPqDh45YSdOrj7lhKGf+rGGwcCQ8TfFCuwVHXHNF6gFn5qUGU
aYOVo7RO1wr1aU1hrd8C4FfQrVoH9v6xe1K/I0tRcmKuARiJ3G5NHGOtEUDQki09
Yld7RRSmRD0vdmp0qJyAfRxqPs6vkTt/OI7RZ+jfsK+Ot1UM79yNMn5KiPh4tYnC
yuUpnnSM0VhyFgSxtYNsYB3kAOA7gtpEF8azmyhopWurvO6dfzV6dhy2U9fxKq1A
OMvYWIBFDG8Sbj4hg1wwWx0Oxhr4rGmqU5YjRSmffk6JUVa1PhU/ng90kcpb4QLH
7zOYag17qWl1+Q/fNi5OCfc7JZ0dOezUgt3jVvUSmk2KaGgsuw3fKdMdpQe9Q2E8
XxRU4io0S+82CRJQEcTrGjXbIw+EK8MUKbB49/3G8cnzlKJ/75Vd7WuY+ICoq2KY
1UBfdXk8WYuMVZVdXtH6atHHpH943lWsbRBscE3Hv8ois2hi18RvGaFbyL5PSyds
NIIBumjsm6tnZNo/ytPolLJVA5lGbQFzb+upAZ2ZGuJHTVOg66UDaREtSUikLpmy
iqPPH0gR0sgAzDkJ5EJfjExS2p0IjweC5OLDh0Mg+WSfzR3hPxssffTWJ5kwAius
kudt6NR4m/NCUNHcf+Ms+u7Et0qRuD41WOJkMReSGmduycv92giuhKoQPGHesRWv
vi9mE9LCgvNKiUpaeUt/jufRhqCFClO0mp93iigQTbAUfNKCBG+8MunDPRU8hUA8
M+RDPMGj3Lias6h1Hp9XULWUlv1tquUbcSpTsv271zNJJ7ZlIhXIqhgYmBxLYd+7
N+CMnX+g2wsUj8z1EXPgNknhDebAxUmWp60wniAxxdaq9MFT/WrqDgc4Up5Dkw/t
3g0Q0dcK5KT1eqxSAcpqN4+RVIIHWU97lSSi2qDu239GGP9rnWtVQe2+54p4HNnN
aCh13KvMwEyPyNNRq/zi9uykeUANIsxiIqLhx7XUElPmocRY2Q6WHeoyOVpb5TfD
tDo9qNNNuBJI8tKYMlUt+a3WGq9StxNK0OHYtyZYuH12BSnrRGjyiDD+bxlKy4Z6
mCZl2EfdU30D14ZR++HmrSjc+jkNobMmqQpa9tbtP4xth1+ldJlMCYus8+QikX8I
Hecqt2JsTlkT/13/qZAkpCxxU/aK9HnG2qWmqzaWZ7Jysp1z4Rm1Jjbr/dtvorgn
EdGTQ5INuoXbNH2yTxkPySVhsvJoqqJno3F3QPLGqyuQ/tK8VFlAd1ClP+4+a/vd
Jdu37t4QxRshTn2UfRKVgZz9V7LJ87xePczwNYW586mGqBU7vB2zcS81EvLNe9A3
7St9s7cYBarDCUXgwqC4V/M+tcY1IpRIbepKT1eKqcbgNgq+deYbNZ/rio9r2aTM
teD09YAkOTCFpmM0Cnz4qphlVeR/APMhD3ESZrN1uLtUpfDHXCeWNyhHJY5CeEnj
cYrqkHxWLedwqtvzE0a1M/8rnepvozAHkPAZ46k9FnaYIFkDFhsUKp+UZqxpslBh
iTRhaOc3ZTPKeShqYljZFf+sbxUCj+KKHTv2d7vBC9i8Rxdsr328SG2Z1rlSAZzg
B1UJh3UP2vojGecchz0eNIpfIhwQZHoEn5gRinnTtgLdiiT4M0jR1QUwAAYm/q6F
68+Hf1iXUrFZDx17CQMDJRRW3CIwjgd08BdTSjnorQ69LWhzQd8ryLpXSl9geetH
KXKlnljz1fBdega4UEiVeyi29FelfqUUpCb00dmEttq853Vp/QiXTilDRRpCGF8a
lRtWxNCRkTSma99twlDQVwm/yPNxEgg54zVmEd91rRJlay/EYrSqz0Dpbt3cqeVy
vmDWw9PNClGbdlKqde068Jfj/k9Fc8t0/117QzjMJnMEAgFXITb6ncoz5olXlTda
tEzjVM/MYQnUoovdxpT6UuiiYuDjxOvcHS7PD4RTIOZA9ytj2HqJ+FKuDUKqew+l
14LlJvMOt50skwCKR6kXxt2TlbP+7iBraMqvrVtuFk30dbHTS/WB+XE26+dSSV86
sdGeni8bxtcZSzNgUMqQ+VrIgN0hlT/rl74tWpP55aOKVKVDoiWvFp0CNUpgMi43
cItxiMyePUeJiDWKVi+27DBlycmdHhU0P+8wi3kryCFpjSshViBbVZ51jkV57lpD
AiecZeEzlcKBN2Z9rLP5m19/WEZuaSJvliZcIJWOHj/caf4w1umNx6WMkX2ChtC8
CogqF18GWJTQP3VLX2DRfqXdJ7bam4K0r/SjHM/K/oDRZYy0p2qyhvjajG09ADUV
GeC7HhMuX63GBO51ilOF+v6us5/8yNqwLM6nVqLUkXVmk/ZERAESHrnYWsdZAet3
l4BFk5xRrcqu0sH3y5bj8EB1WQYtTCIcZY607M0c6PpUi9qPGsHsTU85606EDADr
8YJF7cQJoJ7oehXVrvl6EDAXqCogY9/vj7u1cSUiBAc4YwOjUX5K2j/b8/W6HPY6
FwLvS6UdxKsCyzHNuc+dGW6LWPJxUgT4iebU4dwhW5Ieem/vYAmKtGNVLKGhre10
asWh6jNkOAszaeOf8hTypiuABmwSAawJagv2WujAo1000NvSes47FDM90w4VWltx
nOv77W/P4sQZyw21iAV5tM5p49TTfUrlL8N17ef2eHFwipYK6if0cFb21Sijb7t4
Kgi+H9P6HOKsqCFIP08OXAh+/R+i+hoDxIPRpTAOVxWhHYzAnSDsJlf6aRurXjTr
0U+xnhaXQOX6Pe0CIprsVy1IfaBgSCuf7v/d2wlT+4Y91O5J7iBiSXooGE19zmQ2
wgX/ighZJZuHGNxzOrkXxshPnLyiAb2Gv6tybheriGGOEvjpGy/No+/1eHha1cHm
BvtBLVDhKi9JLtPHRJrLJFpQwW92tyVUXC3IdkjvZ/wY/mDFoqU/bkKE/Sn6TJiF
AjzUNB+TyIa9aFNnGQ7ZYJoAdNWxrYAgZRLNNWzX/CMZldyjQMm+HvaIdRP6USuJ
2CXatPxo+A1naIgWN5sZLIG26JFTW9I+LeTzow8od32fFbdTMEJfwzd+rUE1BKzp
zva/KlFecUdACsS2Uk1Pnp9ZH6PsORf63GHiVZ37VfOPda3k2WQt1Fx/88I+f+0k
JmJG6dMFt69wyin+mnXgZGbKoaNi6Phk8OiiY/ljM9BSfVwVc2s6HNlHcE/1i0H3
wE/w10ykOfqTmCk6XMvCTH3RUoAGxUlci1HY0AgBOE6LwOMRoRHVJ5QBf1547tCK
jc3XO0hDpv7qeb11rx559ASz86m/exBPqpPTujCncuKV+PpnWPmOlgSmCXwFDQZK
xe3u//nLhG6cq0rL7Y75HtRQS4LYwNk88zkNiUGh7L0EEIuG2BN7bVOR2bVUE8Fb
y7ZE7KeL9OWzYsn4QTbZbU6DVAM/juXDH7801mQ7OLzjat81Ii9NpmMD4urQn77Z
eEFqwe/XtrNaqTfjM2Q3WDWaSG/O4QrIdbksFrzxRZjsCXLEx/vh5cTkgdnYx36O
80N/k37KnqnCL2W15O43HiGYD2wEoT8UADLpBP6HuchxdX3/1KurOOsgIZfmj9Nu
mNndHeqaTL6mMDSXtSKyQS4dVajRClv5Qp/ZDlvC3V5ZiIX10ojFsrfYPc1Dm0/2
VRjraGBTqKrNBugFIb4ohPv8RoR8eg0ECQZ87U0cTNrruhTge1GAHQ6dR8tWirKV
OVXLmddQefeY3NTrmsWswMzo1/D3GsB9S1OjHjtUfiepSm2M8/TLtZH99JnN9Q7f
IGqXBcMMnQMCnszmLdAzHUsXomF5AcnZjS2vD65qBFy2Ftwhwq0+IXVozL3vMp7I
ug0Gv1hHFZnG20VgTpJ5C+97bz2RB9h/CU3SFGFODqXrZOAxesUzUElf9hcfBR0d
56QSx08h/+GpjM5iQ5FxgbtS0A//6jrlvfy/3VvriUCcwxw7XlGPFl/Cax1Uq1kE
cf/kaUd5ipITghVEPi1vAWNN3yJ2rex5TcS1yCYNwZThGQ9xI0ZPGx9heZcgX3YH
gA1N/dP6ri2UAr473wonLgKqZATdClaEy6ftXbjmuP9m3+lXia8LWGymlhn9Hz6d
FtuJzbq8j/dgmA8bYy7CiTpqKjwwgwCedzfYQksnrw76m6XQigZoHjojQh503eQv
d+qM7luxbt0IgACvU2IBCfPPGKcCEo0PHqQIXUfDm1J+4OGwzxd5D0xfR6eGhWQy
P6jK55MCiru83mAQkINEsuKhlkmqU6allDBp2/EssmIqsJRxSew6tbYOMApSG0Q+
S+b2bHGZUe7273pqki5HZGkSmSMay4YL3ha65/FtI3ccOFp3mbs3kOobzdIiyMTg
ZpYr1TALCbTX0R/RSSBnke8e57JucG10AfkXERRsPOKdfzYwrbgr+dY295w4/Mvg
MoyznyHOg23nt/qEHE3qjZ8YzLkgTe37xCbt8W76rCrXGbaAW79D4MFYSrLe+3P1
+hcdxus3ns01A8BfJJBiMfRYc3rA4ESciXadTKmEp5qhkss7UoSu6Ez7nTLo7ttR
OlqhImWSZTfEt3K9iSGrjN7Hy94+DiJV9dSiPIS68D/5rhlgB6krfaurNgPyxG+R
KDsdhAAIkXqE7B7xrnNP6Pc8wQWIUycTiLEanKenVThFKq/rmiIlCLWsszPVck/P
JCrkJpQ0aJxF1J3Ct4BvHQoYBR9WsDyLF2U0QF1NsUQCpFLBTTpyfrmMqzCBG1xo
QAQNQeHALXlrL/npVV29gjVWIZD7KlFNme/mZlDdsHkZAvtJ/GYxbjbL1E/1ms+i
uZz834SjY1AJYLqIj7jNoHNN7J6ZcxUnMnSG36IWRsW4smL6bMDXMCFu+0+SJwDV
IfOD8p7uQcivwvwPNuztn7YmHotI2g0v1aOgrXNDgRIZD2slzgvctzvfhWTcJgpy
xM5R3Dgzvl/ScElSzMNysUEkWHz2+bfYIjiAcI/+yJVmys2/T4gq3QBZslfV5iau
UuBGfQUFxAiYw17mk7Q3S9Dgt66SPWOeY0atWy2RI35LVWl1ujuYFN4W4cLfgHZo
rfz2waCFANCbkxxQRb6BoeaOdzbyzdjjBh8DMtZ6WM97YWYAgqO/FY0AHXpWCdyu
qoPSMHsjRwqjYv5ElufS/2ggMUJ/g9ggzd8MZS1pKqOnt+Ibh/YLwfSkj7sRLfg/
3+k3rP55Fh2xSm7wgDWSNBLkA93sZGn/JNz+EYF56AceiMOJjjhMFMeRX1GnZcrL
SnxJyu6eJxa9d65k3y5g1FcXqzDEu4UuOprRl8EXso41ixvJ3n1qcgMsEPqi2MbS
v0yQE0NpNjK2vXAxNx03j9pMflLuprHH26S/NxjWlO768SdNr+fm9BwAnqB6sZyb
gLHzPCgjXnKKRq1z8Dob4tJQ3GBWOusa1LQBCIogNIYs9WaM3KyuTMPSQZxawY7V
sHJcSEHB/bVedjICLIcMHYqVPL0kaG4UFD8ii2AsENPW7hnvxnX49eYkKfNbMb9Z
9c7L3MpiwAb/s/G2Mwl3QqRC4PpwmXHQPi7Y54kNSA8nGhyOJFP2j66IPDE1Enik
X6wJuj6yv0dCogLwT8ez47x7suLaTCZMK3hLWu30ezddjQtiBtgxnJKa712mo6px
4nxnfE9poU4eRcIC2nI7Tn3mOCssqlvWgy5l+XlF12qpTkiE2pWduh5jVvOKa6ck
10ryZbJHI5jH2cS0VHCJ5qmmiFcnB3OSEc3ZsnktUl4KhTgFocDdoJjPfqkuAeNB
/VeZOEqVAKfjgbjbNboOaqubpRXC+ieF1iriEDPcW+JwsAnUfMcma82+ewsqhdoO
OladkNVS62iv72g+gAkdSVaKvH+Lh6iINA0mHc4Cl+eueLdiYYyWMS/3jL9AQqkH
egK9MT89kBE0npXPh+NmhIurQfzRBUd+VHOIdsKZ89fjVj0jb/4uqpPY6CpCpr2k
KlmY+/nK2g73ZrdQ7hCrrKtyOfDpL6ZMJaojyo7+kopVKx/YPC5bhKAqQ8cgolR5
3p0LXsdlM1SC0oBSOepPPrYNxe0yjYprQ14CntqQIfx5stlpuzmFyuFqdN7urHHe
8RuJ6eEQuIxcTwLR+qPQQIBWennEs8ICsbX13iQkVNwK+E1G3XOkzZzidtigSy78
Vz6PMHWowbidgcYeMW1wfBE8f2GihWQsmA8HZkMfbMMev0+klwzL2Xac/8Wvt3oH
YRLRaAAd5ud09XMXEj3L2sXelBZAPyJxOTfi+gzZ/8/BKd/dr/CR0w+DHuU5SB7W
y8Y93yhiMQXR/wNstKxpZIXAngT2LUeTGt6fU9ODYvXLgj6F5zC/U+1pgyCx/jX3
B0tAFqeUK3cRKNk7gPv86MhqcD0i8LRuueBFrLcOGElAEsW129HGoGHi3H8mlGiL
4EfiRfk6Dxtf1xL0227gT/o9U0faOtqkic6Slx54O+enK5XTSp73+vo6sKZy+iNH
s6R46QlIBHNYw7ScGSoUhVhg87JyLt8tAyHQeRMIVpkEyZ5z4SPIl/PT7XbenDYy
KQ2z9EwyLmh067gVh3umJh1K/vOP3h4aWneGGTgEP0Uh45ViiXSe2BZxuVVNiFMN
cB5kBNTTTp0hZVSpGQbhCcL+hY6ip9DMDDgFb+DG35v+kLx4bFWuSYvjOZ6inolv
CiDs6cHtWYpiOp26eCWr6HEiw+7LyVh5IhVWt6R54kLnItT4kJaWaLmzJvlu/Ojb
s9tqVRvPqViDZ5J5uVi6v4H5YdW1ZYvtEqypYCRpJzwPHwWIjOumwlUWMXeX7zQs
uc4SgfcE/1uP3g5mJ+pSa8fzKuv7wtkmmdh0gLBnE8vvt6PJLPBC8uhfC2Uewrj6
/ogXujJ/si5yctgVnGkrBNtv061WN5zicBa5w1NLCR0C0bMHP9jH0prNg9/1z6d5
C+QGB82WPWgIrqPltmxEKW1So9sd9H0lG9n2vdsr9T9UOnrF5EN1DmfCaHDMRxVO
5SOmJGpJPZ6ngHNhHUCCKz025LgZ3RRfBwTaqBjmdV18TbPMoHeXb+zbQqmEuD1O
zXXu0I6YCFUQPH5a/tocriOaRl83WrNgvDLm3BGLqypuTkI03sSTFah3riqq/503
Up7siM2XaJVQDFkjqqgUteZ4grjJIb+CQN8LNF7umGReX52fOeqthXRTqgTmbE1d
+svE8sIbzyryq/7XDeUJcfpVMbehIo1QZWgwbywaaRnMQMj7b5gln0VOmcXy8TAR
s6ZAXvcrVf4LhLCVpO7532vTgZKyZw3XpJR+1+JGqD3s4O5NUfZxr9fgo7KSBMxb
p2b3XxrPISjUx8LrWf2g5ODPubiCu47M5WA9VO+1Dnfwp1yhmnIfn3X1uVK5ndUq
Xs8jEUbvI5nNBzM7Qc4k5GATkv1pnlIRaf5+5U70VeZCNi928MbLX+RJZuBwc2wr
IXlbctUEimIzV/LyB+ShhrpKQhcpVqOO/c6LlWhOU+e9LUBXpORLYX+38ZKxEr99
xmcS9+0QN79XqDQ2YSpTXV5dmiCOFmuMxlrUcPQO+2FHFP0xyQ0aV+KD2umuLo+L
qaUxpbf5cDDbcihymZJRxH6AzlUwRWUEYP9vjgTynxdIx+gg297ltOqASmd17+h2
xTLL+jM3CyBHv4ymFszgVxZOJ6n7YwPBmOTHc19oWMHFmgED5JI9Z14m9oz8zc0M
KGqU/aSKizU9VGUE/VVlVQYx9AlQQL1jS3HLlWs61yjVQvZ/EOxdOhIpyb4q3HOH
1zlv0EjpjNyXciks/KlqUejSrLPOxO0SYqD74V7S/itY0M0E7OkXyffBmTtqd7uq
YeqaJ6j/FdoJWCScZMSThuVCV9GYR7OazjjPfqjyEBBuEWhbnQfDx+01aESraTdu
teKL4yPoh3D/z1VoFaD7H53OsV7/g/SO1FCPd0ModTX9GHoZzWgsiTpoQqlv0MZt
pavuQXYi7BObiwgPzHtLsADJGdxD8Kk3+FEIifncTBqhFtIp2rgtm6PHdv+/8z9A
bOX3SYnV9Z6Dtlvd7c+r9gkxwg+KM7BQmgzPbdBDyzuQNJPhySTLTFezbxzOBhVm
8Jei3amrqx1JQ5fRf+6iGmPalLnlzJCw4rl33JH/BwqfePH7a07VXMSzYWgGb1OS
ozgc5RQLX0oBBMgEIu5EcoQURu3ngkJhe2ZsY6H7gV9dRlXaRvjVVBTzI7rW6YbI
xBgLVra3hJIIv9uKsSePxETePrsiB3sscw3YP2qpAcjHpm7vRB4eApnWHMD+/+of
VKEbvxEwEsTDTtXjRpxvKoz3T6Bs31BQeJKHnuI1Z/NHSy7Uw+dF38hDglhIBDuR
1SucHPFJE+lNCILCBy9bicJU/33rPCcJahxEATPm26z6N+DVw6Ps1qmerkUk9STS
7VuxxQyf32jsIL81/lIwKPJBWvLxNsb/xOkWssK8o11Fqh3anrpOF3t3vUttiVYj
JZcvMzD21kxmPR3a+SPu06M3Fj9IJHojyLCjkRmVV4gekL7q6n7y15peupOQaDwz
KMKHombjaH5ZUr9FhfS/bkP2G8J7j0kYnM5iZjYr8h404d8gkyswVApW2l6TXEWM
Nu5+g2/Zv4YsboatWbGakkAsIEJDlnoNgBab0jg6f7qoubmRa03vaKcEWWt/8K+y
16cB96/XEiPyoECZEghiAFDHmmqnLCMXU3J8RO8syYqCJJt+otVpV8+5T87w7pjI
4MWa0UfEs7KU4W6hw3469VUVINc4ZWaMosN3wMcBGEo73Xs6lAPpL5+5xB2yh4AB
Z0th+d4E7x8YqnEHZlqB0kGwTMg9BXQfdA7l/MiTOt1iAgdfpb/IC4NKtZ6f18My
gLoPj6ASn2y5dNkpfJ1h3SpA/W+jfN8CBVmK8ytdIzkX+o/uztuRyuN82mACizsF
D95GvaZdsmgMHEAvatCCHeflw8K4Y2tcFPa9kcqt0n1LVdhlLs5VdOp/x5zzuCyg
LL1baoceqybwTsOcRoC771pK+hy/NHwHnoiRL64To1tnLEQBXgNJ2tF/OlxsO93W
yWAjn3sWHQSxtw9qrxdm1+e26R1LWV29bQLZaYfcgrK4apGqRDnbjuWpW1SLkUbU
Nrj7nyNvfg1xox80JSoIGHNFHu3E2LY2bxkGd6saI4kb5r+7OXyUCGgbBEa3vZS9
b98Hoxp+up5610KOyu39qxDCYUyvDO/IOa7XJlK+jBLapwslB1bMBe8STIb7u7Ec
UZY56OQchs+30roVO4d+/AfhYAf9cs4QZptnI4oXl83LzsCFdK2hnV+8amLUUhEB
7NYxO8lYi0spHTak+1104yL2+FwkkReCVUZg4pr/m6IPiP58+qPymMANSDmH91gD
Ss4pAIhEAbCW36hgMAWEcMBylfYiwaRPcAe1g9jTqOeONyNKqy+RhwV59hv0npwt
wPeT9Dbub1Ukv5VzuzcOy8QtnlitQQcfav9ki1se4Gm3m3NNnohEFrdEbiZ29HMS
wshVO+GqRLCNjyhkP+/8WUw+5dHfx10vxuLGygn6w4tBxUB5Tijm+NM2QtCIhUM4
zuJfFrhmY0sDyLgmGbkx3akLjH8LAsEWUucelJOBO/A/DEOpj9J9KRn20ozHegGX
fe+T+kOej2ngxIXZIPhw0AB+LY2UXFJ2dHwQ0Rb0xaNseMVWu9OZdyvAlxx/i3D2
Qn422IvhYLx8/3SY4/q3ScuuAETNehihLxDRiojBrZOdqcQhLtpKYnIrYu6Wk4po
ztluRAQ33vuIRFMzm0ot7Aaip65SbT4n03vI2IhK9uBdxZdGZehr0gv30vW0BAVu
vt1ydu/XAhz+ne44/1MJHark2KEWKQCcRtYGdZ8BoiVYO6umMm1F3GyaCMWh66uy
Qubzl7HVoqu5+9njilx+8/rHwdmjtrE4qJDyj4ywGyKy64Gbf78jBe4LLoPcJ/n8
EphUe5cvSRMxwLr97weWPt0bbgCzI7nWVtMtoBFjDdl8dA6ncqF2RK0gBO7ggPuN
8uCBMBxuGckihK5qApfDYaXVKjSpareUTpiGGRsqtgwGGIaz97q6flMRH25C5pIq
EuoE6wWr6NTAUvAXkdqzTl2HERzx8YLWM4MEXOzDxqfDNB7iFbv2Cd66/kSg3qAY
i9S+E4P1B8gVgByD3MhkJH6lyJtHSDiGtEgNbHxYE5yjmng+PEeKXTOx3NSuTqCB
DnAPtkcYgHVSrG2hFxK/9/SWZk6xwve0WD7Av/PBZ8wvCb49V4kiIN5bfUmrLnlV
lBp/qHe+NHh+gUxF+ZXUIq+3rJMW1UrEAJsm7zVMfPImIS6tKyPuSfVeXvQP2Ero
ToVIEZg2RTU+/h3zp2bAYRAxwDKwU8CjuqYb/zRtNr4SJn/w+AVYxI4UHCSrMNTh
VhKA+K0PXIv8hWb8aGnePPLO0u2HXHvK1OKXywWgfR3gFNKnnPPzAeKa2vNg2XAB
8nG9S/26vBxf3lGbx7Lp41DqmSUV/pc2qWLIEIs2cgDeGqmVYUva7G9yNOoGMjPB
3Elk/tCpWARPWLL7Li+s3qIoyp6Z92jx/hbdUYWGkzKG11QPXCZN2OtB5VWRxfFO
1si6pE2Lovwd+cVhStgGITeg9RV+otpMkHrHh2frM18vh6e2OaKD0PlJ4pQNGqk8
S74wCmWv9462pzkuTcWTbZNaczab3Adj0xQGOnzVovQRw7eMKZc9mpUCObZ/Ch/C
pHqRoz2C0kD2oHiaVF/Dd++bXRgQ3HVWOLhVl9w2Ut29Lga2zodHW+7keZkE6Pe1
F7OMNHnRI9POciUMT0rBr91KxHhU1FUgr7zPWPoiU2buMjuf/xyFNCZn/VjJ++JH
pukVs9/mlb4I9CMQJ/D3eBry4ISHjrFfWbyXhM2PamridHhKN00PHcn+2sqVySlK
uDsvs3SItZVqgkwWTC+mtesKtk+lIM59mnkc53eaxXjRlwBXQ3M+MmU8Lc5YjRFZ
2IC0yWYjyy8C3UPxzqbCY8FO1hnPG98Sr6+RvSboqOPhaKB5Pu1rHggMEmUk8sNC
G7JgMy4FLkZvg17zKeb+NYOa4MZZs5sc6VK228luXdaKdToYxmCkmhNgp9tNeluh
lLnErPEyUtKlI02j5288XMLaUgyfHhroxU3QnZt4JiCS+uc3CZ12UK4TsxitJW4U
0UPHI0PdBtzInwzkA2TR06cirvHklBFlgmOJeP/EvybS/oRoiuvFZM98/AbPyrFy
qmdOHrWsn2wZLaxBH3BnvDbnPcuTlkaa0wHgji+XqHxe8Fq2ywJCscOJ6MyfvybS
sa3QPIrzcKs4/tTyLjNFcQeW+ltMucBzVLQk7MCzemWaAmbqInqvgA7M6SeHtt+b
GwLyVd25EW2TQyGPbl5d7hgUefKlOBbOqkUydf0yy6mOC7efsrIJFply6vijSW4+
361r1yQe5lesUwlPIWgIczA2SHGUvlh3O2nAqd19kDGaE7cgsY1yyouvoWkVAlfY
2hesT79q2lLI2U/JrXBJjthsSf82IEynDLRNF+pcsop8xMUCWRPSRAgemi8japyH
+FuKZMvCGmhb1rqZ9jduAt7gJ5cS0A/73b7yfs0rp2HQ5CwVeiF80YI1VDos/9Xn
hh1qx0ZRxJ4hR+AiJEB/wS5QtJj0/k7ZcxIhuIDTPk2LhCkE1TJbYn6G5wrJmJiu
jrcInOrLhNN6RKNtuzjTUQJEA8CX4cgKQ0vtwC0fwmsH943Sc/3pXv9rbM0j0QcZ
3wzq+VbJ5dOWdmFaU783OxJ5STHVgbCiN70ELWWercVcV74dNA0pF3Po12TnqC5e
qfilOEEUb8GTE1CbJgrrXGiS+43ImgmYYbGohQ9jrIQ+P1FgO9YK0l9gvyQLyshK
aT6W2eAOt/ckSz9Hsmnx9I41XmRjeBDmmkjht5eQ2kwpxXtZeh+Xnw7qzj8XWz41
HATVPO2sUFApsoIaEgbLjUu7zrGwWsLIVaUVjffdtp3bXDF4+jeHP+5UyG51iZWz
ptPoCHh4qVlj0dYPLnk8bKOdHFqCj/XvTZ9jGt7G/YW0g0BBUgig8lm3Eis8W61V
ltcqdjrBuZ41fJ6N6gjM3GbT70MrshROG1IBw6jJZtUQWvSN05W47tvX0E5vFA2x
P/sJyvrpH35sUf2wlNpimsAsY+ggMhsetcuYIWGAnEnfTl4l0ov5wOgbGZ/IIf0H
SIHBR6p9XBu2AawKGHSQwVywGC15KPPpS3kmYwVu5WV/VQ25lF2HJoSnSJsqM0AQ
UGFHg3lNaBGoTwv0Pyn3+0g/3mrm2n9P/u6bDK6q1xm4vTy47xisjGzItwkuZKSx
wKLz6BfLf++frkwQGIbexrpFNAdVLlStsoksrA+HkYKyAa2arnDP9q+rHvrACx2b
M5zpFHIrnsdvRh3g5DMspByCS0nBmu7P6mSG6W3px9Hyb6hacu6jlumqrzICHNqe
vk9Hw27Zbp2wc2JDrH6LV2/1sXcEIfl1Ok0vE0BYHPA38e7lI9+NbpTf614NOIaA
+wHosaNfqkc0NhkJVqnpT9/kl+4ipjeM+veFaMd/MqorCudQ0S4olQJnFNQ0wV1u
vBx1rAouNsw7aE9JQah/7stjxyOCCUKU/KZdr7Q5NvqtOFFpOFG4ne8xKOrKu8QZ
VI0PvY7heKnmfyU/TQzCZShRrdgPVj8YwUbt+1+dATgEgKgiVax+9fJzz4gNDBzo
l1+2Uc9ACnE1gWQwXu0o6Sty79hsJ6yoVhgZnlieSeBKXS7Nq8b4ZpegBhMxYEa9
/L39Lg5C5uMXlKPmfiv+bruqPCtsgKVWb1MiOtDguPukzvXyD/+ZQM6JTNBKpoQJ
An938jIEtwLfuNwjo87PP3+PcgSBhymLDweNjovMVvJSGXHv6AEGUiBe7H79QWHz
LbuRwBL2pWr+QiIEdwr42XWqKgIMLMkdxeFUmQtkGF9xgmugGsvV4hvq/Ez+nJhj
4rhccB4ZqeCOUZIlDU6vgSi3uuyX2zav2VdkT6f+gKzNH2ozkYseESR+MLbbe0tH
95eVCNkW7HIR++WR9wZP6GDBT9RXR3w2z17giF5/zDorroU0xMH8lR130rZZ0lry
eMuMkbP9Psh/J4ymlO9HCaXUo2qFbT0Ul8iDqoeTmUXXV/bZBYynXyvw8JM+lh//
OWyzNJnfSoAkfaLx6bHUnOoUsUqRg9EIfnNGabCNNsv/mgLL7uua/xmBNj4hiCaY
8th3DlpbkGeH7fZZ4bIaXo4G5wAbL8uFgdbcB+D8E5QcwPrmndQ/ERVdgQuOyvv5
4p37JaGay5vaPMM+MIOJ60bhBXO2Qh7hG2fwFH8+7IRntG4piA4znpI0fIC+xUwx
QbdfDNhczOPcvsBb4WHnbE4S+ir2xNJlcYphFGB4K4XYPFoTRqR+zG2WETbLjquL
JBeJote82pMaJr6pqb1ggoiCx8B8lU01n4FnoFtMHjTGz8CdZr46IBcW2yFtaSUR
wkMLu1kfWQZUaCoyrVF5ey0ZILV+HMm2J/uUA13DaQz0O4X6QS4lBKCLj6r9mMVR
yAA1qB1+DLteD/O9oC3h6nN+gKCPPwycCoZ78I5In8GsJxKznq67doC3zwx17Qf+
MQ2VdDDcOIigbVeLECblBktsFve8Jz9rJOEZJ7ltuEiUylq+m3lHfvfNgIHFXx7K
E30m2OnxKrKQe61xMKPQIBlq6MOr+jplkB3Q5rdviRv+roZGTwXN30xK9tWiZI5F
ZSLTNdR8s+Yjaa5vHHhvI5/C47Tofzb9XeAW1CKqPHB41B1+oXEi7aaijeHL1AXT
I7uBYpn4Iv110l0ysL/f9v6cSVdoVa5XuFPpF/V/v9tXoYmVK2s1txfYGASHEqcb
d9O5CeyNSPuOt47DlBI150IzsKw0QZbzup3bkn/i2d5WbveRkGHGfjTFQsYL61Cd
t8bSwhQ21tkMP6Bc4+fHuHD+fIkZyLcXOarPIU/I1SYo3wyu/+9BaSHwIYJyVpMi
ciZSkTLIkTx5oiTyr+tP3rIi/1zoOCPTNizdziM7bXpNjRtQgdgL+kwB0UPrbkVC
vtvThzQHt3CfxsaDO0chd7PCHjTKImCavem7QRaSMjUV1ymgE/WyZJgCAhFDQ6vs
qm6UU8Tyv+OHPQr4KNHR5WrJidnhBI5S75ly66QiheS0qckWqZN38ZbDoZ3NfMxy
zyT/pjCs+BCgs4hccRDl4b5z+EwwTX2FsnOxR4s9BJguPRdxXaRplB/rPaj/JS+b
FeqPVRvZGz/XfFdc5SOGADgX+vp+A8jGpH1ZWBybod4nfw640YXCe3HyY2yLG+B4
YEDFr6nXuB5D9WR+9BUYlZ/ov6/D3EEE8svwQKvvTdU2B3TnDMuS7TMBSOUWcjiF
stbTgnJ4tx10rOJzg+PiaQ8eTbagSnDBQB9aCG7Nn4jz+4UfV3m6L8gbyg7ktcgJ
Sc2iV4mL08D4f6RETkfHXcbCeqDY4Uv65ASbdeKOhFLWT+gCm0IWCy2/7K3+9uId
mkwoCJ2iT5ZAD6Sagkrbxdl0ljpPr+fiWjD413E3Yo59xo6cx7iL/rkaTgE0KI20
obdUH4kDyHry9tWizJR7kXdSirTZdzChGxTxKdJsO2xgW7yFvIpX4lUt4yQ3NUXF
P6+Q9lPxpxO67Urom3GDb7FFvBzNCxe3eqH5r32U/q8PFFeRV4o+w2Xg8S2wljEf
L0exx33o0pk7IEi/dZSoyOjE3Houab5Vc0D7DYKtALKndx9exA2hFccHrX37UbZ4
Gsy47Y453dNFItEUh6wiFyD7mR28TWOJIaEYMsl9MfuSc/8ncU38E+1+jeTI5OMq
2L5A26sUXdilarr9NGQ4YeQXSBe2QPTIBchoTp7RBSqe+jEZs/0PlG+4jlO7ngF4
xZ9r1zd+8IjWsSA+i9zFbMdNZuqIhbiy2dezO1hjkqGJVa4ObuLQ+zG5aWMKQjgs
LyxZxM2/wu3x6EJJNJ6BsqgeHdF3CMRc2tKx6I4ptKoq2sIO90O2+o/u3BDk7oS+
9jQZGj2pS2WdTRa6+8sxMJVBWzE3vG9p619EXoGG+LIO8BGxFlDUfsf/PlBmCvtn
egqHRoxfBvCiveB8tHdKzhEofgxwpF5Meb8WjuWDyI4RbS2AVCl//C/K2Lphgz4v
4V2z/5JUiBSkgmU2tjoZ4PN9BCfedDn5G84imlut4TTXQvF1Mci6tN3FY93G+z+e
9uC8aQkIJ2wTiX0RfDvebg0ER9+f+7l/gCX6zAiYUh8/nTnn8xt/Wmc1QbcAgIzI
PjkXXktJGiYR59tVuPjlsPVNoSGRu3MgYeWnJbazVu48jwHu0FHi7hTc3deie17c
2hbFKqcRIsQNBM8jTtS5fJUTHcLmsD6VK3kREosOBGcOXUHSoSnPA9IIOtybP/rU
xdn+TBGz5P3UfoBreDQ0V3V65lVYFMEsINZJM0rF2p6HDMYIYnX0DWmECkeZ/3BD
GxtInqA5WosB1kDhFTDsfpKXmerTybST9ZeypCRw1vfwZNLoDD1xJfghtgY5XAfb
OcYZmB7cQSPZXi2wrXteN2np5bIt3/RORS4FrSkJfMu/S1hT0eeNzk1C063Cm7iS
AutGlwgVZ/a8La9op9vdcHEUBVQX7gip7sRFB56p82mNSzCqdbiwgEYvA5lpJkZ4
KlDUKmPTODVALnRgxElFyNFi5+APqnR8s+URQNPVm/69bUj2kZu67pRWS9Lp2LDD
KpSEYwDyqkBf8pxhofDoAce/JFzE9a1osXRyrOgLJDd82RIjoa5kY63uZ4SYqjaJ
UrTMqXjfBkX2GgWW5HIhlNp8kHr++3nzT6WSLos8UBk0K8rLyuOI0RILrwVoA6en
AjEVOBGMhoByTq36CcpTpjUowgHPIhUsvY1DhiNAezzZrUoxChhncdSuN4uHIwrl
TBouAp2XVjdKE3TQ6etqSiO+Soa+Js2U9aQVAwGk0Gq/cGf9kdAGJlMhg8O1l3Q2
i1z54w8TcJsaQjvHNhs3MNZUCL3DsHTcPwwX6wr3dWdLBgqob4NAgzH26qgN5k6z
jWkO4PFM5OmBOmYlV0BI9EYFuOER06eaNCIwLA9m7La+Ao/fiyB3fmvRWXjAysGM
c4kay1BjdxlC4XfcEGNniaNMwnQLtiQBCk7l539fIeWTxMgzvDdaGW+AmgaDtQ30
tYereNJ94dNj6yrmf6rSTsuadEyZtHRWRTyLxYA9Wy25AsAxLcT/KEs1zHQru9qX
8X5sR4Y+wXG9V8cm8a6bYlmVM0OnrCNh4bLxXaJk2Jgcllyx9TvGqbAC+8Q2pyOq
b95XrdATh1NOZW/tISADIbghtbjTl5dc9JZ0syofi+HCzLfrEwYT0BEevcStJOSm
uRnDJGHKWFUbvMkAO6b8hG0NPOyrouccNDuCaO830SpYnL5mk+zYkf+ZhFxKyA8w
bAEpiYfAHYMlXI5ipU0DI9YYqCdmyHbSFEX/kEwjzRok9YIIl3BUT0Sbyg3VRbZk
1GpU1i8SGg6RRvHfipWkRrGkxmW7B38pxdRdYldNZ/pBmLe9SVVK5zmxP/yNXQ1S
Sq/UifxI6BDvrNXJ3iJWg5ndS7P9RhenqXPY+MGF6vBCzHa7NscelwKlCEG8zCWF
X8G7VEa4L8uq0GTVYm6K3g8PeeFnJ3UG7zkDHVB7rMWEMtLvGUaD48kHDTAn5z/w
DrrPlr0uNCXJxCVS6rFue+foF7n60Aes4DneWILJ1sXmKItW6Ad0q/O57A3rDuE5
RvhvfhRO1moEbklRteQF+JcrRinTszDTaogEBCmcvIKcuBm6JxSFVuzCEgJf3r9k
KecLgnlYquLXdD7XhiiS9RAqHaMNAXeFsQjJxiL7WNuTs2k2JawX+661Ayn7vAR7
DbOm0g+wvm4lFmYT9O95AHexv/cpfSdxDItSeisbSYueCXogFzUI3nR7z3gd0aRZ
/2RWne6xjzSX5DdQVOeXAdts7uyPwmHWQp8h1b72AD/iKhEoKMVLkZchA8BP1mbN
SXMu/RMsgXuUOzWhS7BAHbdW0euJ9JF/5Uyetz3GSuVvLRTQYTOrfY2bSonEbGXp
TjG34bhMQbZzW/6054yi0/01fFprcPRX9h8QyOClz4Gp7/OOWwPjdAMA/lu4urWt
n+A8rjYyjyQc6+7nREDaGhk96puR/Picb7tnvsKdyTu/TcAKk2Lv2heGX01TH+01
2Z5o5PtP2tmm2zmsW/qXFHvFVUoINAmKuxRSSoaFMbOgQ5pve/XEaO9xa1GqaUMc
4jKcA18QAYlQ/TPo2XbFYNHwn+ynpOrqUEXnwA/jcfzLUqouBDTcPGMIOfyJDZjI
KLsZe1VvcJFkC44DeSCV6I2cM5FWx85pGJlD68Yl6LEEY58yFiaINbCi72h7z4CE
hOrdVGjkjL8EmxhezEiNFjLOVffvejO0s9VJtQqgy2dvW4EGVnLJnngDPjW2FCYd
9naeadpF6ABbNwmKEXJQGB5eMjYuHwdForEfdJFiXpe7cp5wPzkjbeH+F1oAFi+B
5ztB+BGbANSRXbJlMI4aZVkhQWS/6MA/73P9hX+Da8Uz+cwr2H1Qf5YmUO/AIk8Z
Q4ilSQIZSmL+ceKW9iiL60CqBP/MGKbDUBmNdFPw3xdr2KxiehuZUt0a7e8GyShe
PtwlimPF2J9MKlDG/IJskkx26q0dfxnCH+3lm/iA4KRAOfIqHULqRRfUy68/OF7/
J29hCOZvnq+wUnAElNo7Za5rxBiHC0fz3G+gt41pjs6+HM5lU2dnfJqewMvqy1mE
DXslorP1Ewu62p1Tp1lAWUv8C65f4dDNc3lc7XbI+H3e5/HSz/m+9xCvcVva1VTU
lfAgEQDyYXigzmFxNl9/z36y0eg9yrA6O1HSS81yBK2YmWKJesosHlps71Bgq6Te
YomxxO1PzmE5h4sSXJofK2kAA4/rjYxRusZwFvDXaGZ9FxfpKxEPttaY2oiTP1gR
kI6zsPIU8Kkt7vx7F0TvXn7hkSVHC5FGc+kOMj/hMFDw3V/e9YrYLQPhFzjZ2vDU
aG/bahJwqlrWDLi2m9HZjqgtwwWxVE9MRXFp+My0MWxDL8z2Gma7sVPy77Bq/tEr
ihZCll7z+ljbmvjYqJUhJEQRS0ujY1R+I9lC3YjJkr2ly5ODx8ElCxoAhpe0Iv3F
pHllblNxJpJsBhbRrdY8Huu4OLotLSjazyElhPA0ml73ipWKKg9F1OyGBcO+sgi0
L1VQjbDmd2OODHIXDAhRO+In63+q2QRNxfYeXlpZvCFVW2VEkF1mzpHf2he+nuPo
8s/OdsjQMekDHpJHgsLRJai/AjK5eHuCqqWLYB2lJ+LnZ3cmP0K4ZifIGjvui8di
9SP8A+xJDv8+0lmsuqQVC/W3AVDGhyz68yKa+6/cVDxFXRPzEthb2FDyosboC3az
4X1tfOfHH4xCEbGrnQqvxpHKH7GfrEBMh84Ne13+el3dGl7ZIy/699/SkG2oriWx
aEjPxhS2qroBfZQuKSXJVP2kmYtYeZCcY4MaVbbyNDK85Mkg+x0cH0raIHfQBoH4
BimLVC1PS+2AdXsfcCGPp8gtLKcHt0Sriipyd9JV48WHlYKtzWUUFi/DJjMiiHks
eff4S/qU9YiQPqa1N3ympN+8dqnLmvyj4lUK5Y5B9P4Ji3WiXOF1G6Qjknrbt7nw
URJQxsZfF+O91LSbyzkOybw+tv1Jl+Lmz9zbzTcRlWh0ZgBKJYygdp5PnOF/4Zov
+JVdLhPija8PeQUGjCTgCvOj5DM0nt3YPi4nXfdFteFd8FTlkCHnlLqqs8LHUkS6
NgAZhv0phh06OiKunqqwpJxm05qF+ZWzwxz4bhaOkYS+IbzEUqWqQ/1OfTi+VT1D
HmGw4JuaRP2mnAjNOz6ynS12Qwfv/p6vyFwfeQj+2K/1igNaBV9+LKzM5AhaNdCq
dkK0eMqaHxBl7YQ5rV7ABs5ggYI52AtB2B3XSgRsXtp77bgK2dMxOAUBxu8AqrJT
luXdlmYtY2eKpF2HDUCt196SK5NCc44MLi3pF1S32bSwFHjSvTKDIqytx+HQgdvQ
mhPytgdWP/QD/zOT3E2SRYX6YmgM98RjIU7jAepROwf1kgH4g1Ufo1YvSPfJKHxi
gRZeMPU5xcBNkAhHlygmYqKEf+kn3LlPgwTP0DJrE7y+0LK+TNpwReQ/3LWfAKYx
VtgWNZJdY5tiDGUpQik+8be8JL2PDoRDohk+mHQaQjv3H2B3wABLWlOxiaoKM3V5
7UcSxAxd7ydi7g7Wx87JxDtaKfnWbzr3uVqHSztnk0l31iKWu0efUHB3wdqoaxxV
/0KL5FyxZV0VEbnEh3NoOoeAxiNSL/wJhk+x4GaVllmCrq2a5WrDUUb0601CbpQh
0y6ftzLsetlPGl/3sBf6uGUuqN7Cx0gfJV/1qp9UQvwKrjG6Ao+2oD0m1Eil/j5+
EwklxCQk6KBC01I36RkIA/oBEtJ5tcz+zv/DXwmocQ8UNfsqCrATdFVGRYWi277l
ApXnRbytBeSU5VIFeaxy4LYtmjDndi2hjMzIbCxeuf0SE3Iwq3hfXD+ec5nG0UVV
7TVqW6rlLGpLbXR/vWACqYoLxA3Yz0Mi8fR37V8iaMdeNW84QUNGSC7e9PA094OW
pcOLrM0Q2bjnBUo7jfsy5ZYDOyRi1MnE07QYOpxfWfZNB72Zb6Gick4Hvf7eiRFT
WUpSjhgb/CdkzE8QFPbQB8XiitXK/35eyEJ3Z4FDlqjQBPHw0b2DOVDf8su6Lx0L
UapSO52VBPUycK+4YWu7rZ4hdOZ28xqppI1U5JeSNKDUN4ZxlVKlEGCIuFvfwcz5
NR6/saxbi0dA8G0UjJ4yH4OheEVuqB+/mbZyX6XQ4Rcs3fe4YWHDoz6rq1vzKWia
aF9eVXKMblPhBSpCBWQxPYCz6fa29fphmImo4ikliLrkIwKI2KI/Q238RILTcATp
Rvn/cAxDZQzULxlo8vmCQeKBhyFkTfH5PjVK9Nso5PDlWtmGRDB7hPdEQpcHTcUx
0fs6w0ca/urlok71tLSDAhtUSR73tnFVG2MYkUSQjv2Q3TD+hktBacM+/wKAHRYg
IoM9A+muyOCvXAwX+CqmKWnEuJNhcs01M4cA11HH8VzWZqUuOvJKn0zje0Jk605f
pAJXq0fPpWw/D+oAUwhQFd+BMCF/+5TCkhGieG3hsMYvyH9X2r9YfrkUUTwkoIKQ
S4g8IjVdqo4jwFMxhiNILGo5lDUigi5t+tav1eBeXLht8MsW9hdvHQPJnkv9mGqR
hBBlCoqzk+zixUgNelZ8dhutx1HwRBXw0OVN2U/FGoD8rbeqnqi27Wa3+u0OzcWj
N9ohpaWCYylEgmfaGMosmaN8SFUdXdd21Tb3yAGoV+NzPpBKW+Ae5zin5V5BCDYF
I4rKpQMU5pcbag7klzT7ojPb6zDW4rUt+46Rbh7aIYt7WlrmmTCMtFkPwH91MRUR
kfpZFPHxHgTjQNN86atxDjMOkJb2NL+5nhQkgOQEEIgRGoSIYcEFQIkw+8SfG0zh
V+JABH6PfbRm/gz+4nG1kX+YFGqnrwH8GbF7uAb9NbTys68K8BvN9UiSKgmV9Uxi
6Z0WbtWVeuHFPpcQfMvbaKvLsJVVenzDd0zCkae3AHgIJ1HJLlfdoiGsnHoojnQk
hwXxzusQpPU+9SbxslF5wvSM7gfZLufZv4+dLkBNfj5jdOKaV/3vBNN5xvvZfQu5
4VTklvFYeCxZCY9gDQAKqec8ry/aQRN/XfOuvmTWlnBuX+EozTlpKEKqz+ceMzKl
uMlKlefVTIDUCrSfLSTo9Qw15pkABldBrKsUtiX+zPXJts0huf75IhfKunygB4QF
gZ+7US+Wy8nx4dUIWz+akwdTToQGC3+VWt5+8QqeBJ4mjf+ZFz5BrVcfw42ePEQs
2OARSPVXkz4sZg2/xo+bl1waYVAqDObxltCtwsYVFReVXgkThMPgNFqLbrJBkcgp
H770wFh7Zo7JIgfzPYQzXubE8TpvxpzBuD++WV2aeWZJZL56jC9HYfDGzQHEeOzv
KxJdfq1yrrB1ZPbLKOOOCBGG2I1VkW2ocVePV1MLRXvlr6Jixoeolqn4RJySff/M
bXUnJ+5h96AoZFOP/8+jbLtme3med3+/yJd5CAXvB2tLZZMb/wAMe0Ps+fn2n9EC
FFuL+b+e8KO7XIQf1yI6vlhaKYrlsEOFFz5dulVSOYrJrsrMIIwboGXUFc198Yfc
o0BGZwgxCRC3SNAKlY1oUZYgcxR188iD2DemPpouuKhYqhhgiF3gJ12+isXee57C
JfpHivAKN8KwVSrXDbrS1mnksE85cGMFv9dvlYozXRiWkD/0FZSR9I0LwAws8hrd
0RX6nt5USbM2jGsQoOUrl8ysKDt6iWRmqR/7V1qVK9YgwY8HzufMo7ETRS+bCrKS
xpsI7L2xuEw0SDkjGuc8eVvO+Nvi420zycMBZaNiRhjnJRrWj2JIuNvAl2np5NT2
7BzumrqCfXXdGXkGqN0dVBIJv7j0ZfeY+Z+hMaFa4LVq/PSsyLqc1mf7tZz4w6og
gi5/+kfHBE/mAyvbW0TsFuqdevTKAu6sCdCD0clxv2rzxSDZe+g5ZSyqCV+AKXug
1LqFj84rofJlnrMfjrzQLYDGX4uAL3HsgCOmBAbkVzMiR2KC6c4O0ouheIeaxtwe
y2YL1IMnOWfWylpztR62VyjnL6/40+z7xO1CuNkrxif6PR1RgBORAc3UT79MvDz/
8pgemR5V9d48YA9gcHiV2mtwW1UrwYC++7/R9P7Lr5tEsgwrP4oW0gns+ABIti4o
de8AWZi3XYr4JYPHv/EEW7jXhEaYGWLbQJswLdJycf3p7hKRJGYeShl0MWM6KVAu
4PFzYuxss0P6fUWI6ncuJE25eVZM+0l22OJro6aUiWUk2NT3R/vQMNyBe4YvExPH
n3kPd9YzL1P6LWAQCkh0aGgdmKQuMAD7IOPy0HXf/R6efA+PYhFps7IOU7XFzrtu
GsCvXZAR2Ma6wc3EHmDVyheL1UEzXxMRN6/BXqemYbtcKKu85JA9hm/wYNOuRapu
JAH+OvkTNiS3Sh0LD/5Vbkv7k8iUussmY93GeXpltDXCGrKQYIYb+Kxba0Gq0vey
YwkuIgqHf8eANCdrIhwwdDFWXjMjs6Ok9VRnSwmtn9F7Sn/HlFEWIvKBrTxsq9AQ
5saJRZ73eG11kuAi5qvQesBUTOvNSvxsa0eEli6VRobNOtBeJs6f+rC4QpKEDMLC
hTK6cwjdHTmOJKppaXUjSZM5zCQcdhCEv8/5YiFBhEZgW2NvcTXecWzEmia28gin
k6IELBzAq2y37QRkc8QBFEIP1CZm5COun6Tieu4OxfGcoVEUyVhk2JlB90hB4rYn
j6MEUog3w2KhEnFYcXSwGmgMrvg+7zhxEnzeY7e4WqIv49MCW9dQAojAGG1bj8hr
HO6XjXW0XNivbXgsM3lNTf8pvfOqvx6kmmhApiUxU7wj17/WYT/RVgMccfreTApe
QH7d2NYl1l/Lekk4fQk1z2Mwga468BVrYoD42h6z6X32RV4A4+SODS6aSoTWVFe+
fQEVfv40MNPgbqENdtUzVu1JASHDA7t3ep9u4W0M6VFIIQSgdcHxg/w0tqPdId9x
Hh2rmbSJeSx3YQzyqZsdC27e7r1GyzKsUb9d+xcSDYiZw/I8OjJXWys+Bo/UFR2t
C9R9jzq+Xy8mZJ5vC71bhCSDmX2smz7i1ipKRaWYtiLRlApP19acuS4ef7WQJ1Ux
tRkhP3Uq5BtEZF0eUWjagbo6R4mZEpW7pMjWRqzCesVQRCQanGJon/uv8tliApcI
clJ1GTa+ggKyDErPahWLxd7jBjC0wpxG8dCIgy+xiTkZMOCc3xqS5uP+fJYCYyqy
lhpFdv9JnubncIRTwQOloVrUTtVJ9KaUJ239bqdQluQK2phgqVwZs3nhy3tpIjio
93nBadjG2qY8FFZYd3bELwoeedW0cx/bCJ+2/wOjnuAju7t8TzPYw8SxBiLRcnFC
tQAvsg2lRAHPmcC8o/ZGbqPLpnbEShVHsbb1uZVSxxVEh1eWmAEwsBI1m402wQ0y
JL8pURv80G6HbSG885O0RFUTPiqT9Oe2kmq32tK8piLZiXU4mAmvDlCCnqRbK1T/
On82uemtNAb91nQE3JmpSmpQcv9GUbTTxwWEKywWDxd9U/6Vhv5bu/126p1rjbxf
pPRiTA9TuTHBBS76cl2n/+3zceaeiYoGtI4yIVoWwSkDHeNEuxuUh40UipuTjtIW
G3E/u3Y7k0zvlYC6QMUS6nYgjIQBqkbn5J01QSV7BiLWY14Q/PZ2bJNLV8VoYmw9
YSWsGagjjF2DiioYqC79/ShUusMw4HWDTqoAt3tD60JvfTxO+/9wEmT81CRCbC5F
wCFENRVh1S06cMfJinFVSwvid70yO/njLhQHbW6PsycTU4PzRvTfMxaoMD1pM27J
ps+zPcpoFXDsY0aYI4GMWXtSZTyQlDwoDpC+XhHnjcMgqGH08ur/mZho1ldQLly0
d5qqlxE6xKJRmIeJIfyChXIpGp9y2iRVx2WbwDBCU8ODz0U9IVLjydGC6lzDrllG
K/Pw5kkRnQG65fRjbPOxtDSes0z8ADBHW2+o8YRFm7CqackgkYk5/2yTVHjObBbv
XKUuuTPbGkkUT6OEBIqygin0zW3crld1ia67oyrm8Jw5TLvKQydplMjK6PPJPPSt
1xtXKOqHRWL8jDXG6iM0b4gmFa1oY4nUGjC9Wvyqgx9jlyzacBr1W3XhEujZgW9a
RLN6N8ONeXxViOGBHGw4GSJyGMi7EkDFuLLoQ+WtUszHQibSmH939oWhiW8v5y9r
ex3FJyIWsCy7pHVGeHwgwmO+lt0ygci4Q9goTk9lefzMW2tr67vVNhxR0f5IOXUF
WgDF8/C8hMR2tssX76JfYyHjKUVJY5UXvgBvA1enMAWXTxPobDw0Azl7AjWzvfK6
/ocdTIbZ+m+8f2wEU1qKPpfo4wSgdeddCjiL4gKN141H+EXi8R3z6F3R1rflcqNx
6kTxzUUbEfkMIXTZ40kkzOUmOGXmN44SPPURmG8O9UXcFNAqKPa+qkNtdbP2hGk+
etiW6O5SyfbVC6Hws8d9G0p1quvWtW8da1RpDKLxmAVpm8k+USMeRBtoxwPsN0B5
qItYx1XQjElBtItMV8yAJ9h3OmdVITRNpoOqvB0h8MqkqRxAr5fgZ9RKlH8q+qDN
y0CCxVSfcldeeNqhk4AZpjDSmZH9NVT6y1+QGtpp7fVkJvszQSkiohJH2FvbsHwD
o2/m+N1vWWUDhT/OclNom94TiSu/LjvYewydm2n0ZV44sjANMWVx0B/5kmdCsV/n
4DJpEvsvSaxfq0pL3OueZnKYspx5eYZDCO/xLFn/+L+mIvxmnscQOz9xMFBtqrvJ
ie/3rQpA+J6GGpYSAQQInuy/G2NyfVb3O7rBc5VMmyVAt7kT5ugTfprihYzT6+TN
a5PjIlosj3LgSglPil9r+Jc8KgmwjQyaI6URf9znUa7WF4kDHIUdbrSzXf83UDnk
CZEGbw4AGpy8gYJPML/F8stWmT4GldFPK/bCPPK+lcVNU7c7gX1oaGEEcOB2Shwr
3SCdZbp/xDmE32ctI0xk9xnS9219H9PAkt5uhOESYqlXFuUSrsUllZp6/ViUQ1Um
aaGjKblJ32mCmW1uo9t8sJDtzmP7nBPBUOiRJ8g/py1KvGffFqLlzzOzmU8kIveu
up0zxj7vyJMtUslJRu5UHNdVnjizCnnDyeG600/AIjgzoSVhP6wx/HLBllynP3Sk
s5w7nKpPE+5q92CL0V3g+wHqCrT+hp/q988cFlrGPjHLdnlPs8xkhX8PKvVlJD0M
ejex0ADd/q2i4X8NfA7VIliFaKyv0KHhUGmI1PEXLkEBQeyB0tUHRpTXU9CHxZXy
OpMZMHgDrWrxEEBFHSkbiiQo20a7fqpaF1JNL5DokRxdq+S2nMTO+BgWBz4M9vP6
ba9QICnbssp5GQCBk5Fh5UDHg5uhQtbHtQcTlirXyuxhcK5/DIoRlfDQXNzHtjrW
Ci8zXw1cp0Y1o3qQRJYZ3a5dxlaiKqR0tTf+29TefSpZFCXhJ5mskmyMctIdTb6T
ZlAGkOalWbbXfXt8Sai+j95iWGv7qMxZBAipuHxXL8jDcqC0Xyd7jH7wowqwKtPf
f/slNJaFYFEv63F6HglgeIwM7SsKOGLWwITTJ8pR0KsIzhepwten6WI3lXITePOy
qcX6p/VS7CZRxmjAcS4PFxSnlkFxgOyeWX298aShyEk4B3aY4RvJYfilzNw0DtR0
1D0gkqqhwaK28f6mWOv83QPgIzVdjrpvANDan3G6Y9ZmInPblLwNYUl483qpYJAQ
F88GF5WhDeE2FZVkvza/A/I6v4+lwdJFSIhAnqCy1K37UDTK81fR09+T4Q7FR5/s
1TaWGHzM9tWHj2/LKin08AQ5DtBC/1Hzgn5vTpRuzDszCRwF7Eq/5rFk+xc3gtxb
Hs8F2C9+ZAWIvOUGNPty9aBUjQtJ30GQfbotPs1ejKSX2kU3AmUn1ZTc8tmFyb/u
6WBk4gsk+ksxf8eSaEY67R903AYUM0PUfzGtcrmatg1ahxV4dffqR9Yemc5j0XWu
InzjfkSl88lj5XEj0EkV34ePdLL7nw3BzXJ95kmhukQFndbkFBsvA/6cILuifkwp
1Le0TSziD2+jreO94swJcYcFuwss1RYpgKutmzYo+5bNdwLn660Nspx6DVzwu1if
NFgo+OJAmDcWUl53H+jDiVx0Rn9f/WkbJhNJCykI8j+SnXCzYzJ0JVmeQzsps51y
ix9GkIMd9ohv9mZ2V5dqb97IV/GYQc+OT0/GtuigXUc25A9BEAk6XXYQQF20Xk/3
P2bCIwF1EbBVtju9teYbCxwN2aq4cxWKmlqz+CxgDQvBIAPBZZoGmnzDp+4bbIjw
SL5bhnxgBYh3PIGZ+bqY2aTvxkSHcZm3RDoeAlAHKhQibLffCSlIkkKlJUEmmo8x
9ttV0YLicNLjH/UmyPjxE11fIPG6qUjY+qyxH3LZyLf90GhTrTRDsF0W5QjdHefB
Te8PhKjbS3r8SWMgAXTt/RW1gSuxtXra8YnD8tNq4SKxBJuCGRdqyvuR2piTmzn6
fX9qaIgKBJin3j1ryM3U817R0vTJTJd1luH5fVKNkVfkZL68dKk+ZXXkCbiyTP5M
RWjYwF5NooVX5ZXxSIXmXPyuH6fBZNbY0FUm8dXUoSDFP90ddlGJk/BDwaagxHlw
pZnNClqGnJ/iuzhzq1TEgCMxbZry7x5r0g4vUtr7t+C5fbJiwjmjkP78DTfFEZSh
is+PuEyXGIXkDj7tIZTaW9v29Mr2+FTke1NOEOpsoTyLqbIPUi5Y0aOPzIYD2Aie
`protect end_protected