`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH2zDWBuK5P8yo7AX7UTifRtgjHPJy94suZmLcoRomtnF
tp0z/T3lV7uwuAODOc84OQJHwoo8JmkSHTcs6PAQAdE9H7oGeabXqjxQDqI0fDDR
M+nk9RmOjTzQjsGcenH/mKJAsVK+I4eYFR1rA0Uwoi8jK3CR7mwjichzKsoN/l59
gXqxitfp+w6G2cA+QbO81Tc2sYT9wUc/tYkK3kvps6dghC+fQbLoRHQdDPJY4jHD
C/czVXZDW9cE5VUkEby6QuNDSrMnSUxh0zRTuq1dd52ehlGwvaw8NQWOJLudqK6f
lNrx+kF3yOulR+IaPacR9DVp6UQ153FeZ6zgCuP2WBwfgm0EZUgiiEjVRc6kJexx
yYsb7zYPfWkZs9axSBp13Xk9FLX09Qv6jaXLIz9FRxhddbNtLr1Ra59FSBfSdu+N
RMeZdC1ZPNhJtXJUPbhoiEJSD1GVxsFRVrO2c1MvcIDOE5xm3DZC+yCHKxPnC/vO
tP7hVHCruZDn/rzqcU8FhKnwBHSokMz3suofCgh+fnMyhoo7XJglfqcN+4g1DLeI
LwHfLOyhGLfgPiMnqhbbSSm4Q8UKbWKJ0xisjYhPEWwCraoVtrdulcxK8ecEzFjP
77lyWkAeZpTv6HGch9z0z8jD7JIpSYjCQKBLSl2HFNanL8Sq6xsS89PuICS6inUz
6hP0Y0a3I1KBsl0xTxbBotpECJ3Ds+h0GgkQaxu1IeO2U9/jCeNiQdhfmXFu16/o
bLBGO06oCB+hqDw0rAxcZoepISWuy4VRNU2L/dCvnzI8mTbWCS5y+jIZhfLiZxGj
nwuOrC2jBAEuhqXGHsQyL5cyGY9vLrjxNYPgnNlfAp8Chh+/+Shddy3lHyCEMWwn
1dJ8sIf0TvQlnJN2v6REqKSkh3N/H+P/gBz7azTn5XEI2XzLs5ppLfl2BY4ceymh
GxuUEkBFDKfRA4dNKNfV0detVCDXKAoLka1d5kMzmvxqOPbjtsc+Wz0deZkxN5kF
UcdFIsh3Lr8DqWsZwkq7s8kb+hKRHM52pb9tyoi9C/0K8yjNA6iM1875gnlIA2cK
LWdVC1eOGdmnc4Uzwf9LFc6YpSsh6z9V5IetfhCmDKxnO8tdxGFcWOsM4UuOLESA
DnGAxlzSOG0nM3qPDhSMvABXTKpVVBWPCSsHTDwJSCnyoCjPY1yCJvokXHU1WOCy
11UU40sMEgQl+pq7LQJd0Ashifl0aH5pDK/Ag1zUrlxB9I2v5GxPzweG2/Wvy+WZ
K1ajKiK943p0vxtf+a+gSZRa6nkBVHL7xyzFQDsLfKXqbnZPcUsleNJttzg4W/gA
xKFwtxxqU09i+tXPBkFpCMoOoUUtl8L5WsTnDWi+7XeaGGKXa/BHDWULiDlda6Fb
pAau3jHhSWtWNjcu4xTE3iLykhCV/o16sDAK12/4LwRMRQy4GPdPiaHaF8GTwYN8
/JOKNghN2xRpBP2aT0J5pu9RlXyI4lcJ9jp1bmBLHGz/KvTe0Izmc14clKnjB5QO
xFVPY5OmcestQoTw/8BxkE6hDVtuUMRJSm/aw0n7/miHoEV/GMD2oMntHEA8wNQW
tmFgDapA/B2NHGR1+C28o6Fju6zafYbP+os2fwh88qMyoXd5OjO6shmRNngUfaF1
BRZZXADaTg1QVSnd0aiP0lpV8sUkpGZZ67Aln3VuikfB80J6r9vC8sW3gWxUtzR6
bK4p30rl3zWfYZpU5J9WMgO835OZkTKqMGzplC9b0aDu3Pn/4k5jr0doRbMIVVxx
RYNqLQlcAS3LE9/hGv+Ra/S725RWy4+01aPuFGB0O2YxFAf3nd8uneHg80rpEEVy
XYSkJh0x5N3utIpkEWdWHzh59IO0Ey7Bt7O5g/4owWxMMAVGXA64gpqifipoafPf
wIa453l3Pwb+YfyE1xk8o/uc3gRE26XyGxUuTHkJKu8F/Y+t1m1671V64ilqdxp/
bjBISCtC/Oi4J/fPjC7SvaJi23FQhlaL7o/McNQs0zEljcj5/C74DwQey8/ZcxT/
QXYyvDbXXXtOPEihpBxgyG7Ql1ePIoqiSW2kVwxramib9opSGhFXbwjauKVl6XdL
PJWHGp4szO/wTAb2i5W8NfyvZahg0EX9RRCYRRXEMJwQMHek2etZWtrumBzA8k8A
ggX2Ox8vVMI3nrQnwukXtc2zUuDp/TqGy/Mfv7M1ickNl0ZMbdUG9Txm069DU4VJ
gmxe7mMuDKqYtpR/pwqqIa09JpYksh+1IY5U4ceJ8+wtJEo0S0/RpzM4hcM1DXfQ
TjxpO5y+85N0n74KYN+O5tS3IJ5jVWcHm0jQ145nbdT84vTHGdXxpHcZq+9REMIx
iu9f0KMdXm4x/2MUbrJ/IpZp8DlKXz0F676G1z5A7DWbwHhDeIL63PSMPjegafZB
+sH3eBXEHTu4oRiHZeYWapIe/dguohlcWCebdPiGSXFTfBGRVFc06ySRWKjK27oU
GIYzxL7uiaTtdbBYgKdYjgbhX1PxueQCcxIDlAsGZJsiCXIjHFAFInBp+Et9nkQt
I2F7zKGS4/Y6u19fmVexIlqmcrJAKYQ8Jn0mjBmbp2d4Ml5NAlgb0cMtpPoUKQZz
Vf7EGjlJ9oVWcITUTri0JRXZYjiehqCyUdkLWC7cQR7Wc/gUarJul9U5XXIrUBUr
k/ub6CkIJmLNwqH+qfLHXWPqobYJ7OKb2RBPXlGNB97adamTjdylPKPOxaIIPbnT
ZCZ0008t2zTrv3+0gjqIItvaDDniQgcaVPN21A7UCPfVqeiteSXk+tQEVWLIHaop
Kt+3D7+VqXc+FNZOULDdZKIEGd1AsnbV4VDTjI0RCaJJvKr0B+ttXJMVxaq5h1a9
3xtGUinxTxTUkYPpxYx/pnjb9XiOu111SFgclvN5+wdYKLAF8wdukHy1L1e1fxDh
4aY90M7QtUFGAlDvQbvJyTZvfX1dZfChCLopCEgPkorduAI7v+aNYFTgGprzr0PR
bGuz5vfG5Auuu6Lzm5gls/Pack4tZOcr4QgjHcPAC73Wcdce+ZFhO8yWhoE7b6wv
3NDbSqwxba5lX+/yG6WtpAWCsGsPEXFsOZxodexp/m6bSI2dZyzVB9jsDC3iVxpD
UqwTM9P0CEjYNyPU6ODjoH4dH4KRC4P9WdrpUiqtf4FXOkUoZ/8kpChUdaCBZCPk
IUAvQhXKm6rhK+Fj/cgB1DhNUH/yoEk06h3pJuGvqVQGWnctF6dA2GKXuemgwhlH
VdMeUldpq1GG7O1QKuLELEGK5oIdFP0aSTH6xa/v95UMLyvzfmLJQ69PTzKqy3ba
xLzLLQCQLpQoqMXGb4OjKIfspDRsfRfXRyrFBwF2NEkns2RPtjDvw3ZkpS49XLTM
7rxnCQpXRShhC6AeHUSixs+nh1m9g2rJHmepPjk+3qafJODmQXxkA+ohDHvCfv3Z
QTi9jjm6MwKIjEw4XU0qHadiQmYZKhNWFyY4eX3/4QSiy53HQLsx1l8ztUg8KYLG
nSbxMcJK30VSJqqK5MOvMF8bXM6nqLWomhds+4FYhtRF0x3uRQRXHJ55DFctYE8i
oIszlyQidEjUVqVc/0ktu9FlK+S2aB4w9EjHwgxjWNG0SgAmCs1edu5IezwSLhOn
qboSPfrC1BocRS+UpbfUK83XL/NVZgyoiIA/EHkJyLUhUpPyAxYpPXLHEpaJBv4I
1sMGGEva1rf0D7v29pTM7cJ7G7/br605/BxU0LO40w+e/D1uhqEawwn9IlNFYyQe
hMY/grKpZiHIQEc8z4LSVMoCB6bs/FXHrCejc3WQPljmxEWquaNGa5AwmsnSAihc
5/eFyUw+4z85IQg1UcVGDcdCIzpPQiT6oEgoGT9MycbhT1qsV1b94oqinuPx9uqL
0FCwjpd7FK++jqyzd4c7WUUmlwNVl3oqPDtkZq+Euap6bFBPtlLNyGLxm//qxN7R
zKGPWjfPcEIOKZrdCxPBv/oth98hNxFL4UI2M0pJaOqmCgmoV5NsSVAWa086Ocw8
5KLkUqeUbGOmriuUOA6vpQKOJrtxED+7FokekaiukSk88SPjlhaeMPDZ93R1BMIK
Cb5FJKBvXckja6ozMtxIaA09VPl5ZEwpRV8BKkirrWfRisOjxBZ8+DcOVB5f/+jm
nBI3v4mwkMkXBZ9GA2ZKKRKFU8MMfUnw44YW6b8NQKrDGakjnyLFsx0PTCHeK/9f
7s2ErZoIj2xYyIM+87GlcLyYrcWH1HvDhSXhtsY2Ce0Z1nFfdClQNY9UKt06XuUg
euET1Fslh6+CW7jRBD7d9n2vpyvL5i9btsXnkDcOTNfHNghMOtWzZh2qpb/oGA9J
3gD8oj9ssU7YU/uRxhzDjx4v7LNUzSNNvBjwGpw6H6/08jQ6RLyCVA1JMRZQK8CP
5K/y6MKUEsbhV5F7igAg81QL1CEoUrBmvKvpzcTiIX0ap8oXOKhYWhIHgmw35L2P
tNR5cw+CbFjvpON4ojfWu7aPTct65k0gtfL+hbq8/8Nj4pLyQtqVrJGUgrT9+TAp
Hdi7cQ2zkK+v4aI/HNGwEqDgjFN8NBqTPlkPkaaJrbDERAd4MjSu2oNeqeNdyhl4
z/AmsYMQwuZpj2VY8RqAsZhJZbJ8Z7yPLEEd/fuTbNoKkTWnSICh1E9eeSSOV5xq
v7vBZr2OUOtNtDAZXX2hmy3XB2F3AeiTuJGtzzYrtBVP2IHXdsbtlAwG/aKGg7Uz
oTUs3O7szGCCDa7P/G/Fu9ApWiAC8bPGI8s5Znba9DynQNIHDJDXvsZeVHd2ngth
0DDTTtq0rwKiOhb1bgR6zhfaBvMCSnDW++2kyyKoZML2pULrshbAlpF+ZcjH9Gjx
pNQar7saSQVSSd6SKsYzeJinC19ZLZVcHvNXIAsPWz9uu2fZQYUsdG82OCTtedxX
Hd15riK7SDjL4tMgMpMQeIWslcRJ0DMYujg5JhjOs2k=
`protect end_protected