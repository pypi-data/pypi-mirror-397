`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
ESp8jRyPtsiY+Gb1bQiTICrBDGBuaohyJmfd/xowZR5jiCGpAs3wDH0hvN4+IMSC
tmuAjiFIOwnaYhk37OifpkxN4jNqtaAfkiqwvX4bsKyx7O8i8Cymvdjt+FvXEvcv
m5Q0aY3m92Cg/qgi9MOqt//xAL9J8Lp9zbdh8quH/eIIcPhn/D6NKD2RZW0+PoAJ
jQhkxg8wgDWKqlnxb6WuhxrRij7kn5ymxJjn2XDIOLdbCgvq/LgZVRSnMZdAbR8m
U7UNb0iiusTxoxnOlnZ1u0aCaxvaI3Z1EC1lDYbyfjMcn2RiXpm+HOBATMm+UJcv
Du9Lg0ZYKwnD5txQ46f1qQe6KAi+EQqHKYWpJKtT1HKVy+b4jXjLQ+n635XATDTc
XV3eIZD4NIEC10MrD7KX08Ywko+6pkC1c+0gwd5lqRsn9q0ykXIMMiWMhOry+miP
wuOG/5U3BHA5LTMpkIRP2D84U/Odx9LEB+qIEQHKJauDQLthlCIEqtVgwQ6u/znr
/oT5Q/KJKb9/9CQmIn3ghUR/KeAWufXt9E15ZP6+qJ1GPGKljZR9vItQGSp0Eofs
7nEpMd5KRUuggJab/sVMXy6tvAVsVFChtewIwnh4lwjJmnqazPBmKQP43wPjPKhE
xzu0lW1T6rwZuLkpmNLozprvZi3j5HcVUq7ehT1djWzZolSpVHkMCGJwokpq8JXL
jvzxe5V+Q2k5zA3RRkglOl1SrgvWxVwT3gb+EPufQAE3nlvDa5cR1d51aSQMpe30
EYNHygGCX4cjoTXpQFA4zOmcYrCsmFUigIkXMe39xR1TXIG3o4ecbP8vB72243H0
PSoZa0NvoRerhfdQYm7B0ziqdPTjRYhtS8GPXc1wHoxcj0Q2TnUoICyTw6ThBLRT
+sYaqLkFM7FdGPWZlalVBpRgDqTpcJUKAz8vd3MF+TEu2VGtCw836Ad8NqecXFJs
r5sv4FZlUfFayh8j8mYd0P+uZGLQTKYAw0FGM3FFwWkJz7RmN7Hg3iqxpK0CsprO
mEVJqIdo//7EFn9oENzqunujAOfO6BXD0Cj+pCHpkOID0ug0IQrmO2NJmBtWTO6H
Z0/fn4heZzqQTdgAEmUcyarIGzgGxIvZ12HdONsI7alC5oRZdKCXftJPFP8egZwi
kz6M10GZXpZmLYccFuBPwn0+UEIfzd4eEZ0S7ebjYXR3ZGkq7noe7CPuDF7maRnR
5fQu1eC5gOR/jgz1+oFrx9XCHZL/lxIv76obF2Fqw1/wT2o2XnnR0Ra0WwGleE2I
RxpvSU8e7ZR6ZK9NHPkmjDCK0jHvph6hDrlaiXYzOygtFFxiPjBecF8tdgteaF8E
JOLc3BHML/eeN2YppD5O+gnwSb27yZbOi0rwnqwaz32j4X5L0PobRtnLFPGUVF41
h3gY4X+buOsHwlDwaSJcrxZT0DukrTz5QdRhNSQczj9D7eFiVq8q9jIHFkepm2rP
kOLEX7dBRQ6b2s9tdvAkV9iNAt8IycrzyXTUO2RFHaQUo5z6gPsvg32GFzDysTIn
Epet7O9th0Sda0vTSANF3VC3Voz+RwpQ3KRNZzkvVBenI6LXH0paD99l1JbhmiMR
8bZX9tZJVIBwuFeh7zWMt1lJXGP6/qaWKiuXqXApfSHeY52M87ELSu3J2DOwOwDW
HgGqUE0EVTsMd/2Xo7MREjjUMdsTLtFGNAmWkiYoMrb1LYFucYHvE4uwVRzpeQdy
26FiQzUlcC82s/1JAPy17ge2/cKaSeNwmX6A7kV0MdyWlrIFgZ7gQoFsLiKlAu44
l3QoYwYlo75JNwfObFQXSftwSvcf6Dv81/40cE2+YmLAhN2sj25HVOXiymxcweLZ
Iq9VIllrC8JZgOEJNhxZNe4kUfpTvhhebyyRFjJMb0Yvkk2z8sD8dusoh67yoam/
SU2+ZUX+a0NJVHT9wbNEeTiR2PcdRhIP06LHBeriSzRMqV4D+JZC6edn6KLsiWBD
ncEUb6wnh6f7BfaJ6Wuz7e8D6Fn0xOqY1a++VEAeezGnqwwagUz2iBm69AsfkAvZ
o8zRNDlkPPzNABMAeIB/MTQ42426ffoZvEpgnrccs/excX52JtKMsN+yRW7YujJa
sLoCYZoAGpf2XUahz/qBBD+N/o6YYfCvQX/DXj3sAteGZdBoYtZytf0BxbSTfEzL
isFnKe3Pj6Tz0eLR8oNaTvvC3lcXjWjHQYmeP39ZF47uZu6rTE+n+sItYZBeeXiE
5Mlsja5QkWTGupywZa6aowtAFxlZPaCqCy8yUte5gl59jrd3G5L8kC14k+fE4QO9
XlLN9TqXYYpICVI6ggkIeaYzEVNICjsvaLKpOCC1kMlT+WG89V9n1tdZZm1wsg0R
y1WJi4FcFZDK/j37JMUiQWxx91QFq5sDV+jyH/vnvoQbSteX2rh1iTwE8Usd4893
9aJx6bcrVtl3o1sMh9JkXjt8NsHSO5JJEsR5pEZOQeqAA4PgWoyjuyhQ6DqzZ3nS
1XQrGoskk5BGrK3+h0XRC04fOyTybyEAt/l5pGpXuGt/CLSGoH+37P925qtcueUP
DNNVgULYTXQiPiMoLbZHiXUldu0rdasyZJKErfrSueYxFIGVbSz73OePXr4kK5Qg
Qvm8j2/sCf+2dgkHH4rrWNEEjSGy0/1K3WNcgRiEXuCKMfI6gSHhLpFCIkbq0u3o
5pkvY52ivb3y9+r/wSQN18dJJ6677d8yJ/YJhlg/fvNvHNRm9PcSAHB9SKoDJCGx
JNxRz8OkHindhkPU1B13W5ClcvNaTTTkeaPNMVfQqW74sFV2rvZs86wxlYHT2cNq
j4DDG1MHTgx0EJM4SE98pVV3oRk4jbaHQZuAd3PZOyv9NRUYiO2zzWqpfg4NMVuI
FEv/rQCKb4jQP9oi5SSmiAyttI8Lno5VreHsnEGxr0ZEyXwBmXD0wgzIc5o3b3Yo
Tk/ZeY6BlKVyS3eY6DpBweQzQxjSQJMeTSUX35cU82t77uYoeZIjjqOxexEbBsFE
3vTnck42KrRfViTuBUbyNGRsnFkKqh9eWUkxHaLOuNhigYlA9dCPPXP6Dt7+VWBU
7D/MwJdv/lw5C1mDLOygn8BfGmRjR+P9cWnt6Ity5dpX/6ZLfRq8jQaCtkCjlWvk
+9zz9Z2j0Mn87YTWsgFrHvHUAgEtn+yMLxUx8XItA3uknrJKiaIEFSHiQfW0Hsn3
e3fAjJ1ZUdtTvfPwrH+n9HftynEX6JCGAr/cAQCv/Gd1qovZeTtqtdcBYs587GnA
wAHSQ/MNmf5RFELVmi+eN/NNgZxFXEaExFUi1STX5leEII2tVQbMcml/DhbCnf17
P2yaorBODhuID6twCCQEnArs8w+s+sxQ9A5QCSyxXOyOf8Hfg7yOtloqoFuCexYN
g+IjyDUiYlVrrptyM6eakSDy+AYftD9uZSjGGoBc4o8hSq5bIVGT1jcvT+87Yljw
sdrHOv/5tMqSnw8W8owY9iprGTEZgu0Z63pCF8+gc8QVBhH7MWexS6jPDU/gMCRm
kIa9DF3YW+Q1tO8X4r3sSymPOVO19E+GuWR3AJkcrw6cynmvGk5kI6InkxSB2EQI
isnhRcaBl3j29XgjUMOSZBrvyW+IaICJ8fRRkmp2zkOXlyE0gM1uJIWw7MUNlp3Q
4WKZ7FowuxavsBbPOMycp5iEmIIf6vS/8FhGXp5BcUIe5hPXKXBG3jItHHXM8oad
21TRh8jkNNqTS3kf+QxYrItrKJaUhGx7ryNPeStOakBXYPT7hMzHhMqaSEE3TStb
UOFBEwfMMXUfnGFmHJktDwScG4xT2HuaMUjPcSHq8DJyQKPMKw0TQERwT3OA8x8l
Bue/LjNpbCNS8DeWDQXTIxkC5SVsWtzq6amp8Cil1ZvyC0WGdMVrEd4Kr2O5+Sg2
3uc6gQ/XetRLJ5cW6lLnUA/y+BvF2Ji99dShhy9lerLFA9hFK11Ed7oDN3Uy/nGu
Jc/0L40gK6YtE1ndZNVRjmkW6mUPCQyuY2jtGp+adF7ADwrhJ2Q4itlU9PpsHnrI
V0KFQwpuplDK1EJbjyQs/3yctK5tdkULDlJN3J3c22etmVWygOE96w4uNGf4jmnt
l8zG5GYc1uQkYpqon6UIxjmFWIx6V0432J4LHKZaImGqOQDIws7/aA9uer9oaT+g
Z+6Al01ES/QP3dyVGGtT5zstl4CFz8yA49VQ+ICOPyIde1TUFX5oG15v1ZrmC3iN
7YsxxKAocTK9sNFI2LhRffEVPjnXu3ib+KhSgBKaPW16Ka6ZyxoHaCW2WHZ2+CI1
H4qOf892Bks2yfAAm5YTFnT89T5UiRkOt/xHdtXSOtHq/gYk/8/44R0OFfuyS7ws
zj1K/9y8HSmxgXhUzIZ1tT9OdY7ykGJ3JBrv+PEhe3DmmDopJPsFdN1kINj2ZJSt
2DfiBxIEIzFSZkXN0/LFATc8kIK5iIwYnJHPExV4hUCmp/LZzvdpzZCvW+Y1Nyc9
IYDEP6spipMWV/BQQOI4B1mC8pgp1Qxr8kU0zANdVmfNJn9uQTHGquwsvgZBdBFE
gKCYD0rG2ye2HQT1ydX6rtcjeGt0PYbX7HNptYGaurPJZO5CkvRYX1B/p8Usgl51
242Lor6ou9+KVN3A2i8ap2DQRwRVLSSUmW5KuGif8jsvRvxM625z2Ra3nwrhNwaa
gTR0U3Ij6fdrJhv5PwpX4Mwszwe2kNNyMIGL0RZ6gZh12wGaw7i8Ff792MiVgByu
Y6XIA02h610CBhZu27seuuTLnZqIssxAj4P/H0oFZZD6Vuu/HRG55e/Ewr1AzQYG
NwK9UF+dr1aRz/nHn7NwM7yaXm5QEkymJARFZXzw6iPg4H8ypypEzpdC0xbjy8tb
/nQCVpsiH0w88Z26Pwoyayj7afbt9kbB29mq6dTLN025ljEiTx0xAWP+EodBkiWz
HK7m0o77spW3HhU8RJhVlsStlP7yhFOFY07jkLcmT9VpkVvu1A7i/52ZRRE2+eUJ
Tcn36kJp+dPS4HR4oz7igYT1gqirCLeMeW7UenjALq14Wf+zgeiFKB78wR7mMhyR
U8NSIzzTAj1kHhS13bP9rmfd/aZsD9AMluOrSYm6He1eGGu/SXiJ8q+gVnRK1tP7
boEYk2lKO0U0XLhWl0JXzHEj8sGsrZtVWYDRst9chhz6v6LIW+hi/fTMGFwBTjDX
UIDz5h+RczZiUKLSgXVR7VCnIXAVtKEgc1JkcRju8WZzdiV7a3FFkd9MCrFAZ0Q2
6EKWg372K+AcBSHh47j5mCUMCqCMkI3xJxFtNrrLH+jiOxdBdQo7sohmLAknhGvv
WrPYhw8ZVFs0o/zCWFCrFu3ecUxqr6ahjLoAtr66GG3G/0EbtmAkl46j0SwLHJ/G
iZqw1mWop833UHbhREv4Ive/T5JP9ZBUmp23Dpf6SSacOZwxiTEbWiSEoEn0ZBH5
PYV0WUq2vxC7SoxlYe0/NllvAj9R23nUsoG68omO8UOKKTcxRUlKvpm7RQ1efox2
An9S54zCDKw67JE1MV3MYUIRZhW9zPrCpyKESSimTZJTPw+r4HM+fjBxNKxSYh4S
aaKc2xyGqgR3QDN9ECSfx29ZpYz2He8s6k9LULnoV8McLg1IuVpf//TTNVE8CRbF
EOKtZtvL2BL2oE1IaCc90heoAwP3rG0PnxZ6KNVRzYd7zYn3nmT81pfBsTNsBtur
5uFrdiE9YsPQ0u+GlukOjL9b0dVa09acvWPgqhNumR1AoyzLqgg3pgB3UnN3dzhW
krgd023Nkda5p8D9ocSzHw5egxeQ8b367k3cmRLT542HPEQ1rhy7BZXe2KY8Joaj
mpy0mbe2HuEXJDz/Gow3XLoG+yEj64btqL9lpjFHMlu6+iiwmpyJoP6cWEYbnteS
GBIqT+RA+d5UCNPdJCR+Y3KbZmVclQqTliqEJ3uxIMVXlys9SDTcWuLkr51lWkon
pKtnAeHEVeKnBS0b5ASn6tzzu8ASKql7yzUGw/gjaQw5yfM0ARHGc5zzG8GFbUsx
+eH3GLh5XXF+1s9XYGtkL4sTiASyKwcjYp46WNoyvroW3hl0OIkfeGddLnIkvjnn
g4ym475Bri0S/rNn0LD5ltCcZ+oL+5mRyBr7XKV7KyBQstC1mEmRpLXL3JZUBO53
uuodKv9Ir95qzo8SbTzf7o9SkyBW8yeLARCsKn/UPh81dKAPayrwdkh3yI0PNiMk
XejBe6sqTyD3oZdJ8uSl2wfxVIjhmU2Tn5Bq+Yl46/wK8H8mVtffhk0XHJMtoj1v
/ov4FvYx0u7s4JAp04GvcncgWXJXxcOB/v97wdvYOpmbCVXasafNDxM2O0kn5VMF
NYqqGNQ3x6hpjDr40bqOg6QgEIJEUzEtBuWIjh7Jbxu4sRIW4it0y6YYiKHSsuyi
Dkg234ncyfZKP70pp5/gCG7AfUD+yl1jqtR19wpOY8qp54jDkrv9LPV4d1H6lL5V
jJaNLoDN01N5QUJXy2xgSdEKK97SnqcVL+2kcxFwwCde8aeYO/arMMJphb1GzExc
8T6VisXwFDOqRTbeH3TWgvaBDP+IEQTSKzInswdhUa4x4PkR2XYXCqbsJ9BTuuC3
El7TABj/9Q3OCowcoorqy648nuTHpb/8XQ0T6R0XprG9fncg6rY+su0v5syEIIlp
xkmOy2nEk0uoH5ehXg9+wC61MYQ5ELYhpYHf+vIvNfcyqXxsXtnB03Vnlt0FRKXd
5umy0k4S/uUOSizhGBR+wp80H8se+Nci3J6qsRaw6ZMkC0DFpNrlLywZWQz6tJpi
WeLtGa/GLTyDjsohSdKhCCvEbV+U9SOXTlgYU8fMqdA7+yTcYpYKxPZxy4loKB1v
tos7eumFCrHoafYVuGeG8022PpcmbPhTThhaiVSammOtvzu8nEFuImwheW4cnySA
YuEpC+x/UmigHWdIeHK465r3Nq6UQJ/hwu9eVQ+YS8Xwqz5yXuj7rf0GeXrace8H
/wje3Z3qVissw8Oa24dcKzj+x1iCr9pz6SNvfXDo4aNaHQDyFvNGLv0np+Rob8YJ
L0qhWQOs2MMjbFlaGNAGgfs+aDympnCsRy1Fkktn5zAekJEszmXZxZCAiSWzgLU6
jy99gC8VnGbBUDOknLz3e816xcBV7Ifme9N2rzaPVbFRTRedGWD2d3t4/u2YFQVv
KUttf3cgsGC1V5JOm1rz2f9BMGZq6xAinlZp8Jp3c8nBpH7mj0fvkjOXAGqmjlLW
kJo3DrJl/I277KllnlSpbsEZNMu9zUrziw8lfkmqIQpwLfB8JdCtgWjqDRgLzrf/
jCJYiLhBUQrOYEqppz5BO86ZTsfoIxAbycCfcwICYz7DtAWSNi2OAJm/BvBmYXgg
IjDAFqezK74rlYUUAuAn8nZWxnojhDWqdMUEefv+dHza5up77K3gRFAwENMsliJ2
00KQGzeEImBbtZy+gtISgSduPCmeIBbGhIrdSeNu6WzJz9T3FbxTAHxqRsSE5lX5
ERk4CtH4yzbyT3k09Fy6MT3/014Ob1nUnpneyFy54d7L5b1yitrXtWKpOIlukUOP
Sr53X7lfeR50vSm1v0/2mvsm/GYMj+MWgu6Lg2lyvlhimFIszpz+k1ykjpYn0iK2
CM2K+aibS43U7OaLAwvuPBPWoZ0SkoH/YqE5tmwa/EL20sFEmEtAowEoVRf7B9ms
j7qZQS73daieku/71XORtBnRKrPnPvKPCc7i/xcrem+WRxgA2Rb7ocHH231Jn/IN
SZa1H09G5mTykMr6H33xV6Ry1wFdgjZ7e6W2B1ZIi1kHhw612tIbGWf2Xb7hDKkt
Fh+XVVumHAgcHxPxHtVcc/QDcA78IY4emq3zDDKzXrLeQ9+ZYbLV9CK9GHsZTmIf
Knppnpxv8Ju5urrNacp4ofBINGX3lFYRsNGzWsgGZ7oHyx+LbVM8wflM8GdA+ucn
NuP01042sRYEUIDfe0KOvvpMaACocFg5Qub0i+tOjU1OyHgtsCJUDd720mV1fma+
36qKCO0VH6iI+zU3yfYZ0uFXri6iFAGinJPPAsXceT3fqnBiOgPeM5CuSU963g4y
sMm7sZ241u/PplayvOTwUp7UOCu7um2te4ZNK9hbWe+2rU52R/XC3IdY4bN2jdMv
UPvQ/g3VSV7mAWa8ZP/VBGTsb9YqOo4rbXsreBcy8ooI9wZr4iaOdiMhLYUR0NIK
aB/f7JrjlOti4ued9awsqIjNUhhQGg4Wq0rHdyN27FLmEg5CjtYHxlJiwsPA2Yk/
UKFPGaT249F1lDs2iD6mR0L8SeKDkJ2jPEo3Z/IvOi7tx9oSl6ySIFeSKy9x7Lds
A2VKDuRS8W+ClfF1qf5S7yGHNSsBHQPtIBpVf9NmM4RXi+IRkzQuyTDhIYfcgM7u
da4C5EUwedgwio5xCt7HSnj0BFc/RpQufaimKBXXbroIdJYhNapzg7/Cy4gKWfBZ
8pzgRHgsdpxP6ucLIsjTotHzdCReM7ZaNWIMBhG8XM6HhY9NuKFJzNfPUZoiWhxW
rEPIaGa+OV+eFLo9vOkTstiryrydrVwVpix6lFN/MHE37INUHGlwoPtHNa9WRCwC
cGq//+8iLB6vDS+CoKVNwmgHPmeSYnpMdfAsojWUXBQBGzkolhaucxIfdbz5saSV
ZAtwr0iEz/rMJHPr3WmxKiihiFgYIzKWLrtGVzbvJOA9aT9d+F3iqlLRD4FPOIDi
mOkIpqWiLwS8+rHq4bviPMmC1DKQ7cm00zAeREFsOfL6ns0DHIEy0ea0RqvBF0J/
kR9p+n+X70XPknLf1aL3H/g9oEj0VDRjww4gZaKHTOhdzmGLFzqPWJm2V6HytZ0g
YMyGAUfu325WA2eyh1RgDYAXAY5USVSVaEaE6AAsLSE3GeD2QU0OqFZ7tchBEPrC
ewlgRjA3pu0IRMuL9PQISQJkKYEzwYzGtobgMAApgIFYEfN+w/n0cXuHS27ipxJ9
p3sqaRm6kt37LTFe6Rz9Efcr7u1hdteEM2gyTjMaUdOXZ9D3daO1/fm1QaSS+Li7
tua5vRS48fcHizL5MCnaLR1VY+Qyqi1kpTEoJ7qA+wdaopwpThE0aP0aL7A/w0Il
r8HtgWpehBdFlev7GR2ge5cwux1g5AHzlyEw31LvNNCfWgzD8704CxpkFlQd8iGn
KX8mpMwTaIP8TRjLkMcWcHt2WuWlzJyq83DnV1sH82QCPLAzetAM76O2nmote4RR
JPkurX3CTynzLKU1yzcWeqMKogvGKC1X54J1LtrHbatY4SSSv9zMEPqevM78LkaR
vePLVfPOidKfL+Gyvg7GeuyZKK6CF4SPJP/WQJOrVFD08zc93K+1/LBBaX5DjVYi
b58p58JIT9gy01jl8lM0O0pRxksmL6720KAzCnyAYhZ79UkgbiM4wEFA5xygUHoz
75lz+5uqsetoLiAE/qHLWjAirlQMhLqVG1bhLXrUf375wz2RNp7oaJUzTKVugSZi
5fkPlM9x3r3xwE4kDn8bIsqXteeReOPRCuPK2xcKmVvuNvlrmHUEnwBndEbDyadj
W7UaM2Gr8no5RI2SmyBCm7pyzDti9otghG64P8DctmTt4F2dhqZizTppJw+PfCNp
BzxYD6ai0pj9pppbEUEi0vsy3pmYg4yZ4lZH0ATv1MxDYirtjj1oGs/QhQ8gwzMM
1ePwkL8Xd6TavIKLevuCF1mcJH13OpaN7wZxjuwger99HRmIaXJTOftWm4V90H6x
BRtwlDU44jbEMwRMLE4caZkk9YQ8LR0qbRHFsHDqiyo+dd6m7EJrRWaBxv6SQbNZ
u7ZDwPZ8JX4awbgxd/95sOHSnLKkG1nCRSPQwVDUfGLARpT53qVihVWCQiW5+bN/
66nP6qtrFCSgCmveXFqr9pamSSoTuaIYgjH0yAQ51PZGVqyjtrrU+n7VWFjpJjZy
tk8T05/2Lm/lzvKzp9lDwbOFU90HIVWijzAkIaKdPwN9wr/vqcyI2vmyIhk/0bNo
1XH8KBk7aa6+7YtuY6mzax8vsMIeRNK1tsRuqN/fe1Rm5bJyywNIyiWpAFR08663
AC5vYR1zZ3tL/eqZtTELavO5cjj/ImkQw5WZDc88VlDmvbcHjPAYd1b3Tv4c+SHv
xdA1y/vt41k3nA3q1v7EIx1hUECSiwPMUVGJ6bafo3ooBjvXg1NU9IHgneq5H/ua
NZBAGae7TVBMqA7Ar/aDNdD3dX47Pvf/zFYe+gu8W7dgkTk/ZDQCpSkg5OWUiecb
xhb9DwxKsfpo65QoyGshtzWDojqXRRn+pc39q3u1D9GTZI8eC4mA2gh0Uw1PTK1Z
itrGEiAeNqjgWvuOUL+xXj8PiE8XqTdJj8ZWoIoPA1JObtMfB4w2V+MecEdToZ8N
tgY+zbPDjtj1AjBVQI7ZixSP+HkNnSkMzKAP+B1PTk6ZHFvz4NfQLnujMLBK1u1F
M839UwblaeZ1/ODvP7zWYsnuRUEesY6O0yPJTbj71DIHThqOd+3Jj1m2MxBny+pF
tGt8eBzCemlP5Jkk/w6czDv52IB5MQWM95YMxcovUtvOagAVdwiLN9x11eRv8TGf
vQWDEvmDXnxZuGUQYzzh3B5CsPMWzACGLWI9Q29npXhEXtsuJtQfQAtnAEcV0Tdu
ewN+ZxSZu7RSyckZkhurA4nN+kR5nxYoIK/UtrkvZpXmfSAMMm/r2YwRhF6ezlyM
Lki4PHubxxa9nvfQTxx4CcnxV597b/x7z1Me/7sUAcCOx3UToU7JMYZ4lSh4Hdy7
BmvNPchJc36YZdBKvMygPTVsSrbAgQT5eOQhwXh8/Ptz2uG/2sy0B5nytNJDnSZt
tX0fBb0TEc/HbjTM5gaP1qL/FS5Km9cKE8M3VF7oLD+KeKawRwHBK+ghLi0LkXG0
MdjqAklA70INLfzrRmCgRRZ1pewhfF21K/k4we7cwVlCLBb5G8jQm76JlbPSM4b5
kd2UIwp+l5M7eTbT2FJHPCtbvP/9SUl3+e+LYHMljhW4/zBqPCoXp1CrbYd/D2oX
P1MwE2igVndxFq4KYAHMY5WIKucRhcthtYnAsBX52Q7tQKxEjNSiDCixcVcjI6GF
dttJ8s5+gvUs+5ggX6aYF7iPhuymzKzW0ZbGNoHWJ8jdl4cmx3cpiggiT8GAYyPT
lXvUQSTB3Io0U/aoBC3bXd26kPR+OUWNfxABO1geG4NXC48wuFzaRIIw7UzbX+T7
G4jP3tpm6USebmhE8+SREr3XAlysupRxQ0Nuxwjucq3QXYFsthrEKTa+R6gU9+Im
7wiQzx4EDJJMTjTrdkcLNyvUahRMGWESPaU0NDdFsodtY/AVycgTd97bV7guwaNl
BGOwmVLyljLeofwTH97vLdPUpGxvD9GUL+ytCc50NgVS+SqJi02rtjTWIvCYm2jQ
/qRwoqdHlkCMhzmF3my6uX9aiHtte+BtoxuYatsGVYXMo5w8JqqYt/MZdRsUtwqd
6plaXMPdckKenZLXnEqCgdrpjvaw5n33usem5oExCw1eTIHdN/fWGaWocQ3eSzMF
ZAu6HcgNdRHt0sJDyt30PQ191PymPSUd/nWEvU6hyw9wvI8CzEC8YQR+iR17Zetx
DF/UZofjwbR9c8tEOnZKKDDHXqYqA60caYTp2KxQsB/BnttgwGnGUsNvswwcJl2k
zTRZCmHdcqNyPQIqR6Q4knHT7W9Y8XQqcwPKCozpkHlKmTV8CdJprfMxjKQG1Xwd
AgnVvf2OE9QpnHppVYViqmaqlEhC9IKxjz92gb1obqu5DtrktXS1MhN+pioLA07d
pB1y9MvIZD4eqgZqcqq+jroIO/51rHfLyHPFMD7hjG6spVYmXjQ61r8V3dl1WR99
y5eXGD+vhay1rrNF0uFLp3MbfM/xZncse2ns6oqqtC9QgG4JFWniHa129J1k28fL
zRx0B75FuGvO4owvulz4NX2t86KAPxPjTUxjDlhCRTUzdVEzh0VNieyDHwRKS495
alMj+RYAPtLy2E2VettBZSSbAQhI3Vz6lrDZjpqWS4DfDrKvn8ffj+RG2pX3fiGR
Twz70U56EoX2SKqw4TzEqKXGAhhEukhXtCwjf5q0E5x5inrLrmTRQx3XYF9pJ3e0
4lezvJgDG9zfuF3ZBMdRRtbwMA+cwfSar5eLh90pijIFujI3qL5cv0P1SR8f9mO6
H9CNSCBsFG6TfxcE7ahF9/XZKm0g8C9Us8OBSSqYckmPkQEzM/TM+ZeE2F6oPk+J
fyhEBYyl2b2HBOZdFqXQGauxD2QHAtr3ZaQMyS284sVkKe0uwnjQHAnwQOyO0bYy
Y3QSsVD9eB6UGtu011qdYNmpR0HOxXjzRBPZMntT0ZgToL6VivRaedXAtcmhVMym
RFZn5VBA+RhJkHtQCt/0aBJcBonylnsFS9Az6Ikhy30++4v9xZimXnOwjMpxFbiX
j5eEetmCdPoBlafEr30oZw/qkTI9QvtUjvllyhyiaskk7HkVROE3XMq7pq8yLdub
g2l82m9NBu2ZqwShTgWa1vKDVYJ0/yDlIH9e2FwKhilxMFW9XuNV3SPzoIS2zCs1
Fgr4F6vYWVq0MEfnDhnojzTOB/QC6LpLhcsoby5h8IpJVnyWMKcZQgYYg0h8xAWq
AxZ0OlFlj9W1AwFNYzNiGxa9hX5o9/FvJm8VtrJBoFko19F0qzQpQcBBpWUQpUEw
MVorLeIw96O4Mw1dpyv0EdJLBw9X1lKWD+ke6khfvn27FCm5uDAZl8FRnnbgtxUV
7Bu21KWaW9qfzsrKSxIczK3T2Y7Wyp6LIgG20qSpgHEp19MGSWHFlri+c4twXbca
OWTWd7Op1RLl5y6JBqT38iIhL2iM7703vJKvJ2EfBypCCXKHq7TE8H2gTnMfyt/c
fwLO1jXNJNGDaRKuxpLW6hPJtn5CtLQaq//ZskGuCtVspHTRT0n4gqa6KtvucBlZ
1mKeSjZ54gyUoD9VXmer1ThEdKGVhL22JmyGUnxHdWrtRr2UmN/K6nW4apzVoL6t
1+wrqlVKFZ2+bUPVv6yOlcEZdHVDt07TTNf59tSHE5i6I0TkUIdoDe4/sQu26FUD
L/GxauZG49Yi3fqwKNm+0z3m0HqNuqbe+v2qOogh5IIwp9YNAb4y0O1ed0BO5X5k
q8oiLGlzFc5YTKrApFtYx1uWBkqyPpg7yjfRJT1SfmpGxTD39twGrIoHDe46iPzM
566bTPN4Gbvtq8s+VqE6jPIJZJY3KDlwG1aQks4XrRiTCaDMv91b+3Qohc+1cAG7
VkJbCHAL4JxUgvKHQLbAe09DKMrZpX/fEq9z08KM2e0WYjFJe2hNcDpZivcad9em
DxzoT1fewnc413LSbJELEZQu0tUvrIXFvwWdRwJHL0384GMuXGPxYfy6y9X6wEVA
j5iPknz+4EJLx49FYaqZaV74zfZvpIMgA8FG//A/iJEs+TAFB+n5ul7/2wKCqiqi
kX2pnDkRyVL+aTjiMonhiV2QbYByShw2IOZIpuFwFVQc5bkvJtB1Y1sQxAIgmgWd
NoBqxkdyfF7NmUXdxlc7ZZzO8QXgrNatR7ssPy1qq1A6ODML1i6fE0TRKhC1mNxw
WDnU3bvIbIvY4SDC3sVwb2HbspJdsgnwV5i1vUEUv62gOIiNlWJMxh89uTWQ8Ag+
8pCHbWmnucm4YhZpff4TX4J6vCDX5ZXXdDNZN/TH2VjbPGV7GnI+kKotLj6BNZma
goTQOCTi1jcl8a4tHuaznzvtK77KLguFCjsAGO/fy21VhfFd0yZBmAt4idFhXY+8
NA+J7+xXHcvNf9GRnFUdkAHN5nZMeY90aibt/YOArFCnHWc8q5f8DjRQhuTRLnGx
l38NDNCl+DIY4Tl85i02duF3rTcvSCRzIJF0B2vjJijawd/iGuFvjBVAKSNZ36hL
pE6yp4DhAKtWyZ5NmeBnsaVPE0sqKEXiAeqoAkkjtPTtGKUxi9wXuSytmdpDol3s
07nQ8JAsble0P+o2V1uRDIbDcEy3uWXUqbd8nYT4KgcyelWS1hdxoMyzysqbPoGj
M1BGrrKwIqeszii2znPdZSaYJ95BqYRt/rXo5lrswpnQ/yapHKzmqox1vCTGT/bj
fC2TA4zOcCi32x2sq+JKggyCdpe3GXm5mH7T2PrEEwjOTLCYuP5GxoP0Sq0LKu3m
Ss77FOATLJEQv5eddG66NHpq1vIwTR5kBaOZ8wfibuAJnXmkO1KFXwdQ0sNw3WmL
Xp/v2s7OOmD+BTedfHiethuv5xYPm0vi8b96A1cCoMYvtgupiikFswzjDcz/Crbw
PNPuVoa9wPGApftaup9GFVncnDJgCAw9HZPzoNURxedGCDYVp+qhN3n9fU1mSgZR
sW3ViygnZdxBbtV9lLHrChUTHmJpmqlYzN1s7imES5YFqN71D2HevjH5g4ZFSTWo
alwt9lmZp4CVUjwK7YqwhMfRUeekeRl76BfbEASJ0Ed6TaVuqEqXwiQ1d5temJ2z
NOJF18JamadvrYf8PRIAXSqejJEEO+vsarHbWCu1aq8Dsi74N2HDymYkY6CnDHhZ
KAmDmrJ6EKKkxmPkUJZGqmEJIqnf/bFrqiQXR4Rump+497PAgdlTF63zrYjaBwQj
PXSqqughJqaQBF94w1lI0J0UO4wN//KLK+EUSDXLr+pKKHdqUFpNyLPoRyHT5l74
fBx4E2jS34cNYn9BxI0v23afgoEfUXFnhYGSUzC59WpWd0Ug/KJRbwhwqnSvKysv
VNH1DAc18yjKdXdURXCmWvFKMjNV3miFYKEPbimfZPKgXh27b7s69S+ylN1Ds9qc
k+Sfu0F8P/NTaKoNtgwUPwEBvhKzXC0R/2ROaJJO6hq5pDbbLHTvsvoS6Yoabf+K
SdBY3zll1fc15K0npY0hqiySVuRp52SJSwOmvW+J4BMqvVDhLVWYmvkXQzbJVF4b
KPGVcWSOCcAApB93MKdxkfqalCk2ZjHMPY7nUIuprcbiEkw8D+wpRWog9wUAInBi
N+5H1I6fdO3FMajJKAQgQ1/0jGzvUTvgEmcnJRXj+qxG0sNMXLRbo/8YBxsWZuGA
/+jyqi+G7ZtXxcVOFTAMqq2+a+GeeGkAOqIJIl+YUNPSGnQ+LbAVo7ab5bUQo6cr
XqOcnWVkOVDvDz7l+oxAd/oS1xY4E1++TPuMbOnn2e5t66Ht6OsXjAkQ+Rk3MDDa
5OZJuuJHz0ibhb1JlnTGM4i+I34op+MK4a2qdgyXDyv0Sc9YJ743zFZu72+eHok0
q7luRQU0YGNazJSSaC1EyP7EClyC6BXdQM8QRDb4itpqNl+neP3pkunk362zsLEr
zK8Wk71AaoJ9IcPbKQaCXaVbY24zGLN/B9F6/GuD09fNNdctChNZvltbEPmSD/Js
x7K9OpctyDCq8TdZh4V6PVci2t9asBkGU+T/QUa+rW8ynaFP9nqe+IkaanskOlcS
G3Odr9mBrEWvuNjmvfx8tfgIJO0OsL6fwteIeLJCawNmM7Ky5bzcVRK2/KY0S2na
TzP6kr0Rr9AykQG712XtpNrXzionD743f61BsKRL7ckuVkQVBEAydXlK7A0ECNq6
0rqV3k4v6niFlEbtkuoXVxGgFl9UoLd8nI6oReoyWzZqUDnTKAETBS8fCrBVqLAS
YIBNmrDzZBq8/TJzEC4uQl/msOz5HHIweUkbSZnn7+a5rH4BbIZay/JrwpoYqBNr
/lrgm9m5qiadr2HAYPp4MJjk1Zdxq1lc1VUI3vdEZQrIsmv6of1sC8UOjywh5SOW
/9dWe5zY1WJ64NN0p4psfpICVMQQuoNdvBe9OBRVdexF9Xi2HVlfhhXHOhbF7Iks
yUdYisKcew1b3IufWgcFgHUeEgP2g1w/+5iBN18ZT0UQ7B2sNnxFlgbBeS1Flj6U
DPzMrhFs2u+FCMmiBMpksxi72giXIoc9do830Iyje60zahK4dtBRT7IuIGBtfOv+
pOgyneJDEgYteP3gAYV4hnm+tDPB2n8+WGm9pDWR7Q0vTotaRjO5CetLfpcqvnVo
wyFV7UWpZiqhItJQQ73gjXUCgz2gGK/D0bAoEI3n1zY1ZnMc/mm5HXcfUVqiySgc
oc4NgAXx5qAU4AAFhQpTG33LzHZlqZ/fXQQgQi8kxwsfoFSlLoWTBVFn7HzkvwKo
ln9V0oKyN0PARX1A47WrLrLs1adOtD5gZGnhE2GiaOy08EhSnk85hQJajWFFK6Dx
BqwDl22gV5S5dQJrBvl/sZREzqmGQITSM3hOefAwxESUWWJpTYw1v6O3H4JfQO9q
xQRq7zTnDul2e5ednkgWfEja5TOJt5O6xdZFtYHLnUvN6s2Zw2IlASTPhCyYwKr/
Mwkg0PKm4dR9cU34GZFak2HLLKhfrd/hX55OCS9HOKj3KeR7c5zBHltGCTjfTDzk
uBMFY01q5AwPGoQ+Dfp6w1HXAhtL6ppHrrfjVHZklL0MMCGJYfBUhilkCGJHAcRl
vnB06wRqsCL045FT5xWT+p/yMBU5qZ4XP+Qdd8uLGmhOiBTx4EHpvekQLVVq5IS1
DZ7H8cbPDVr/OERUIK+MPGCvoDv91In7euboeeezTF3mjyIQmZaQIj2tfjzn1cib
4w9IynEvZXZoAKKtpfXyfAa0u0MUttVPjytlllzkhh9tzvHUoJmHGF0OBySxS9MV
HdCKoT/FuEyu4NLFPOwrymi2Ur9jw2aa0JpLDtSWqOw7LOD1r9iI8c5sORFR+30A
ZJWQ2p8YWJeivFrEs6ZzOIvBXL15hORciAozduuRxxWK6fvB66EL7yE07CKbrhxB
YKLPErXELvjLT8s/+8XpFdlDTh5pwV+xeolIW3WxxwdqzOwhqNFGP+JrIQYAMSHL
7+GemYBb7VlPpm2nPjarURX54I0BVkvp7oCwJUgZ03bOqV1q9GpiyRwWAzcCkWpa
pxUpzh7KeEsCJdwEqY/u3t5udH1qPWHbpRYdsnyWR44UhNirlGyRctP6rsnr9Zq/
8MYr79Ux8yB4fG1VlUJ7E5zOjVv7Z/LoCK4sb9Yk1eClEETO082CxrTbrmKjIWm5
wycuL8tlU47uJwDyOlK0NtN/3avBgww5EJDqsiNiiMFSPSQLUT+kqndA+wiy//Uv
fo8AmH0kax5Jyg9EtPEMO5Dgd7ilVHRi7G8Vz/h0/Y7qKgow/jgdKeIpfcT7fTZo
GHTdl2XSwsm6g2Ht5s5B5bIqDq2z3O3KyLb1GoOaTLmk+4inr0n3UzbyhqtnlrrQ
Ae+2zYR/t1vWmNZrNW8mjIfZeZhuNax/8/jJwoAIUKTcoQzrZ4eaC6w9oINwksPg
KYrVTcA62LPlW6prPdBfmvEgJZMYkxxyBNafJUvu2ckcN0R1A9Pzvl4C1AykI5+z
vRXGoTZZEngdsWL/3QsD/6hTEiRrx8hG/sdxmaZ+sKSF+Tj/bOXRMLxi6X/SJZTT
x9dzgAEDe3UT4NHN+EuT7ziMHh2yTIBfRAGxWL6cAkfSfAXJhO3l21i5iledRSJs
HFCEq+GQOzpSQC7Z7hth3BAHf6dopewk7tWMKfBfj3jVIQAmPDdyqm3UrtB/rYJy
epSR7wgZpxt3MvQ2XIqqU4PqwZMqqnBhWGkOtEOCNoQwLPcxsC7yScttSK+3PEhu
yO+A5XFNm3ihvo6CNDKuXWSNQYYPPM8xYWB3hqTOMLDTCU5B/whB09gmgHhohFEG
2uEOYS69KviGgRmWTg8RJkrqdF/CaD9kO8O1jrsySRo+o1c4JjLOv0JiTzWCCHnZ
D/BNQiIAckf94991c4uLyW8IicThOmV/C8/aDTm4QBVB5+JPUnue8J1fO0ais4zP
XlCRJTxuj6hK2rK27es2FZs49zCt42pBTpFRxQdxKmqVcIN2YzDVArSuA5I2Nbl2
MGICua0RsF00jxa1L25nMI0MLAM3kiXcFrsZpeNM2S3f7KX75SlN0BadhBmkN7Gb
vec9aeLNRZjpkdna4mcQuE7dHL4mRo0RSVqUKsOsiTkhZ73CqzkDbO+nNFmTir/y
q1TBb+39rVl9lXesHCkF8IK45tmEKKozd8KD/hvhlKdL9nMGJwD5ZzXo6mIfa61D
xSU5EFgkXwELdZkkLBRefAkdXcWWA/ExsUqFQzF57kruWt2v/0y/IAYxTD9JTech
vIGbSwr2j95Ih6V/WdhIi1RvkHd9zuLS56teyijB3JNxBNLxpj/qQQ3fdduP3/5v
S5rASzCfhT+iHOGrNYniaV0kIWIbp4VTOU/lvpVzdc7K28vItxAf8BThdp8cR3yZ
f/Evfbwrn/wKdX5zolxm/Uv1yQoFmKmha4c+CaFK7WrZfWpJg2m+lvJe9nAaQe2A
3VVcP50Wkn64UOMMmzex0Ty/oRV7VefMEYyBB7Ree87ubY4e4KxCGKDXotFOKHeV
hCgJOlbcTnsMyZ/168pOhSSI1BrpDq5jotvIy96dje9QJRo1bDgqXaDQCogGOuPe
DCN1MN54XFTjUV0eoRJ+XLzAhP6FFVOQeFwdwAL6znKrnvsXTF0n2BzqVnEI8PMK
CVzAMEGFFDiAo6GWEskHBRYhu//SXc2KupT6mMEo52n0fAaEKmPb7+NpVX0MSA+P
Ct1pZS3Ipei0I20+ryQFf/ihNaGZDYX9+8rQo0A2Rf4CLT68KWlyfUuDqm0MsC9Q
TsIREvHooU0PQgMOCWXIcR51ONvw2fouXH0caCL2MkkjydyldlJMFCh3J0kcQtLy
BQKRJKpUyJ+LVrB/zpdzc9amY4RKQbRXPg1Y4vomCDx90UcMgzP5ODAO/JQQAcqq
lUTF1t6iOqaIHLNSnY/WsiwD559/9DiQJALUO8LM8aUIEXzrFBvjdyD97M8uOdYq
nCqmJgoGD9d0jFR94lIUjJTE2xZj/D3Gz8h5cuz1MPl8MGqTEp6imx9PIUInco1v
+7SFTBuND2YD3kCyO+ayWUZ7yF1usXBIRoAECbwYBDqBwl27/+1j0fIwxsPoxdFb
go7OaXJuSX22K26jezP5fYPX3U2g+kgb1bCX5chBPKNjabnuAnju6M+tnlURw16W
y+d0aNe/bnEpoGUJdKVXitOgl6tlh+S3HeFEY7nH0U0mHFzXy3b39Y25U/8ZV6ZV
ZEz80aqVGf7kb/dCCKFa9dgMnGSted3DL8e2dx8+G4Nq3V+/VO8Z2OBw8TnlAW16
O79zf0EHttiB/qfMjgcGq+7IS8b2bUKro/13DfGBzfnzLN36DKJ03SGBQANn1reD
CXu+vBrIJWTJVNGoJ9rzPHZPz+8G+8GV/VyCFNBgj2ldzdRC4OujyFgGrdvHduKV
5oEOnYkld+2U14PIyS8gxQ0k+L9VkDZi1+6KviuWPgm9JcJ154oiC+V7y+GRvMEg
KN5RF+e4jNinGmJCRax9vPYloSiqcaVcZhpb4OLwRaehhnPdNFP6PmwjuW0TBXUV
BWhU79J0dpTsEA/m6mJFJ+11UuGk1VBqe+JGvmXQes2F0nFtCmrdOkoavP/tY0BE
g4W9UG5FJkbljeFmW8H+gBP10RQxNRPCbLAPtgSkikAHupuMIewINvF/MhmoaUcN
EjiEQZb/0GUcztzHmAgHB+M+3D5Rh+1Aq1y8PURRfQMQ4uBlHROZLUEJdqsqdoeW
Al9aj11efhaWnidHdMaeT8YkKrm16i4408DTVcGA8I3E3Bnx6suzN5q0xfN5qvw7
4sS691OvmiB44rZz4FO43YEcR7EB77Y9n+oGxdDyzg77RC/0t6bkNB32ZhmpRhDl
bhWT9ZL117ZkjTEhcQI5rvDwavM/VE7MfJ1hbvjcYyoXxDwR0lGtPFIn2UPC4pcT
tjPNdQ5ImKX7lqi3L9RaNPqR7nrGOEWcI0WhczUXIIp7SRp4cihy3TsUqEYhKtit
j52ZPZbnY3gEMB80FctcEq7vyQrkH2TxtnnuiwqhOWOkxKSRA64mdNQR7n34fnRn
CQS7QvB2rEWK97NVdeTLt5zBAS73xSSXBYalvgA2BrqJo40e8VLzYo2Xb4wT29LN
uanVGf6W5oxGmMeQJNKg51oXW7HcHZDJDxkJYF1zTCF0UwU7SBy9ghfhAsFrPA0H
7b9hDZAYJ7anxW4RyUL9wcRkuRaGe/nKnY8OORWQeqG6SaYbcP+swuEJTbFQHJiU
E++d1tMnIzuUj7KboRvXBvhwcofFCLA5RRdyOWDR1zbyadwsDhQb7A1OVfDM8+Nh
CXpgYpD1L3uyxQYWt4jPtuIFJV6kbm1jr178W2gmkSdNe9K13pgvGvfFYYhAjauv
4l4BB4lGT3sm3Ub3Ph+gBWWiYa8QXNmhYecLzhV4F2MduXjlQB9K1ImjfsT/zvKd
GK4/7wQAmZVasM8aidOs6KdIpftH+YJ266Gw2ICENCsVtWDHdnU57RjT6fW02EHr
NDYgfRfkUxRX2btZ1PFXjp3omb/vgHESmZQ75q//Sk+pA4liDFJsvhqIaS15aJ3J
yp40pSDubWM3UE3GQ+xzxpr+7E3v63QwhvLQXJ1WxYSOQWj3n8R4Ql7OTvDi46hm
rH0tvAD2aibcNf1R9zPcvX/Gb9CtQeJ+X7aBPFhPPncFO69XcAk7cI0VXbpcWXRv
idHXtvbwRnTayfkaiuRLDTfp/MeOizubtD7Yxt3i1RksVefy1f4SFX/LfYZC9NnX
VvpxdNf33fm0IOoJYhHUbegzvtXbyqfgx35L5d/NYPsFfkPeBuN6qi/TvYFkxqbt
rcawijSyd/cIj/7Dn9SF2IFZyLK7noAr4oaQUyabv5TzPfVkY4t0qmjlKbV5igvY
T/qfa29HzwGTV1drd2b71XIFi+J0pQoAvwGDJWhQ1y+JcMKd3S3+E1F+ZEq2rqKz
s5Mbn5cn1sWWmvuXVVPJxdrtbfIBD1pP7SA06LZWad17tzYWA64Umo4DsoFkL5O7
Wvmtetvo95uLEkOY7fmLD5UzA6qeMTMdX2LQ47FdDqmrY374+8Q8Qa4xpzFqMH2v
E2MVCFuly4QK+iy+S9BvD/lGBCusj8bWTysbKjXT8UE2iGfSCr1RvNNZ2OWdzA61
GBFxPQ7ukfkCSPJXR7DiJiyan0DJHkFBW004fWTCpou2osN6v5J0PqLOGFvzNB7t
f8dEJjQNmJCyKYb78SvUMb0w2mD+OGPvtVH7paGoZstoo1PTrc2rRXR68D8+CJ7u
OQkolYZxz3h3tMiYBBPYxIPPAsnE6GXW0NmS0dLaoZOwJi1RL+DIx/dihbMsAO1f
3yQ5CDjgwBtm5akIz0Egu3y8T+Lqt6ixc7rBJgVT2yFfcBAafGUKugkcZ7fdL4HK
6esvNxWG2AAp0JNfus+4JCu1a6Q8YnmtJCtyr+aPhwoBsEx7FwSitq3fvM4D5TF2
Ib0DVC3sHwT1u0t+74xsXctr4jewApcIy/cHNBTy4lQqmXMCVUI7tKAIJE0BFbZc
LfzCG1zHqEzCBk+OPs3PUo4uKAJCf8XBeVUuxEA9fH23Av0NabDT3oNftSdE1jM6
zEhQNQ1BrS9xMDEqjVNvMxfh9D0gySfdp5Z1EIiPZ9bc6sapfMqrlz8u8L/NO7ak
pH0Iu+kmHfH5OdaBJFG3Xg6t35bCwSSbDlGKhPDcKfkfG9pORjgJyyPpIgmOomhU
KrrZQpuPEf4rzyRDJ0fD/QuXgEyuHWUDmQa4kpbMacOjxCEjj/JBP4bf9LbGWwCT
TGW79lNaxLIyxZPC5tbWA563WXy64fOz98hNUGX+QUA8Q6ne3g5prAXllPcTXSxt
pCECwug0kI6Dw9S/b1B3v0RX5VWJEYQA4Mo8Ux4CIsKKk8pTXZz3MkJr/yGTB7+Q
LmWSI6i1b+20mm3TSSQB7yihFx2hIclZZRS7g3mTa8+kLuIi6MY+w/LoZW80zwY+
5o3+Gf2EQ/TYaTauyAVOhS58BEpIqXnjHnZHRLBaQ/Vg7c9g3db/viJeseKV5CVO
T4QrAq4ED7HGFqUDx76sqymsBUTgqFMG/PcIvtviO6D3kSE8ZywVrmbjzSYpQZct
P1JPFdz/I3kx84tjMXUGhaYWZRjlBbUquSmLF8MOKrpnh5n6JV4oqU+A1Oa/e3z+
oSIVK4ItZ+iJsHGTWQ4kMGQfVoIX3Y1mZVV7h5CX6NizrZZ7I1nwOSDSK1wkpkkL
WlDZCKlSjxIJ1BO1Z5n/0MW1wiqI05BKQTd4XzLYJhZWTBjcQDAzvRgY8Ta5/iJJ
azhPltkyHeCGxdChRVHv8ju9Ra5hctEP+va/enyTYjEdIvnRpR/zaJW5Q5f47cEw
XZZAU3tokJqngQ9LWN4rLgx1Q/Enaivb1n1QeqhBuMUl0DiJYDhUH7jUp9QaovYz
KtY9OPgQvfyrV0ny4fJVFxueLxauHmHFL38H3W+2jiUE3P01GY4ILbc3ByLikunb
yN/IDUgagbp+EP+vjv0ZFfwF6kG9bzz7KxyW2HYxPBj8JKu+wfCnjHOyfE+Qszh4
iEA2fneKMS7sS941vpStylUDK1WI39tVBEQt6rRyu3MQH1I2XSJVensicZog/t+R
nWkde1j9yhffrTtYjAoUzzB8zFgmbeltuVHC8f0LgB7S2zJkOQfK/optQYvoKTTz
pqNLgXmGR/46VkmSj+d33m/yR5+QGkTENPcpTu13KZ6GuiiBUQo4TwTeoRmCyGqw
Anu0DGDzTfFi+q3/yAjKc3FsHmRBRvIsNlpeosyisOw1FQEJ7Nk9VyEL97k86wev
L8VO0yoKwdHGGmNS4OmylGl7PTmMlllp8kvAX1/hgtPGowjrNXWeWrWmGWW6U/O+
d5GDWnKdtr1lMYYe9cT/FlOHeSrwvSbccXEp8e8yc07o1XIJAnEempWeQHjNPXM4
jztovHiry43pbIICCr+LVm3sr7qggJm0dutGb3jNizhfKFqTCsyIG3wUI/q+sHlW
c5FLmFm5BLnqQ6g2/GI1EdwIJQSiVUHT4XPTl7zgrU6ufGX5iXhmK4a/WflLHQXq
iBvfEleMFuQnbrVLEyytN0whAiXCHLnt+RQLZNQQJ2TxWFy1iWbziqo90xTnI0Mh
KV6QuqUiseub+RK3a3mlsNHID+PJToeE85ICUGd5LZz99Bo9eh6CVWbbLVqHpgDu
s97FZaGRxU6h3o7GkQqV6v1psbmbQt/l0YN3xqPShQU/6apfMe/MhkfnwXMgwSMr
KC9kAnB9V+kREXTrX2EzjGDSExdavRBG4v5MB6ldSnOQZfBZKh/sM06dRbXFFFwz
mvbywFsm1geXgq0oVz+1EmLcJoifsl4EL4NEkb0EgyETCgoX/dhdf4HYew7ktkMS
h1CK6xVTxyMlNL/MDEXB1m0ZUHq+0qWZ6Xl7fMoGrPQ56xYxZGsRUmniJrwuiR5+
wB0jfVMx3NEt4O8KmJZjbGNWbetw4qWpTACpcBtAXIWYwVzqLy+VkSPbNcbMg9vg
Y3YhO0lRovWBYdcgkgYmPW3YxoJ3782/VoAtsOM9IHloILccWI0y99HJACD5pJ7V
8RHR4ONQ/BITR1w+QcwviEFPbzJQOafwrPU1BAlSansF997goBnHAvtmqg2TdQzT
kE63rZIFA85qES/XYfPTyXoYXfgJ9+oay96rXIq4ceObLkEoelapokVVOd6tKJyn
hMcSpAx79bnCM8dzSmx3+WwVaov2wiUFHVceYAhwoXZ/j2Lul3rQTJ1o+ciEZZ+l
Qx35jdSM7Tw7LHH6Dh+FUTxWKsxH+mIxgcBlK72mLkKGN/nsGB+tOkHqHDJbsQVp
UERkXBASn4AaFEdMcAKjAOR4pTl3oc7WfrBhln2tHfU5Sc2mxe1PzIKPkey59hwn
NvuHnHkWqpqBPUxnUmuOb9r2p1LOidFV7HWR04W2e5sHg3YOcTSmLp5TitTelh7s
PLtX1oXu7PgrF9qQymIu2Bpat8e5GMwtweGJDz17Klky7YEOYTlJwccdnxNw8BgM
kAq+fK0dwuZg5pLKtTrr9LB5W5Ji53MtyIYYUKICddhszMisEkM0Dn2NvSpITdfC
QAmG06bbV9AjKONR4wZFgiI5pqlrGcXreg9uXE0Rps3ua6cdr4o38Ev38yEupFQ9
pVa7xvqPgijkLHjC2cWRJe+qBAJjrXT3jru/7bKJv1DUX9LUPmurQE8BVAL3avP/
UE+c3RrCh0oNrPeDtPCDewv/BDiZkzO4UDWCcOGi742wW/cygSFlphT7kHfvA8dF
rJnw3oneX9284MrQpFOOa5WUt8NcKBFKGno46jQ4HKhH9G+VUGtVMadUG9z9GYb6
T360fsCv6APPWxOE2fEvJ5fuyvhyIy3zsQ6dtDGxQg6zg1Viio8PofNXtCTIDTlK
WHhyUFvC6e3LmIkxiKhevDvuF3iBTuf6xTjFgm/BwGxin2LsWLKFaNUSxrYyiO/N
gL5fQYt46xRrjxvXJfSOySjJl4hN6CrZ9zPHVmKaUMdSzpEWPkoF1RjqEYdPWRnL
nUx4x7v9O/rdzvW0slcE/VoYvPNmRN+RYtw5CcyVMeFbbRyiZlh+ehyfRHXYS0Oo
F6vrrDkW4Q37yM67V8UbeG8oEZzU8x/BYAMsreG15zKUMYrmRL3iT4BE4ZWfbeyZ
3B+l3nUXege740dB8iL8VXyk1dlJjhDQat6S4WjuPY+cpO3QVw1QhbEtrk4WpI++
u68fgMGSdqM1zCE6ziEe6zWQP4adSnVNkNhGnEovSkzFYwMb/vBtk176Di2t5z4X
qENZ2IcXU7Lgu967TE73L1PnNqQabhvxZfZaQ7xOkkZEj4yxVPpBFU/I/tROHdJ6
0uKSAqBOe7z6VnCq0b9CzVHaCWa6MDVxUCv9/CcSezH8QlubqmIsAK+KqEJfTvdb
eIEmOqKMT4wSyZLn+S2ARgNWjL5rQhKyRaJh4/IziF6E07ZaBFySt6huV2HK53nq
QOjIirlIhmpN5jb5A6ZuI81gnNvLVn+QOi2R9+dVAAgr2x0B/7okCQ3s8WdhL9CD
WhA/tNgxmsGXSbsrIwmaidFJFf6f/EuA63DCG3paQDl/1mjsDSXAtY59HlLLDiEb
BqVPkQra/BppsxpduQnx6d/E75dcmj1G+ysqYatdi5ujKsFWq0zNnEPsQY2XYs/e
1Y7ZEOyc6f6llQx12VxFErFfDog+02WFrOWmF4B6OYG3+AVZFBrDNDP0UH50tRNK
kRvpmtMH8Di/R64WnwW2EU4xE5VLgOb/KMq2iFZO/ZnFphPFWQB65/Atq9NKhbEB
t8H3d0/BrTC2j3DtJyw1vxgl2M3EkdIJTuNzy+mv0XqRHwRojQLx0iTMwFw38vIl
wiPuQvPPOTER+zJ9l3GZzVnybFQTNHi3sVhyuOa8oMHLvt4N6q18M6nipBB7uJ7M
6oL+wTD6gP58vpeO6V2b4gurUCRvTR0ABg9LPPx6xwPb78rOCXM7uEHg0m6OO4o9
kwsGfSo72rD0W4BxDq3T72HSkZUSEOp6+AFVu5a3ENAAZ2U8EY6MBoRB9/Lxj8Gr
rgbB6mSYv5cQmR0B0cOZb81GuUPQ5T47Q3WLHew4G2v6D7VRFhFHgBQuakTwe9nz
zX9rFlrvx+RyF6DRlh0Y7MmWa4oItQDHbYQ7TtbMxwMdI7UD+NS+Lkp0ZkdDDFQO
+ej959THmyNJhZVOQ2JW6Y2jaFxr2tIyoVpSg9hDCQ1m/5SYvw1DEe6DK4PDooym
P+V0u7SrCCghKlenWy3lEUhDSbjDbpIxltBVqEY5UxjxCv2SbyF0f7QMqKTwjrJb
d1Wz9LFxLp4B4aCU3/T1/ZlHr9o7yNNVjuTGxJt+kv3UFNb86rL6hmw/v+mKX7My
jix4S4Jvzfg1HomUsrQA2SpX39J3h1kF7MuAifL6vzr09g3fgb6K0hzIMyhMaxVT
gl3uHUhScSYh25kDrOV4/OpN4axiRTgewxbl2ZMu47agI+xsbSXLcieIaN29WFtP
t/hoE0rrbaQtDxEiT2YSo1swyC/ZYSQ8LGrUn/VcbL84+dFsBIlwi4YtKjpU/cgE
ZH0EX1/sTfd7Vtr24ePQIIC2OpIsSdlhXLFAY2lemoEN//yx8LJwoqe31+eqacko
wCXKKn5hDbAikRNf8n3qqOu8tH2y26z3qnJQBh+RDUYVyMPnVLyuVkH5EnWMLSOx
YahXtsxluWgjxGtZUE39DaamGCRGzSrosvDLlEgKQll2j+CmqzVSAcyW8itfHL8O
7/iUilTlPzdg1aS9Kde6pdGb0ovoAwBPgQuLwrZRXUh3EkFRRcYK0XlzCMfJPTOq
UFiDMdBHLIV7RhBTJdx/yQweJ/JSTDlS+bco7TJ2Nvmk2Bn6RU89nnMvf9otyhjn
/xg71ncGdp5qbAOKOIxQu04CB77z8Wk3nvh0HBug8izLuiOxZzu4iMcUcHgNKk9J
xECE7A/F+8bq0Jz0Gp4xMLBYQOEOs5v7k/r4EqcY9qNSvAdCY/cS2cPrifExElL6
2+Ze+kbsNqJuklT+0R4KlJKCY37Q3YFvDnvUkMEJGuPPGGANqCluSp42nBuQkpEE
tgq6SyB+9/kGbhF42G9OgcdgAQBRsiVvwrd4qL2BTHUIDHIpgMmQ+CBElYrJ75mk
x16fMjc0/pn9mtqF/tbTo2p7uKKWeq1gwy2SElyNtfFPvV6keI1UmiSQBpu+h7BV
UxzElBoFWl2x9E8BJiupy2RYwvfdTObRYUg9EnPDIX6/Gcihyi9GzE2nhHEevy7J
j5GBwAEdHHjZ8LixEfieAMutIaBHoS5blZdctyjZWwqUayqiOAzaPSLyryi2lBOE
2fE6zMPthni1aejsIIBkxQ+Tw6UlRicNZtEZgzgjno7SHWVBSVqVojvk9/DIe9C/
EO76UopSZqGRW1luy3qRPwgz8nkTDApMBoEb+ER7NPKkeczlclm3gnJezeRyOhPK
ydR9oVK0usrolJevags4woQwYs4YJsIGTRIiSruHntwjiP1ZoDxkGWlNF8zOQtkw
C6uP44x0ZSfa1fWfYaJ0zBaZG0uXIHb7BpiYN6N1egY0H5fVh06/Hw5ItlFMG+2o
ISsJOD/Hm6qu4syfdi0tP8b3DkH4k2k76QM080JcKUH5XEKIAgOgIyvdTnN4Sk8E
6X7Fopc+X56ahAFTLZZeU7mfUcSO1O1F8dHH3AcSWVganbmcEfAo66HB9dJ9vDJe
ZWlEJ2RPY9ICXMfH01JoUbts4A5/HIVyHYJteEKnHFBhC8WcyjnpWjjoXboodrnx
kng39fKio2mc+efOYQLEeSBMjIEnrQf5TKT2PRADgEw4CDWU05xLbi26l1k5gQSj
V/usQRixptMkpyVDbDTZIEMUNBJrlIsIEvrzjkyZe1wt6wY3hk4yrVQyHIq4eV0W
JPqR1reQAjG/OkWQJIMfqHImQ1+a89UPOK2g+XfqXNjXnW7c3F8va5LkVfn0aRWC
lwCB+fkjS8OoIHqTLdJRnfIynOVZKetixBoJs0kG+u+LX2ob3X/hHAwxu1Uk50U2
9hK15PuBV4x7mup7rZEsO9TNyVOOPmWX/KxC4XoBiIa1/uEYD4cTifU5dNNcfioI
RHVgDdnHjZvlQ8+guePcfFdHnD9xKCY9UfGS35m+VAMUiMR3LeKbs01sJU1GGXY6
gE1shi1lbBI0GvhNnpEGBgHxGYZ1gItwEbrcv4WAPl2gZjQYLnl4pZAheHaeyf72
macY/JH2Ktw5KTh/m93F3Orc2scuXK2/DA0GEGjygfLcHznZFWQXaO8cbY8MwgNu
iqyW0bDax9yYHFPkds/8j4ZecJktjtnifbaMfOXnmDiFqOvSmcZg8MyinuSouovi
8NdvvkTG8nmHFqxpgOMIUVO44FfKuFPWivqEW5kMOTWMzuFI8bYvK3FVjfYCR6KX
enzmqmuLQsMSBNP+/nkDigo1mp1q1Zc0729kMhH+j5eAVTwWQ+F+/fDniNMcnjz9
j9wI3BqkkCWvSnVkZgZHCr2/Ge3l9PstWJKIPwC6J7nHGZQYpxDNXAsRmu4w9tdr
E6P/HKqumQrvzkI5eYEnrlI3BICO+bFcx/W+G2cqg3/klGgIf5L3IYMI5fZLVONz
GkEdcRssGGEfpZDxnP9bNzHLa3ITYgyIhSc2lIbbRAne1hsopBvVcHyrh69ekrU3
muDScrfcQZteA4X1d4xSE/+0Y/uxp3sW2j0D1MsrvAsGNixTMqy8C9n/B320FmrP
6KAw64seitYP/b/NiE95vURiGtMHfF7mYKgfB4TH43iV5nxUNnmZCPWLRYySPQu9
81oweuEjQ5PqHGHevLj8IpKCovMPmdB9KRzFKX3LqCzlVsFloc6Om5wWVDKItCwg
STqH6AAk0b2zgbzZ8PimOZ3srjABt/12mpPen3t6DAR+9CbsnkcHgPxPsGKmIACL
oKqqFV113STDEif29iq2cS9jkVKDWJ3PHGJaNjHc+aBPEcqVCP245dbMNNCQrSSi
SJ5rBXt0qDTC3KyH9QYCYaG36J8Aim4p9pdvh7VdobbCDtzjBCJuq6QENVIaCHo0
QOihVhUugX1f10hnsAKzmIbldf7JJzrhKTSuHYJMM0vNWlp1XQE28dy21iiewb2e
v2upsEL2W49syaIKLLUoqCCZ2nknsIIihkrI+/6x0zc0NZwh27sFZ2edj1xI4mZF
3GpkM23Jg5J1d4Ak/UzWR+Oy58B/mzXogAsNb0delbWTWsEb2B0gIDwN2gsQmBRT
AEUkL6Z6sfw677GXJ9HLsE8V7O0xQ8oyt4DcFcXBZsn95stgioJGAGd7+U2oamSC
cXUcI3Y2vLefJ4nDwIXM160g+nKDMhoyTZerr9gScGLGZ+33ZPG8y9nMjiGM+I66
3osHIKiyV7KuRoF/rQsHpb5N4VOH3PknYIpebH/5+wg8EWpv7cYo5nDq/1mWYedO
VozcvAR81O2JFiIB2cVNGb9fQGDS7nQ/xMYExRJmsQ5fTryMMVxfd69+2pHBFN6v
s01WknqaKWTP71NN3tGRbeP0dUvufbUmcVndcfMkWxsCYHA43DeBVcLbh+nSytxE
jzRFgmut23w06WjYnETdpzRdaqInt7bLe10gV6krif8mMwXkDd7KfetWCEco/j66
V7hb6gtymmFOKS7UP6bkHT9x7qGWOfOY2JG1kPjJVKu/LzZldAT7CoQiiCvqpLIv
p+lYqVKloQE7U307vQl7Da15Iv9s5MY8QeATSQ+4Im77o54F1xXo37tXru4dIbmW
vmrwpJV9/jZrMoF0QLUiMgTpdDYvPNdF9kCZTO4myqYpEScUC0QlXNuhlq9N1E5V
vu+WCc4fWPM6sJn22ZZYcNDSzSjM8FfMnxGUn5m3gbASAR/ib5256hzoUoEpEvNX
en0RoDoykshpAfYd0RD6cc0/T3tElEHkjUVnaoshWb9RzMQfUKj9knTKw/Ishwd3
DqoMr+oYsx4ukxeLQC8OD7ikwYQkSJ0H023BCQHfKrGL98M0AqrztfDgvUJJGgMm
rlKrhJ2vqbV0NhR+ccr7fb2+SpQyAV61WkSCunJSTaa8tLkHHYXOMEsPJMFfluue
A8hgZYS/a1gDvTkubDegeN+ZRxbqKbDoDF4UcekZMROsmN9S+R6TYraQqXq1p94S
dK3eJ2DQBA6hr5uzbnfPCZcMH/v2aOoEWz5LPsZOkIPdjRcfdVPy1M1Sx9U+V7nw
jXAIYIt3msRbgzaMta/wODlyOkFu8WN5apgqt2oXbvsNKI+3MlqLzdU3dJYr1a+H
HdcjiuwOSjKy/xcvIXWHy4Q4oEEzYUru582UyozIG/XaWUS5Z8p7+4B/xM5yq/UM
MMICRS5EfC1y6yak3/PiM1uCHe6YW1E55Z2TCAWRmBJ3jwvNcaTwmEt9Zt1AU2GU
qbLWtJmYmTsJEE6NIdLQqQbMdjSJKDBy/FV3mnNAXNS+eWEcr0U7sTKo+ZjxuiF/
AKl9mKV2SKt/wQSPcwYpmuQ+mQKl5PwmERfTT5TehEH40e+jR0J2Fa8b9d2r1yiq
cmAPtKmnvWP+rGFoQyvuJSDSPgwOV85mfhmJAALED2mX4Vsi8YjA45XCBoTdTu3t
Ws0Yz5iF2DXIZedWoMV47Y3PA1A6awXlBo0qgmGwpYWI1/j4zPu9I9h3FZRGW5Nc
6lZd7A96Pk3kQi8gy0QKUq2GQLj48rEay44aRvXc3Dc5pMLiY7NeqF7OvGpE5vBp
4NQgv7q3JcN62SbMsVKfnctCtFmIygvHA0k3zdYhxIub8I16tta5LagEqlsvQcxM
zLc8+bQVKVykBXDPa0oLS8iVsRriW5TEcTgyiqWmDBF+xYoTlJiCGHMUONcfAZpE
qWoi5GeGJ8h4u1UuK8/DI//ZWs4Qdv4DHeYP5VfN7OVVBvgJ5TDfj/k8kjzpLk1q
cKnfU9qP3q3VI43PVqpwvsf52EAbWCICO6/hTf9AfmGbbsdbz5UO4TyUeQ60kFVl
R8NHDTJ2wMdQvB6q2pH7nZh/PU6KPbHhk7wscBKwyZMXFoeBM8kuoQ6QcCmThg2C
IVVytLvQcaEMeBreyWz0Tlt6IOeoLAIHdJl39OLBNi3/FptGOTuqEOA6qwsHMzwk
NVxwyba1LXo3JGbsi2IGA4IpsIZySq/Z1F00j7lOkvp2Rcqq14w60DMZ4q629DyB
zkWeAQIZqM32ETmvI5nbUPI7/c4BRW+mTkbkQYYiBVtF9j8igqFU28KxYz8jp3BA
syWACPflOAyteHOGnadMmnHz7DnB8mKum3ubA+AU08eLEiDHj/VSfcOKOlhJ06im
Fy6j2SwAD8xT31nbyzhXTtfBanBUew4//ymROfz98nM/aSV0IKOtHNuOHAJ7EXmk
bZk1PKtuc/T0FX5CcXso4YDsXE+3ulwDN/4ek3b3GC/kTyMlJlqdTRaYIDt67TFQ
+rJ7TVKnUXd8pc307/zbYGRMOiDy2EVE8Ppm+kmRhf+o4uh1sGh0Pt2ZgEXfl6dp
MTmYcdTvnKTBHFbSKx7urO/usqHuA4nxXQ/IdLXIDMbUERewS6ZdgcdSPh8BdUp0
8zyS44R9O+xXRxm/PvjNLwkhmtHmoy7ubtqdbhxAlkDE6zZT4DJekO5zRb/uuYvz
siEWs6G4Ta5ISHdTcy5lkY/KJZISqdrHg+MDhEoL9wEbWbV4TmMu4gaWUV1jEM6p
ZopipZshY0GptMKuv8L4w0cvciJt/3Hcll/cxrv9dfKJh1+xciiU8AbFJw5T+xQM
Rzp+E87Zamvhw5bsWdYDdH6rbdngM/Y90asJdzzDYDUI1opII1JBouMaDlFIvH5G
I7K8J0FXVIArVeY+nmF/y8S9ibLNJzyPKPDVs445iT6EoN+jk2lhQ/aQwOeEdpvy
QBrtYSnDTsxHLY6PLHGgyPvkIpbdd4TpHG+VRU7vUhpQszK0nStcR4Y+mX+mGzLJ
aJc2PEsXwEGkio15vuvNufr+jSVvqwDjPBOpWNdyVcClmALymJEtgVhc+Rdb9Eym
Qj1LC7kP10pB3nWaKsD0rN4urE8MGpQKiNeJimgT+b9za+ZMm47Xk/xyfIBGRf9d
IrksAL9RFlF0lU1dTDkBjWpXPno6ZFVBl6E4y5LB4Kbk07h0/GYETuzOEAxhV0I7
8JbqZOvJCkXKSP3rAtBn/Lp6bAFMX0hmeOXwOFEOjBy43YeW7Pbd0pZCrDatUMpz
cYbwxawK96o1VJJEjiTrCqIBOYaXDDj7Ob8OfevcYhROgRov35WCc160kIvqOaV+
FgwEHbV5RUH2PXEHw0X0I3vZMLd0VPOMnbdgvYdD4hTYn8oz1RY7BeUzZFNAo4Ig
ge6NlbdeV3te+WyHZd2Nz+wtFk1W3DgxcdjejfioIfPjjzxLn5tWq0kFL7IyZxjj
v+rB1J9fhsBTb6Uo3L5yOE6vAT85cEVGc1YQDzWdzi2uoWrjUo0O906We0F7Na7y
OOGQt1ACPAH0xhK7P+6fOnQOlfeEvCuRxCiYIZUUIiaMxzqr9ESIoE7nmKVYamWe
d1tNU+WIQppSAtZHPpcao8inPi3zxPnqnkHrixjKXXV/2VsZcByRpSgzcZO8A+hw
G68dgPiNKPMBUA/PRfANaTs/ZXPvnOdCJ0KQrprx46+KnWSo+7uEy7miimb6Uf0U
JogI8G+HiAEsqc74w+bIZvXc4Aj9ZgPOKguD14H9A4BB8H/hUDgZCArbeJ+ewcnO
0BJhUPeRxN7Lmda2uCRJXXShi0uU7g43mvxde9NNzwcJpPUlc+rR22h/u6DHaO49
O4wNPTFlsgEJbrDTebLJuZfBRrKlwZk6/KrGBoqE0QCxATBgNblyfgMNB/zG6IW3
i7KTjedBr70TDX+rw62xtoCNxJNSbJFeFTM5tlRFM6gFmtsu30TFRXhvtY1H7JBp
XN12kSc+L0gpjIBv+nbekQi6KLOvKDJ+KgnD07KVxXp89kygy+4ta/hgR4zqkrIa
mdGggnHkxo3Go+TWr1l6Qh9Ok7wh7eo7XEW7sdQeHeA8kg2nRTKd2++3HrxF0vTr
Sa0+PLWH3sEGeg5979UChnNiFG48zAIdEj+g2t+nWBhpBzpHy677LkCp/XRQ/kue
UeFbyOU41+K8fYPJksPvr6eLBXgoUswNrhPpmDmN1DTqyorcfTxOUhTHv5KJANJp
DNpIzOZjvCmFY3qScPYoEy+oqVWp5A1KFtqEePA77sM+9qmPmTlbjGIyqybAzxir
Os9wSrS611SjqXf/qSxVfKr80d7EVciJJOXJaBxWaMkZ4GQsCaqajyLMsiqMyZKm
d5issZOFqJPzh7QuD6Gr7WG33zltiA1okYTC91M0DPEkwJLhvjwrgbK63raK5yqn
YTef7hMXpnQ6hwDbWi8CLpnU+qFPF9Qjo2mBqTi9Ueqym0Zx+NE5E2jShRxwwQn9
lJXq35AH/yHyrsYhVFO0o+aplctQyo/Z35i8UoM1yMPfl2bN2ojoYRv3eUj0Bj48
vnCrWQT5fB95jDLcuj2vCcUJt7lgRRoklkaK/ZAmTEJWpAWJ7gV0l0KwU3QbkDMq
TrwPJiW4vfvHuFc0f6k1X24XxS92CAWQUyRG3/W8Q59OIBpGw/YU/vRKywGR/KPm
jUC9BuQXjI4LI7DZ2hf/VOgkp04gysNW7HWq7b2UXKW7IciEU5Gphfyd3fJR2CEN
9DZ4J8jetdFgDsbuabZYKr1L1+lkFnInBsKBd9eESbK/Q3D7ImKwu7EQxljMbOgl
Mn0tYxQZI3LuRrkx9trmbGXAKrV0mtWtqrO50Ns9WCvifIvXhnEVop8bmzcRDtX7
hKqvE79srfH4PwlXsBfeISYJNezq/50De9snLFgQVwl5vqIXnmtLn+gxK1VUjftn
H/vzCrKkhxaoApsTlqtqvIivLGzLs5n0yqM+3vDd6T2HJBOWGfas/9k4BUP/XQwc
Rl27K29r7TS3CIi/pHNEBDPTZ786VRABgKSW5CCRE8h1Di5WyL+jUmwlsYO+/9US
U3HfO0GnVKeu/qCcA8cdoSTvfKxglaNAl2U45g0sqUulluRJhgjtGwgUF2LOf2Wj
YY3YmHTOUyA1AwDG9nFDbKC523TyeWcSG1waFRC5ZDbKvJTQ0g989rCXQzsY50CB
6PV9X9F00aNs1i/fzqjIlIKLDK5sM8RtQZoBv0ASrTAU1MkIPtJRnM3poeiy9ZR0
H+N2Guaf+qOShPiYXoxyr80+5XqqE0qGUwMuG1d+J8pJ2tW5ODdeRbCR7kCKuWzi
CpCzdM5lzKCbJ/ALPNQjk1umJKLjr5u1470GupbNZ1CMVbsnQubISTaDeyN38Xln
sHX0JQrVg9AmovkeqtD3knPrfkY1nazhn2cJfWIj3c30TNdGvoJgAWzvvPBOkKqZ
Ir2mwVh6w3TT0bR65Y+RrjIUkrtDKs5BzRY1NpSJWE4O8LBOw4b5e8+wt1DJ3+BQ
p+x2X/S3xd6/eu666FrxsrEdD++vC6YnlUnjm3v1Z1jMSuE/tL/mmUOLVFsJtTnr
fKybPDnwRqpCtdXekuQQ8N6+VaEZiREyQqAg96IwawMA8YZdvVaNeQDyRzFVyWOf
uxdN0d5qF+ctXP2UGmDYnRkeH8LgX7WdIF/T+o/0fRojNd6pwE2x1TQfW0OVK3z7
y0WF4YfWJS6iUhP6OFDaJvLdknOj9jGzBRdMqCO0znV4JKFV+2e5cp6dUcHUEJXS
gVTgPj9ofoPZ8Lov16o/R15a+vF2KOGjWTTuZMnxH9ap311W7HO9mNqNdfdhCBDi
8wXRaHrSTLg4+zyDMnzBzBjx9VCbojh5aWT3cvdCOJkphF4MJqDh0/sKRhNnOlNe
oD/LwLDHJrlUYBRKC+fHYGg1hCAxFG9762NNe0OUPEdMTvdCY7HOu6ys8kOmemiI
BGHrmENk4Ry1f7A1uVIfsZ4Z8l24Rmu5TMdfyLbiqD0cqo4pAoJznM6StuXvHl2B
W87E2ohlAKZUCwHTmejQrjeBDpEnezrnbPZCut5TdaI86AqLrThMGk+xyEFBQq8a
iRfdPcoPiULgkk/IU8568178dkw2sYS2tkUGlGdfa3jJQKUu+5KP2vs3aZh2WuHW
q/V8WAK1YYCcPZHGS/9bmBmkMsw8B6pP8NfveBcAIdO8XFqxvwGtzeWDV1dWWjaJ
YIWyaUwKDJ+orbn7Rsl9SJHlOnJtKWwEZzlMaB3V3c73h0tCaU2tSYdBIg9x1FKn
IYqCjeCoXMIxnSFA10Fs3k3lvswG9c9ND/quR/Z3LzTXbJ1HJHvNaxzcCPUw4wji
20c+p2+A0VdEAVCCdQlMouLlsegiU+3oPx50hxDRPooCHKEtb+VBs7GD8OtBZ182
LKNdCf5TH9lVJCjqaaWtB3UWulxN/fC4Sq4Nlh9lY+bw7G2ixtwlwvFBfQbbJHwc
QbIrozp6GbCJbwBwi7/rCs8+MEk5LabaNUqNFVbQFCSbZPsQfAjogjAPubkvAJ9H
nnBVgrgFqf4RBlVAmlGzQr6NA/wJe05lyGB4uYI9c6R+panGRt4BV3ZXYh2p57PF
oeL/Jjvaa7vK7k6P33etKkjvuyQSxsfJbd8q9mS1MBos1bJUkQE7TbTEHOp/xbmi
aBi9wBicu5uBasLXuGiWBwBIdwWdy6dwDgSx+XwATmnj8wX/+D/rZXzwwYqq6xF+
0rVi5AWDDYKdDm4keb9SX7EG/qxr63GD7CIKfPOqSuYhYiYHydtekipvaSHywkNb
O2RDIqg2x9G9YqgJGs9TbEp5xx2yGtJ/+bSKhT9WSOFuRlf1dbZMOapeZpgjfuMK
yK1byDwOblwicbpPZT4n5h3m8vdZALZWY5twTO06sz8UB80ojdHFZvv4KkOwLPz8
OZxY2FTkQtcH6raU4J/nLWAaMNCWZi6EmZHjRHbaOcxRwcXXS3f2TV2irFrvaIBB
Z3j0H6RcS/k5nEz62xhqFKdHcsUulUuYmHhM7b8y2kQHHj+cM/k6nq4QBsQO8YOk
vNwWp4rmUfSIqdcr/8GNbTwpCbOsV1ox6DT9Nqx/gsLWcNpkkNQtp5+FREZ7RzTh
K4ybtAje+jC1AyL+v5PDvY2wdRV+LnOi12w2bUL1NbqStf7CVuQUDBsV6L0Q0O3s
8YD+s53qvcnexGaerc7nvhycWuWV3mm0ihZqcL2keoCkl6AFbaafRhmhD8l4AFHL
kzCLUpzbTR2BjAAUPNTApqUEBQl/2nWvHZzl8CnZpx40fkrjjemzAp50Br2jy6xD
kcOdMMX+hMe93OQOqIkosMAOthVz91Mhl2eEDqyOHCcj4NF32tCZYO0c0S7OjQNk
gV2oZ/dOkB+mtIHvjRMUTLGhV7GqLKYpcFA22lmneCEoxH72j786uHu0H35GCBZE
r1f8hm2uMsyoHaWVEkS45RT41D0bLNHtFfXLe1EE/ds1ASmHKPPAWI8hGylLkjGz
5pEMrszHYuF5v1dnVrfq/6jlUkIB1vTGrThHNaRru1lR8zOG3JfTk4y/wRG6U0Ad
An797ppdMUDiNd6FSbvG7sXZQJa4KxCXrJwxGIlm2EbiJanx4OkJ5rcI3YhSZw/S
wLiN+BHmp9+tuskDFuIaTI9gcGMu0DoZKup2qrYLjNMLhlOC9sng/PgAqifqy89G
Gs7vtSmTR26bIb93cWRyR7Td6ZBb1fPtlOYO7yNljsUACAJpA7m1CFvoWkBm45zO
2qgKHelksnNT34SxljpzCLZt820t2YKqU2POEQ1ofBFx8wu5A6dXhlRB91hjdXa5
SF5leRdLc8LZCdcG6o6S91kejIfnlZqJ6HTWtGVrSEEBg6ROzHk5jMdSLGmNouPM
4Eus9zYbOm9ToKmtlDtLN5SvDAg5ilhvZVV0EU+rbGgDQv65kCJvtZFaq7bvAbVX
rlW5Y/DvStDFQ6AXo0W4ov9F3aV7hyYKL99BcO88PLcyQfC/ClJXkKNBHtVjW2ku
s9KesaDfxH+ipunXVmdZJqOTEYhW4MHVFFP3fUJGWaTdmvbdwBxKlb7Odo3c4oA6
IOHyzi3aaLSqtqy1Gnz7xI4f2gPMqAm0NJ4CtSbeqsNliErDIrc+Iwd9mhagC6gS
pe4E+zyg72VvS7D0B7Hxr/BT5TPOBGDWSPsNSjdM/IgPSfXQpV0A38p82KWqyF5n
V6epTpnr3LlB1lKZEE19Dk/wmPfgAEArqN6UVip3vi67EjP5Hd5jEH0463iSTnGd
INIYJhHC3pJr+eDs9DTgsQGt5Nr58owZOVoUuh/zUuUEzlkQ6kb46G9v/AHWPFyB
5KRNO50hH+Ig+2evT956b6R9pvSQeZBMhT6hu5/e05xALcysb8KhttJLFpU2W65Y
kR6YAZju76/tQ+ReVz3OMqEOzkkgegMGJJDkZP1nbH6MTkNNwSHl528QJmj9uz4l
dCdxc4vIvH6Uq2/fqHfSQQkUsRBLkKyr3nzqAcJx5uwWtg7F/gtdvIg34/GZYh8j
z3RFcq9LqtC/z4Q/YUy0XuWbjmnRKCZQ/7KcVAcBVz+AkdoJlVQmnLwq1e00xHMU
Ocfu/GPTR7056sp24pB12KOxhwZx8/LxaIfF9q5Bt5DxddQEhZeYjJ1JJGripfct
C8gIazKXg6lQW8tQKSl9gmaGPU8ru00AJcEvbkygtX5CXX9HOrq/t5PHqFOlTHjQ
A7Mi7Lcu5TaYiVF5W7K9Y+C2tGCf4PSCXC5m4UEW063mLt0LlLTJnKIujjU2jOcZ
idg6agSoQyq12F3/HTtwsjbKEGU1+Bcq45b4Vkl11VwM/PSBIeQ/oEAwzHQCs5tR
jv0bYYcZ5XxpNp1d6AiHzRe6FTxruhYGppkQuvzD+3+6e45lyS4Wq4Lrxoa8n4br
itD0u+9CRh4Mw0ZOsfpeudrW8fhSiTTK71dPWkzcH4/aSOEj1U+UCbDQlg7xKOlB
Em57e5Otv5rrhM4x4CABwNkX35VLxJv3vIb4l3/FRomY6qI6v2mT8clCoJalKOOk
29wrOweew8j/nUkWCUmI2TnX71H9vzwhmDrbvyXyAPxEJ2hP/dn3Xd7NyXteYqfh
K25y7ggEahpmiOoFIrjcxjo+ULdOXz6qJ99iD2TZ4ODlzfb78R6gg72fO6Mqq+vK
MhkbDGWO0X0WbLoCgeOp6le+5PLPJ4y5Dm33gyi4u2jNYxGxD7WFs2PO/dLXX0Id
tFs65L+G5hQxiGhm84HE1VAeDBXKYwDYxgABruJRj5iDeNVMJkEfl0NMtK+RCDrR
dM0HpUleaK2CreLee83nyDtqck/IonBdfw/syIZ1QKilYTWUKMBmVUQd0Xk+L9aV
Fx9pAyIDKEzTeinwRUU/LhT31rnp7yfnRgdMFb+qC7wE0zPUZdj190HmRIySutPC
nZIAnx4DvOzTTn22Cf2wMKvOauDaogjM/GbYUPmLIfHSVsTsVN/tM/zg4dNjRwYD
IwxWh4pr/6zc6+CDNWIGw5V3Kapw8zeA9qhoBADum8DrNXNXAu9mjz7jjczBBPoA
gsiVMKbdUZuW2KwGWz2ijYU5+ZVVW6pqHPCHqeV3VgL2euIGFCIKeB4v5TlbrqNp
dIwklcCkv5HwRbiEBgVpszeYVi8oHmpJ8M1VpOZFIJXX7zobBco5Hll7C2ezJ7FX
+zQquuOuDxWJH2Ho/zjtunTrzustZjiEK/H+11FmnPLXFg2Hg2S3At2DYi747afJ
6v2W2JPu6bKm6tQTeoFpP7PLl+l7eXnhdiu2ESPUZwMFeak+KyspsXeWmnGYqrG7
mdW34VZ2NKMw2m0YGadl3ApUhMwC1V7Ce8WaQSjUkcE1ubt9cvB6/egacUxcYopD
yZZ9A8pF7++tN1iMPxPcufirPT1U58d8hwsNo2O5GareCXCutGAhZpIzHF1GPRkB
LKt3t8yewJHi0l2KmZt5MC822hBEaejxDc9TFJktn1kZ0hTEiIbNeFmRCn5aVpEn
c2S/d/b/n9isg0kIFBuZuwN5w/qyN7eeIUQaHZkuxqTcCsg9t2ORTeDrNMal6qYB
gKSsGqnE/5rJvWV6lN5+pTG0+RKT+Y8EiaouRSxfvLSsKS90lIGsDSHqzL57eW/b
Wq5pVuNdXFC4KvIEviDHIy8AQIvBSkNK4rOHektVuQb5bMbll6eVdN7+djbX6s3e
CBunfyb0FkUDOOg5tzeAWQzXRccQpDZgy9HYCyXNg16VwV33UxD1dQMtZ9rCVebr
4TSRnkVKfaC75ox1VVJOxBASt8EogpOObncJlDV2cf5YoqsH0fZALu7T3V+OkQSc
8yKCFSs6mHrovHc5XbJPmlAPLXwh3XHfks8lj3sCLIzsfOkC6Pu2AixRShF9A/tN
Y8qwZEKii7u1hgyXaxV1UQAR5TFeh7DC2+82/vyocWA6i9mqwfbEEJCiGxPutB+N
Ej3pR9LcRkN0eSl7ZvCSoPTUtpzrVoNaO1FV9fbO/YI3NJ9ClqKVUjFmPEGtd2Rr
aJ+JpxJVy995t7iTeXsvgoC3iKmahI8T9r57KChywQHqab62ShRoHVIGDj6d0K04
sqSoOpoeF5q+sGrG5YR9XgCCkfYY201vw3S5qYUlfPQxrzvqPWmE+70NHW7742wN
4IGCTO82qnH2d8n0hUI+cJgwHl6Rw2l0W3z+M/PyCiBsh5VpNZ+P1YO1rEMX7Nfw
2gBofTwGZO+w36rWg1gIZ0WvO7elzKfJ1YbfiIs0aWKvRg/r748yTlMZ+U2GeyU7
syHKiHj9yJowwlrjtkpzV91ngKLephFx1TMhTPfLffluOe9S0S4FVSTECIc7iAbI
ipChGBOcm7jYYuQKx0wLlJSlOyvrHxQncoS90C7fk7RX/aSr0BjodYy+jnJmSXwN
8dmg0nvqia4+UXLU510mV5MqLbAMDh0M1B9ZGYuZcKX7yj/+GxPqrtq07MfWEH1M
mTdBgxm1W+CKgKfJgG6u2H5UNdiZfvPut2PlgTEdoRV6fcoTLTulqEffUGSyreod
7Zxe/p4joPcdEtt9DGf2pFmcxrypQCKcBr13iRvXBmf6ikpyO/HR/E5DNlfOH7dv
WH4xBOXf/4fkPGUvJQ+DmZKnnFP3fVdnS3EYEROKH2nT6m6DAN/6GexozbSWLife
ShWwsYcGLAG4m1/lT2RBIQ1JHC2MAvJl/0Iv4F8nkpYHcxO2OBPIqZl3XCelOjFA
wo13kK6mOyhVmB1lYfcvY7pi8/wlF7fTEQFmaispijMG3D54EQU+YnscRlAIfyg9
ov77Dpg2z1Nr0E8fn2cCcdcmndqjZ01wzIS/5c0kNxMgegLHvPFj3cM45jJxzsEi
5/jMijIb0AToSgSDTMBzZ4wEPpSCWZHDf65Fh9V2OwVzH4IudlDIZ/Q5KDLLvFlb
Xnv2+9lftdyDDTQOq46aXzS66D4xTkYvwzj3SIBTNJtN1iW3qig5rng/rmkrcwPQ
tbUIZ2oHYnOOLXawKcLQ/z44xkHyk6KDSZmUYoOh7hYl6NzD+EOJwt6DuF/4y45z
TJwIMA0g6TWOofsbv8yE09rznkEVqB3ahFOWWrTbpsIvIep/xkOdNnyxlagREwW1
msKIEVcotwkS2pL99M8dMCC/Z/NyYYq84B87QChLYwtoKYNdixqOK9r3yo7tR8mU
2hcDBOEgwtiGljN00EUA7UMnzgXPM02AaLGcZbZUHPM3opApNiM0HhIvuiWFYsxd
bOVf1583w/uC/4tjZeCy/ChIf/GxnJZRou8mBteyPnERWUE6UEQmQKjiXlFntPL4
Rew4QpEWG0ki4UOy5A+HTCyoBXTSuf8ofiZCNHl5Qddf8QM5KUBu+4R7XaNTmMDt
wqu2YvOZ+Aob4yIWRsG00oJmw0RuXdlKHu4dXtUQQDk86VpSkxQWzD3IQhNiC3oN
UnpnL4PjvbDKUvIwOuMaXiHG8Iu//fPIllVwzW6yODCvixKM+P/eilfJYDmSAYKk
gJBjkHkvv2IYgLvFpbQYMSwrXWZZj6lv9T3LPv7PfsDY5EAbksnj2wZuk+8amayE
0/2h5sXChYqnf3JuhvtjO7dlKLM1ldcUOWYx9fEj63U+jTIXzqtRIGljUVzvYFrA
fZzu6+sNLS4muoCsn5N3AlZe/ZNz+QAjnHP9qOOramNN6gKz/928XoeMyPNS2lKt
IwzjC4zsLfgWDzB68vS6KHDQlCIJrNXL1PWtp1SYimNPIGVElu4MjF9lld2Wx43s
pBHRh74Yk5cpUeaHCIabWiUE9ayTU8Fm0y/bFtsjZy1gLAl3OwxDQrnfndZLua2k
t1iv5GK/SWUxF17euy5xOkrVNU7E9Z9A/IF5RVnB4A0V0XEnV+hzuXjFWC6KUZm3
7/v+4/tR8htUZDaFoL5h/zM6b+raHCBKUCmIc8mRfsEOHTj2ck9dBtZkA43NAW4h
TV1S5t+4+RiwpOHk+oV5Rf4JsSIZSheuhhXYgn6w236vKEosz9Gg0y/gfkLtFYaq
5sMfj5br8P4JfqCFmpqSKvobhF0k4vBqOfD+ZMECmxTJKHbNxaKcjx+djwroE9/r
iwcxuU0l8mmZoin0EuCfDEkx08WJ576K/b3wF04nlJN74ipsC2teVhcJ9wmBaaAf
Zjyomho7fWKCGEiMlhZUxkitHW9eQK9vcRAQLFuGOZwSRaQDD82a1QyiMThhzOyU
k/iWlOw+sYgYnLaKplPEklzOWb+VGJ2bDMSYIkRrDnJcf6Q+X5DmbkZyPAuqO7F6
Vo5b8I0zq2ZmnOnq0NTC8ODrIdOlwbT2zmfc3V6buVqSJlXzm2FEb7/evrh+f+B3
mfrwRobycr2n2tm8lwiNyRlV420hN4W5rVgm1XeNjH96cW4iQ71sLgmBxr6b7Zs8
fmInkBwIgOik7+OV1hF3A3ryemGsIZ7vdv+hjuR0vmALENAK0Vg1SRpmCp8ogG+j
vh2mlgJj1l4ii7EwS2bGCJB0EOhyWSkMvf+r7wiKia2qQ31JfFr1/Siu/CLGDQzs
ibLKiP25tF4yQyop85tpaqY045zbb3YOJqboVKcar2flQFejCMJSInFXwLIh/5aK
ByM1sm+G8Qu9t0NkR0E806qOtFt7c+psrFX8o7n5GCuxG/uKocMOSEieY0Qt39Gv
Ul6ZXwXlCuccI1RFEb6nbNyuHYfWMBvLVm7IF1vxG/Np8KA52I7+Dmm/cB65Vd2O
GN9ZdCTVkEzDHvYRFeiMCUYCbTk+O6oCjoAm/ZA1j6kmrUfR419+bDqt6PICZLZs
axD2sFQhwWQYdPEsCRupECrsm/68wHm6D7mTlv09k8siNmdBawTu9FHpOi2nFQyz
YjLCTmosI9gGMAbXXAbkU3i4E4i3fgX9IdyukqsYZsUzvOswmTSxFwpowTE8EVth
QAEg7r4cUQzqw2XCaAl4txfbHSvdZAK3DWqG5G7Cf1NH3yk68UqTsgaC8cvdOdb+
zu+n/BBVoFEtvlW3Xyu2Ad0bU0Y9N8F+HDyYOGjAZx5O76QFfuIBbMSs2NDa+xm5
+P4CzxSGfqLrnAVPVPGj33R8Ve59cvTui7W9JOvo9Klh0kSU98YGBgzMzQ2onlpI
BlHJlnYVHDbYw5HNIP6uC1DrdkcLomIHJUBLoemUJSlqIiZeiBlY7TcpRCIWoMB3
HcO/qiB9cYbT3YYEcFJBjcT5+uyOWvDY32e7sRJEHQstJg778qDJ3fqIgiLbpsOR
Qn8pMzJelTlY46sYd8mmBF7c0wWoX7aWn6CfWPViIiUAcXF5bUniSeBC9EzdBbAo
JUyWW9Xkc4p/eHcxTpuHlznj+pE6F4TzEt6RLu7J4JFDZ+ztfS6CzYfgBH5EtBQK
8d4ZYD/rEDcvj+iu7EEJu9GTOAgz980tFYmJoHCuTDjyZRl/Z42n8Bl8iTPkzgKS
0x8OMX6B2NBhtpCJqNHlSXrfj9opuyQD5Q6EK0wGL4FvqLZi0AEoV80YW8fhbt+8
5PxhZpmUE+FvJeO+geWZ37PSEMfGYfq6md9EzyHNR4KiOXD6i4fBS304ziAZZ2h1
7GTuQlzIsjAQE74go1a1A+WWj3SWB6o0INqJpbkyonBsl7atDddzn9UiuB+mxuJM
TDj76ZgscDOKasVg0FAJwP53ef7gjMFGBPkdEvFZbDg6STXeeibcZ225bXLScKyx
gaIdpJAmT85ZSzQO1zU2MDKZPZ8L/911CYu/ckqrmNIlNpQqxvkfxrnAsKsVnygd
g1thS4eXSHx5WUpvqmGh2+pPTzGUl6VWJANU9FI4s4jW2OPWQI3p99KtrmqtrnD2
b+Q9vXSux/yrc7QqmTncoc6aIv+uhgiUrb5BubkbPcbojO4mmlsBRi9ZiobuVNQS
+tgjU3MvKaqwZxaXzGkyoJW479qrYzNAKnvLTvXum4r/M9UWJZzFCajelWmBEp9i
3HBzH/KlqCER+JsQy408pnBi+ZUpkfEK/YyQGU3jgsmSBDfTs3TH2cl5O5Zr07YI
m2V3k/V/84VEYwi1wwBZ+kSYJI9OYYrpQgW+uWFYKhTXEbPz4f0+yuc3IkTHxzM7
IxVLVXF01E56SxozNsNkEpQKgce9x3U8Je4W92wd/WJzO71d0Amu2MKb9Ei+uX2R
h5Yce21CN15IWH5O2mMD0TdvdKQbSMyN2ZL/Qghnt5RXChhyItJhw06ZLEwaPBhQ
YYqlnkfiG0qF+wqxhefg8ZoGG/xzuZbGRaisDC8/N8ltwQo2YHuNueFdxWCTiuC8
VS24qJJcEWPL3aoid6MvtSAvENITjsFlMadvqyI3tTQSxz+enmwuMF2c0BMnd/zW
A/qRm69LaCec4VB0jlPBqXacyMPs3cJDA0u5kIrbT1JZ7Rg/zCS1DgPEO1c11Pbh
9PlAo/KAyDl8E5fwifyjGShScZnS70Aj+ta+2yAH0jgvwAH5KZImCxfymupHsMF7
Ns/pGjOdCv/g1o7/9at+4CZFZeJdAJHXn+07kn97eOAkvM6iDH51mRhykYGaba0G
4UFyFUi4hyYOsCGhPMRK5dOlT97zYlw3hPf7KqCeO5bIr/ArU2vjrrNK102HtGUt
7kyklwEJBlgdkU9071c87eN6uu2w1Nod4izkqbrd+uZQH5obTSfLVyNzENL8wXfI
LsWC5LaHmgRwSxm8j4IgYLI3df43l1XGDms1w+xsX2LahlUDB9oy1fTdjqL1KQxz
4/0ePGHdJN76MSiWaj7x5z2u4G7d8euYAEcvLb35xb+0WsghwVTEUt3xpGbaKBks
Hi4cafQmCYHOs8zm3yC3V8EkitpMG9rh4T1kFGtDiLDtly5mtytaCpDBTCokq0EK
s/wQ/X2XfNGRbuMwuB6ZTTou5/xCebxqVMdCNbIPmdTjbJZ6tfDtSB2eTZDI3YGm
OiO8hZJx2n6gMeDfE6HnlRnPwL+QDgTvdJhWJUj/FEN5JqGdpjbk+XdiILSsAcM8
0viXhf4SFc/iKe54aHIzA9ZjW+yog8mlZdiEVrOvdHbv3oG6FjyWVKNp/9+pXalU
aHbLrehc3ALU6aK1pcQc1mAC/G2DFQ+Smr9+XP+7wPnraFGmw7ZxVSh/68OIw9et
SzAeDepX7YDIqEi5NX3R0BCGBf7ZFNDAYA7pz/96CpshShH6LndL1TOuBpCsB2Wh
qsKIbfySeinELeSBfn6RiQ/k6kNBWOd/DaIi+PpeFOXZ4dBTryqUaRynzXllfBDx
XSQzyUF9yDJylVDSlz0S7Ct1UQ0WlnJr6mGqErXXqyO20cGjZp1CV3qSaF8hKek2
+Z1yvpy3rioc7KRrM3lV4SWPDayAmuxZFWLFXcC7zkhmpp4zu9Hxud78CHQ2s8jR
d7M6HWVwpKTVhYWherp/tAs5rRqZalw1F4sXoEEd/9BtPEaCxmagJm3RyKzfC1Ou
zqqgfZQLwzsh8/f9emRmyY1rW6KAqrxV7fG1e54akgxbFY0wbQhA+g/yupyNFdMB
bvZWT+CBRLMrz093Do0NaSGFKX8FO2h51sRpcRrQPtmNENeEHVmZiUS01dp5PJbO
NBoNTPD7BzJr4eeVX1j0a0jC+c902EoiOi4F9VW8lUarhwNNmNUZPdgRh7N4Pyrh
rG8hpCc21LVYCwXexRq7qc5gNBDfEdO7qgQUUjFmUVStxpDZZ9P0YRpr5f6BBUZZ
NgFj1ASLzSH/u02vr0TvO4yrbWpDHH8/Cxv7M0x5MRsibeiyGPWPbxwvdGC+lvRK
sn/Rl2CI4KpDwPQO6cdIBJqTfF7hLeirHfkeJ22gxyjRz0TYsv9JAiTJwyDOm9ba
VKwi3kyZmZRPgbr09COv4T7zBrutbjs286SZxjCPUgUIBPuluQYukEZ6bKRJzrlI
Pkyh781EBXJSyslbtlwR4lZ+nPgSx0BzHkhdmAiKgebW4Vydxv+RbBLCk5vAfKTJ
rU2kH6D7+kBi3LmFe7so7BNwYCWebjxBKH+AQ+/LKgcuzOhLiyN3Zm5u6RHQrfin
1UpRKCYr4fYL6KMEtpyzAY14YVQzq/XIYEaZtIrkx3754gg5dcPLw7tLWdmK44Z5
vUIMtSglp7u3aAmBeTbUNMH5s5rPPakWwYY0/61DeOrxwWYoJDrvFMoo2mHz7Wir
V9vIUkSDfF9E/yGg9VWt+aAWO8/T423fAoMQjccp+LqzHwKqC8TrN2MRAaUYZzFc
r52PCQh/ytAxCeT+Ejnf0TrrfZrxLkvxTFPr2ELs3m3ojpGaFEhbq4t2UIAXfZ6v
EZJ18PnePulv5+c2oK4MqalvutuxGHfLTjzbjuv3FWRMpz+BG7tAeLp0J+mE2piO
p09hqApHEjg0PtyGb4Kt0P84lv8i97PEd08kJPTkopF4wHAp0RKrpxojBd+rYWHW
9LzsL0D8zz9vu1UXLDtfHY1+PPOpnQ2sLbZocX/MF7VlYnoKBEZN0KmXFDdrOR9w
dGNcQe9NNHvavXb4Z4oBJHUE3dB8xE1YFRZuxbbIkH3fHMqqRjlJM8eZ1fpFJS8c
8vVKi2XcZE/n7Noogvqj6dfeWay9Jfzmi0ABtAEECkuhRm+po4dqmXWbvR0mJ1Q/
Vygluda+fKaaLj8n9t0V1lKmjJOouof68bkIRiFm5FDqiHTfd6628zFqDrpA49kz
6EGrUjyMqsrhc4Jp/dhAGt0WmXAeH9BP5ri/WovQghSgW5UzwmiNyjd56Wx+vidW
2xwHgL8Dys0/DaoDQ4FG+YfuxIjPxyQRHgtb88cjWzpdnI26hipyIK2GcbnH+mO+
cPNqJcsJnx/pm90ZmDnS7RW4/Uf6uIMjGeej5oIY5garqWuuyKZ49bU59M3jbkdG
7onFb6GhQWiiaD2/F+rlLavWNphyLWaqdEXLQxCsUDHCxKleCbn87x3tJt+DPVBu
01igfdPKWcabZnfrFqdC05f6uUU1jmjsrD+BvF5sHyXGjnvSqgdHQk8k3RCmriYT
U9lR2SCB7a77Cm7eBClLp6zwX+BZUAfqiqtOIwpHgaUP0/MG+8O1j58gV94jNoCV
y2Sm+tXQwCMS3Y89Q7K84ZsVsE+TirURrBTAwmJSHKMG4RSymbEV55qh6dJY189t
uEQVYt/0n7vrAmE2Ewclezf4vAxRB1TMwlLjNVXRo1WyrNXJ2MlVsls/HhKWlL6u
VrPw+OK1K2WpEeLqBPYpHfy/FqvDkX5PQLDz3KatS1o6noJpp0qk+HL1v8HmO/JY
28Hgg10AvFgNPGo3z46fmypPPcnzKhzn4XHeXcvOzGTPXjRpLpc3YagGszq4O81e
/FpyOn3/+pyhr9+anMSlQmwKqNsmuLjh5bVghlo27DQTfTb1ABcZmowMkP+CCz55
QtrvvaaNnQYats3/Hi51BW9edRjQu1IoRuMpuGl4Ep7LFRF+gFr5ImQYIUskDPfB
fgUIMbOPHE29lXK+rOEpMqvfHEGPHfnz7rqCo+ECRAohQIPXZNBNwz14LQhxSsYy
eBewhP1w8GOwTSX1Ez+0/W033MCwbcY0vFVzAkikk415dwqpyJUoIhy54hEXPzAC
v9h+vciksPt59dJI2LtwYLCgdYOwKNTcf317muby9ztfq3YIWomuwiGfdTQO35Va
SENXbHqUFxTOwb1s/McqYptnFbAKsVsUQWqS6RZ8x4kMuRXFveYXviEiI1N9rSry
6ThpnXRvHpqcCsmXL75uPVzZIzFEZBEtyTtKlA12WZyB/aUoSZt9dDTyc7dJ9rQE
ysfdm7jo3Tker1Rslw37nlhumaNN0+tEutQu7Kay5L8rakiAcixl13ec68LUFnKy
7rkTelk75pTju6BhboZIcLyLnt4ZU6w7zk+PkJSYEEj4O2tFByJYa4Bhtq/yY8Es
C4u530OLC9bF0VICFPyJbRtQ+Ukd0+rV6klBm9CObV1KiWwHN6ivJ5MIE1+8yy+E
b6kdh8Vn7wg1nl+nswQR1zykL+y7I2y4OI2vZHb2ha+G9EQQ+v2ybpljOcLlbAOW
jwqKWmu2oI17gbmXpLhir2urmHI57vAg+uiOBbL+OiYDPCwJ+77209jpGtgBPmjG
46EN4EtIT3iB6vhEqBArF//MpDl6njtTqRrwZIzz/Vnep/YAPuIfNWlZykxgVPno
4XzshjqkGmzfY+5SzrxNsmHVsfr8UOcy2iAw+qhrUacRBkOJpCc2zalfLIQDSQlq
kp3tWqXq1S7d1btc6WoeQYZZx6XsVRwFTet5zaOekMjbncsH+XIAhvhuTmYIPmMx
z5BaV2R1u4oKutzjVXSfXnU1ajOBA8CToWovl/jZr7aZK5oObAne1KHs2WEPt7pK
CWMzRsWrCA5XpFiZenCNufx1Frac+W6etcGl3XU02CIkMFev6hkEOSqdnIdyhlG7
0DoOJWNJfyTPFUOQ/AIPz4ueeSlIM/uNrTMNQ+1tLEbON10p1mVf1Hj+OBLOOV12
nkEbwO8eATbSMVVSRMgxfWSxSMfUCKDkiweDEHxW8oebQiCOVMq7LMFHn5ypHFtf
0MJC/H+TzwP1cbnsd53dQSVmUIKT9x1b/Ys/ngImItJpdJ5sfbFdzazoaspORneY
l8q5TQgMHe8KWJIjei2fQbiSgJqEOsqssf/cHPVtrDtVfy2TU63tkQ/wScnOVdP5
NCPkQNoDbCx+kixW5H1LL92mPkONvYYe/3HLA0ekXBDY4V99/qcFWSxZyY4uAQdS
k8BXBlYggVcmege84gQYyf7gFc7rWLPA9GfUnH9ywkDVdUpwL7Vtg2kXeinB2cyN
uF51PosF9FfPs3PxE9P+xLJbJlyEkWbzaZng3mApQ7HnydMIGU87tV59QFTuhg1u
P621raNsGFbu1w1ItgTYvdGrc+Z4um3G8kfacsndrG7Zlc8Jpp6M20Eprefav9KO
6nSTfcEOOMohZS3SE7S4a8eldaw+0Ow8zIlRbYs17TBNRltWRl7Y6rkzBdqzXnye
wcwauHRpKsIlRMs2YAAqlQxLfAsQvRC6NYQOdeAgQ5O5Y0wmzPQh2oz26mvw8dDq
fZGNdirKzkMXc/HeFx1rVwhcisRtMC6Lo9a5zKTPt24pPuCiUUT+dlEBM0hmJKYP
qo8IxrGRUZKHxmxkV12ZNKx2i4dCz28A7OaCOLgJh2RKgHy2WBIUSFmT+XQe2dsh
Lp9CLxXRqeG1C1mFJkTupbLgpsRHL3QC1IpZbh4ERQDJYPhEZBJXyBTj89rDLSnd
rnAZntsdqa8yNKNGoF5DCaYC/8YRv9WvgMyvdpQ6/KVZJ+lNN0FGp2PeLH+ocqJh
8zs1OOnZd7USzKs9A1T44zDZHLzzs736/tv6Ncr46GqULWMsKcXMaGPUjPxZUNtd
Psr0clZhW/FKZ6X1t7LM1AHbQIUBq9efSZfYYDNdHkOrmkjZpziIenz5Eqheq1dO
SlzvQkTaSuzX1dKVk4VBGJxeuUTEzotDDTF9e5UObcy/uZpPS+E1ktJCdcRvubZw
NlIv18ZrJBCEPZXZTu7IBhcpCwRrwNbSXlmhmqkek9cegaRP2mU7CwhZspjEQkp/
++B8aqyO7hFaDNZkGEh8k3vK2zZVcLl92BkBU+G4Rdds4AXUi21sXypI6vEzW0yS
a3UIYElKiGwBNw+whV2kw5BVR5uHoNslvaai47F/pPclLjndTvaEXGkI/AFAQkGa
8Zu0MLK9LwLqzD4EqSPKMhCM1KJgTNNV7rCtW0/5Yrfk17nXNwBOxiV/f8FoK+Ci
2XVm84VmvZhvYKCexPZQPFJmjJPFM9/MTJzn0QYMId8hNWmIFt5b0h91+1fODqC9
45NutJCOI7DF02smsP4bba9fS1KtM7CB7+rOFcM1AbSCvLjoU7JVEDPjpTBtTLKF
KP6ahvFgChKuMLt8R8Pfajn0hiELTNGTirw9LkVe1UYt9nWdBUZdbYr0RaS23PeI
NbZVdOWMKTqVhDfKEzv+Nd1BhmB/M7MhNl+jEsNqpnOTioXlrNChZ2mGQLwvpem1
ojz905Durq5wY69bLynNOwLpASKMfb2pS5D328RhkBZL0GN0nMUm4YvRG4QhT752
StK3sLRbxxkr/4rlUqWPOM6FzlpHq8jH2EKs4vMnK2A=
`protect end_protected