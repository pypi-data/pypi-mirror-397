`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQMy0Nic0oPYTT1PeBRgvHfGDa/OYtrF2RF81ZRbgQrc4
BBD9bWWBxvLwruISmoCx2jMcu9cgyGw6RCGDYtvcPmrX9v/cA6szpK6Beiu2FPwR
VCJocgXO0eutPgjhqmmyPXgifmEgHmFffTIf0mGaAFkU6ONOKwK5xKzBlv+NVkcd
jOvsdyYzXhPaZ+7Lb+859YFkBfgaSK6yQ4GR/eddSQjdw+Z3W0hrdIa9W6hOafuF
bOQaiz7qb+Xl3tNxcjBpRRoOn5F0PDrmwk1L6hq0X1IdsUfUsOQWhHt/+2mJy5dU
IgbSoX6k01wlfpypBD7O6n/7orjl2eXx9HVGMV9yFaKB9eNmyOK2QhPAsfkigy95
NN2VELxBqLl0qeno80M7w3Y9kALMPv9YOK3wgBIdm/u6xyjGXU4na9JLOGlkpd0R
S9vJrmRo6or/QuEM9kRiSOT0QX1BB3aL8L45RJIgyO6O1Jqq9f7z42x/XvG46i6V
tuaoT9lz4Da4LORjU2I+BU4/iSAD3UFZMiVsQe2g8nyOp8WskYnkjSCVpfhQYFUo
bNHyBniQPg1Pkjzr64+t+8+EC8jdeeG8111jRITyo+S08mBMjzHSzSEJKC7YJi3Y
U2L20qGanpnG7q4ca9F1fgSqIWfdCRIfe51eaOhxkzsTcSOGkZZatPZYFHTl7bEY
XGggGqWvx9pam3D4AImYsum8PNpn3V8dZKbSqqfex18+j4jIrofWdwGewanweesS
s1Ksd5XQexe973ZU6Oi4fZjjm+Vc9bIcVu7X2uU+KLBEYML4tjylfhjgqLVHD+s/
ARfpSB1gZ5ywlvifq3dpRdaw8nRSlftjikEzxjRGGQGHxyKzafm8klQTtjTq1DaH
hX2wXm9wLcoaDRD7Lmec6xJj4q0QcIhFWEUKjwjyT6I3NSp6oPUSrj49U5JK/2l8
d4PC/9aVPBHFPnJCwh/gAHvn7VEZrvTc3QciN7y1i7dG9qDxCqGo0ItHWKRSIxOF
v3rSDs4/rKtRrPKS6ab4/LrOiDPMDG3KW6lfRq0LCrmR6YuLATBkfgimIQhfezxa
jLfoKDvMS0lmE30IzbATAoZpPlZop687Y7vKR5sgzaq7p0DBXIFLYNag2ktSx/20
NW+sT8BMKhtMb4auaVkb9nhEqtQXWuDFqRl4khkqaoEMv9VnJorJbPDXYiCkjEun
gfesAJ2M2SnmcTF82UOLa74YrJfjp6TivkSY9/WqrEe4xyzBY0q6SDK5LQIw0ipr
IhfA7L188vjuVmmcTArVJzKruJvamtU7E3LEfYdwH81au645BHFt37YvAL7dwwd5
uWFq0slvw9j0bahNNH/8IS1gV5Un1dOzooPvF5u9G6CqGl73ieWLbE9neu5iN/Rf
HBU+j4b8N9OpdQH/DdQ1UlWfjTBf3spTvGQSzC5nRA5QKjNMFwRIUALEZ7YR06Do
o2pxy9iCPKJFgvWI3uwMX5HHQzidk30acmkMbamY9dzJTH/djmhRWnmN3x1imElO
wa+S0g0PrAG47TZ+6yavLnuMjZ0c6FA52dq//lr/nTwl389gbKB/9ospVm4GRISt
ItunCFQvDcUAda3cvMKSCVd+NLXne23tc0EDhrHkpfy1HtEwOXbZhmls1JVHNpck
bOVu1OCBG0af9WbZYvNFwUDCzhAhPycefPMv6RRigG4Oa7QsiIksP8ZGuPhciXDf
+2cj9P6UVh1leyp6unEmEfMb6yOcyLmd7uoJwn2LjjHVQYPpFhXkOn8Pn80Q4Je1
9vvZepmgRR14fjeF1Z9LY9UXE4CXxWpjxMHtOW7pzbloq9UY4OEtFm8tabtOk5Gy
PaXbTMLQLqotBuoz2EMmFwm4zaEPR1Ubpq5Lf09cGsHaL0xM0jjAQ7C60OJEAEsV
JxzJ9XYy52bPPeSmztQ9xjpA08jvaoXYSppbHP90yoAXS5oI59AzyBmfAf96htwz
f7XvaVLwqQzxHJgngkRs7QokG5YBlXEZe2N8/T6aBnmIMuNEG3RCVkplgkoZiDCB
cD8PYMMEyy7+Be56kKDCJPJMhVzqGFdHkNO6hMubFlvEc5wvvisAKHPIZCV+aJb7
dNPY3q9+Xr7LdkbrGU1CLKEH2kY1t43/ayraf1cznpm1E8oghzN5LBJ3ltOfmYbB
QbJ3Z4MU8pIGmeI0/ftyrAWlDsBbCdyoi6lhqgrq+qZ2F2/2mgTkSEF/W8Sro9J8
rrfWF6RdexHqmXSz1aVc7lhaE5UWUxzbbTGcr/kYS3JJDVUm+CUgUFo0AdvtoKHH
6O6rutyghqoKuIdhpwNcdT9BPN6+RFRzL2PsNGEFXNY+7e9CaLIQ76PVnX1SLuSK
6/Tg0N8BS+lsoL8eF7/6CPPvHN220wCZg+ITEH7UFXUcR6/ltrOCOxDvHFlur8E/
YpaNUjTRReeMmbdlF1wdmEu2w7F9Eq8dsSpE98KvQKTgj1Xwyxd9oI++Zpi2HRd8
TS6kFzFYR0S6KV27NcDjKsDGbvn3UlhpuhLgxlWzMasXMqDMjNpedBrFDvH3QPS/
0T/9DDWbkBpswmwpGEW29eHCezM/08lBFnpXLYAbg+/unHmPB1KmLuKwiBQPeFaA
7pzXo6yq8KmWJWMhpz4hvBtSa2MxnpdJxP+sZuasSPc95knT39VxRoDI3VlpYFpb
IsyvZ+ULQ2NxjvEP0GwYxiq+WPEkT+0aa5BfXhvG8+1/3vmEqHIU/oI2zma1Ty0c
CNmS59radKwosTDN7ZF1NIQTQRb95CWvjrRJ35KGhLYzCMCIlylkZFLtTuln9raZ
lXY8IEnF8gVjxUNxz8OrWA59BQUhaHpzuXZfgW01BKYQg4mbrwuVZwTHPhOkHZAm
NrLSaDW+nVwXlislZVVZr2tWyQF3jkLiUJ5bJsg8mtGRfZuGkj8ca4FXMwU50S8e
5CHIj8GXeP3olUqCoNt+RHcIh9bARc2lYWGIKnAuVC9z9Bf23sT8lP/FWC+pWb/b
Mx6HqN9pFE1pWKzYLYaAyzzqGfVXDlypNw+OCoUh9p4WaMiE14A6pfu+bMEBTz+a
qq6ybTM4XZi9p8jTGr9MqLBqkdTgyXKzOt5PoBkbg67kQse7P6IvcVt2zoLgHsak
jUDTJr4b1RJCgRBoM09YgXAMaKW43ASYWyN9CpgqMG7Ak/tfEOzpI4Rb2CCQ3nKE
0y+IbvTGBY9jtd9836WlnJMJKGNLmOCI4XXe6URKSt1MlkyLVoXZszVlnkXWi4/m
/+3azsey2Fkr2vhITwJsSqIGiWfuVzI2w1jvODB9N9v4XETdO7WjrNwmiwL1dx3M
8gYDyHHBZusv1qqFYBr9TpYf0qHI8+Spo8JJwzafmUUn7MGmn1LPv+vNVO5hPiJw
txwGX2N7eVew6d4IK+gRdOQSPytN8ErlN6d8twn0bLQiny2LViVyRRbeSoAj2eZ2
ZLGytNPYFUG7RkFb83pogyOIG4AopKZj0wShNk+v3uMRfq9PWtmlspHeDUU+vnAT
K4aPp4A9hELWeXYozMG1IWuxDUKhRQpjMxYsdyrE8J4v16XhT8plHIgQ2yU6OmnN
X4rb1cPxnLii1zI5y2EUTtBjmO4L6PGR+SagSvRgDxlpOkPmCwAatHjUCyBbiiY9
GVLMke+79iznwoXSTq4cZw6KBzPot4KtWCa0L08yon10FxRKLf6UxVZLmiZWPnSd
B2+CnxlkPsG49clvgc39rc6jbgJjCwDtyG1t7Ss4KFYfRfKN1/liVuqqeTzjpqos
uGivYnpYw9H4mCdEi2gWdW2alAu5pnY0pgWWqAd1NBKF43IynpB9Few6ulGrcdQn
prVyjU+DLOmK5kYJ0K2JPcrhH/NtmpHvg02p2PwTas79WRrKMLHbUVl3P3yVLTc3
3AdBhdoXVdz6TnaCQWK1v1e53yuX3DfDWsnGJiwOIfb5QeeTvbfmzDQfDewN8TOD
Nqzvdwe5o6Q8vQnW9likVG5jteLqWep0GgfqX2CLa55Vzya8XkJhWTH1VxyGA0Cs
39sjlA7UOBsP4uDhNinHhaGUzHvWEfs2HmgfvImiiBwfGPP19tZktm8oc2NeKgjZ
0JjpjhgQryxKTC4CTvac9LJiALhBWwCZFKl7U/xifGAz0/OPM1uEZ3i3efOXCltJ
BhN6+1wE/Yxki1cOwbmq18up64glffZQLLNekQEqhCTzRuiS8nI8pfhE73MyMII7
IqK5ds/cvnGwB39FwNbCA55z2+zqyQdE6lqqKBBHSLKH/rqeBBXnk8/v/eKcwr4y
8qkdSG343WVGriXST8mpMPke/GvPDcmZQZmtiLaegsdb0xc9+PuYeoRWGmo1GYOy
4d4y85IjuLyt96QeleF9jbqh6NCB6lQTnUzMzUzvuIwgMz3K/+uTVybR6gU2eYiN
WFA5CIA978fNgcYgmwi/XvZkGICP1y3zY5G6oKL9nYU3MDARsRNRE2b/T/71KEV4
HeBvzEayCqSrc5JBhaATe3zhFrSylFttu1t1iPwLhKyPqQHOndcxDxiXoTazHZwf
79BkUuUPPOdf2+XJUqEfyk/FGX3WcEK3Zxlwv+ww6u7bkqA0xLzncjn3n0/i3+jx
axMbXKF32GmE+Ajti5rSzxmDQ++99ei2pWGMJMx3gNWkUx7bv4G26AgKf5HldZkJ
xYRDStVO88tZcm26Z3t9OmxTe/mDaHEc7MnnWBhRv5TUVSgay0eFNTdcnAzckxYY
5fASucYjL4+MddYKv4UDi2NnHiWeR0zZIrXo2QLNGE8ugnqKWUDov62N1lpuksTb
Hrk/+LEi/1bojjcXI6a/A3uF0ipMf80YHzwWnGHrbmljcYWnBzCV9OBsevAqBQjJ
d+41l+1JC5bkJ69obGcSaMuogBh7yLaAU07r75MuxoGGQ1vBHcuNG5w3Wj7q50nX
ZUrODDQSL64M2cnQYPoLvagMZOXhyFwPVWlDpo1ZT7RwmSH+jtmWIxjmawqWk7iC
GvQdYJ/XFScsLvZxUOPiWNR6qQ3tvV5YIoH3zGHe7P0jeJtU1TMKd9wJdM+DBaNh
br7cvQ0WtY4QGh9iJ4y2rXrtVVZ3arjCkQBlYL8rjXi9Jm0SRRbP0TDiMzFccz27
p+xnb6P55jC+AR+OGQtPIV6HKpGJPKFzps3YcG/ueTv5vrA7fm9Mgbm4J/cAAGt6
eKlV5s4Qd32mwQfpRFAw7DH54k/3BKSfhZzAiNSgbuS8Bluksmn3gvgCSIvv8Ft+
D5U22t5wVYiLaszhxaejSvAFOZwvLwfwxzyTH/2CSzI4P+yiEyxLUUne77exTIQ1
Skl70N56/URoidov8XS01jcjUxYiagGPbMKCcFksxEH4Qst21AUgdolszTrDVkE6
z9RY0XfycJfXuChalrC5G9trUYQh1QOOL6hJ6v7AJegqdMKk8rEo2MWgPUxMTfmC
XFyNsIE6lqglw5ISvXiEinbumLr608Hf8x6RDDYgmudH+eL83xAyBlXf+OTUfVwE
9P+aVfloGteU3WME4TlzBDI+Df6U5zk8KwBXoI9CYbml5zjGMsSQxqopjWdZJpeA
/IsdFCqgTflF6fypAdb6Ri3EVfv7FpPZHtnjJe30D14Cps8rQ8miXaQ75iXzneXf
5y2/jEna9z4/54mQlAETSzBKTanxIFcAr70TVMjn+djU7Dr9cWPHdIAHt3Ex7cqc
ZzP8ZBBYLpHui9b134edJPLJLrO9gywNYMjAMAr+tK3WVDkxQukJoNo46owqEbGL
/9r2+w2wwB4ahp4JE33kQ8FGM5MqOHkyUFzMWPXderRheoZfmQiETyrg58rwTuRr
fDKUuE+isaJeJKVc/qPpLW8qpF/kIJKkO8EZRyVmVAra2H7npqu/iDw0+h4nxPv1
kkHXydBZl8IatnrJOKquWL5lFcn14IuI9mbZO5+egElNeGj3S+aTavR01qJuS0+B
v2X28EuWYBnE3CGgUQyKSJEipaVTnoxefyY5+1BoWxWjlmWQyhVOE7x4OcJufyiE
r/8R+LSoMw2OzUrktLXnRsa6FiBAHb4VZT3BCP05LZhAPKgGqBTClhoNUX+VK5KU
1IPJaXzz3Rz4HiQVcJaQqPgr6ZZ/p+gq3uqdzyUeK1o6xGRPDplTNZEt/PVbiIMg
sKLrZCMz439+NUNfUCCguBgSD0LmOZd2NN+DL8D2wGskOlYLkMhhKYAhtQospA7R
HMpCNGiai7390PY48udzn4vqcjkRn6MHV6gXlg4hshqd0VmdXjywiblrkI9crlIw
FYBbEeH8AGYHTT/tyfNaZJwDERcM2z6N4xETnp3z2GeCD5axz4Ji8vQhwz3aOhsK
73Em3Sihb7Hdns84bO6KAdQSC5qHE8hK8pWN0Cl8tUpbr4QV+abJyh7kEoPNnvFA
XTKebEyD0iB7ARPuZYXXQWQ+d//R4yiKBIJqJv4E7OnnxJoxN4HiKP2QK/f7rC8C
BQp62kYsc0IDaXMAgon75OLKWiG/cbJ1kLD1afbpSFe5E+ksNP8rleFEBwa4c7k8
9UiL0yG0TRqnsDihjtgPD//jZ4KOoi67ImzJKh/y/p67jqaC81m/dRqQSCdflD13
dDURSlAyhem0guUCPqEQowBeGfKHxQ4NERen9nkswt35/zQKreLnod4NxVRT8CgS
4kdNZn45xxvzoJwGBI/qrX7bBDCY5LTsTA9TH3qgbamUx0DwDAYB03vEdgwH8Zez
Y3/Vr9T/JMtEWr3LI4mwFS/ITAT6K6cG1tZEp8jBJmsmuzK1irt1/W+on01pNQYz
PPkfoP/vFcudpTpmUP0XMuOyiJE03SuU6BIDR2oksaslDSFsScez4i0L4NGEZMVf
uJP5y49Kuau/6g02ZqB1IWQmpQBX7uzo78/KxjxVfOJaiIau3aoQNrsfP/XhXAai
qPcWqfgdHfCBSr371LBz0UvYW4ZVM8qBevTwyAtFNjVwL1u7bRReEQZ8KSHMzFww
xiBMOmcqT2aVfudnvKpxm1zrQq1jOaV/3qVNz/Zn63LILY8apzFKVYcKkVmLXgAn
pJ3Pvr2E9fj7jFrsnJBbppSzL98eJMtkbrc3O4qfpJoZlpTk7BauBKEuxQQcQ55+
Y1QWpePKpGXUZT4wrBItZWKstkqYMHU17D+JdVV6bLxJEOpfkhWXgg7lVUR4sN9O
zJ+NoHpnGqdw9zf3mhLTiwzl890Muwkevbn5MWukaa6J/fcofoaeYTOAXOTg4PN0
vY9IlkS8ArMKdavJ80jpiW7tNC1ZdUS7kZhCgVlhTadzp8lCgxN/CMF7OG+X3eWj
AWMaW9Hm0y053Otan5FzfmX50PUy0GX3HrRyApd/NSXode9QMFM5STg+L8JNY4Q1
F8LK230OfeRHjEyKRh2pdvrlOQ9/ur7akZrZ9le+54vojwk9/DfHmQ7TToyPw+zt
g28XYyZ68SSTIkx4L7RvnH78vkEjHAn1RfflnDjqH5+c6LQhMfRYODP9s08lXKsL
Tjl/34f2lIn8fKr9eoDMeVMCjaNi/hammr2KZJBeidZtn7+8kjbXwQX+UYvPFAh6
XYBvXc12kpc+Kc0UM7mmuswakzfPSZ+oqHtnA7Q44WJ5UTXNflt2tXd75voHt6G+
Tc4WPUP3O4KoQBie3nntS+ATdfDqL6+WZGfbieAPWFc2QW8XhREVYHbIzkSkYSwf
w7Us9QGS/oFR+zaSUzQqV0ME4u2mG07L3YiIvk1cp9VnjNnKY8BJ/2iFbSe9zCG2
XZIS9UTX/OGoferFyHX+lxV7sp0Tzz7VVddwqEOr+AELLJol4GQih4xlUe9JFAZP
h6Z5V7pX68d6kvgFA3UYktT1mD1tNsIqZgKvX8MZXq0Vm8W+B8ZHFrglvQaibPd9
cWJ2DKdzfbYCPuRYgf1Zp93hkOba8AvIxXYgYNoJm/r5WkYIhQ2mWDbMXDqeu8VT
mMoIy98Jw1j3/fgSfsfWlheHMD76XBYGwqOGVLwxsERzU+opdBe5/ESvNpLH+J+o
5vO47dam0RHFE01vhBRL5Pxx19CZ5cpvPfrmN1HFkFEgZPYojPEQDqYoahwxXV++
ekd7b1vXgykeEIXMhsFBx40KkYEXCRCV71EnPyv7XRfNmymO6r2bvva87RLin9p4
dM7P+bIhlXwGglbJ+8WASr9G1RdFWEeNWAkugJCw1EPNd1f3jSe8/UoOa6amDllc
0L0nzKf3IiNOtpWjiPPhXAEsmCdAqlocGRx52mdYs1x3ExDZrhsPcU6qHh2tgBav
D2KmrtdVywtTRUmkizVrTX2rF5rp8GEebr1azr6Kxt2cq6n5VDVQQlXFO7yfH2s8
Tb+D4e94GOHzJ8BzKvwsHPoz04upGiehNrUf0pVCWq1hLYJ3y8FWxosJkyNnsoXP
RQqWTpDkrGMDqcc8Pv2hsQPIzyQ2cyI7TPZOs8yFvTo+V0KCDs4O6Q2IBYoXwlrL
eSEdOOXepN2Rbb8PjvuTiIlHZ1B4GT6DLEQBoyuprACY1PfiT+V04vfURMcyRYXD
0V2jtXAZX8PxHGTQVQ/TAYAGyO3iz34HmjwborNS/CiQfPJNg6spTy8FMwL7KmvW
eTl74guKGkeOohpSAOODtYkXXQ7u3MfNt0uaUFtAKYGK5M4YDTydrDCougKa85r0
SrNVtRfC/GcQ5NtOOO4UByvC6V58SGy9RTBInTZRY0Sqcn/Wx0Np1dm64eA6qeZN
cvZwfJhJvZnfT8PC6liedVNst1lyPcKkwygrnwpbSyg/gfwPpr47wEmxxf3/rVpr
WC9UvCcsTGkLEq8fIEOScKbRnWpz/Hrf0/OcuDg8Zrd8PTxvIUC6HkpRcUHhoE2d
VLcnsZ96hI5cOkkKtoXEOd2NM7Vq9sBQ/rN8R4hQl62TMHgM6Gh4OUzBjD/eQTpq
4bRcUpr0diE+P/ZY6VPLZnmX8C7ryC+onSgyDi45SI3GnKXygmkXCWzvx+aHHyoK
E5ha6MqL9z+ZbRSbDcYEBsfw7p/ih76HD93SW7lHln6KVzTFbM0hlvCzCSyfWuN2
571mXFyYNSSMcqt+KLUoW9H+8RX2o5LXanH7fCvgoM+ORu8Wt/6WaO/NquXpPsoK
LyFU8HvnP3n1Nf/sSE/HlU4DBjDcTCh1xkIDx9T3N8D4YSPX2Aa6h4ivfOQDi7n4
FsgyodxFAONj8l+r0uAPRMlzdPTnWIFty1s9FosjHSVC+GlTIjk2BxUcN2uFLsjS
QTVg8W4aY3gb53+E4flHE3bAdkovAVR/pORSZJrnJluw1g7/AclUspUH0Hqn9/OZ
PvCcG39M7USxgTE4cRImez+0lv3HM9x0pnKom1LBFkXNIvn+gg6ordQYKBQhMj75
+XXaY2MIlQoELDXWV5N5xDd4Mu+CF7wMrrfv71PJ0pCAvbDkI5G8iQOT8cs6T+NE
uwor2jr0xOBgnMb9uQu9elnwotkCBjyeLypQh2MV0HI=
`protect end_protected