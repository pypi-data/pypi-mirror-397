`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinGeoFAw4tUtLz5qPNTzj7T
Btai0kr6dutblJw/QBMwvDLdJYtv+Rd0vjXBgrx3ap/l0Z1heZZDAiVk52q2qQe+
yibNC05kE6x15xG1A6mXL4lH9aQ3s9bF+ehRZ0ug1wz7L6R4+hzCDtpwrsTvot3u
7aKHN4fkj9HDFJw1aR524Fw6ozszejNgvQMFvevD8RETzOC5AJZ2uKRP1ubcFqZO
Elnj76NF5Y4S3nBYxDqEKgNr2qxwg+fsHyci39sOIfXnkh1nEs6X8Wyp25Tl1Ubb
rs5ocvCNqoM5Vaur+axXlY8GhKh3EDx+EpEui8nsggNORAPm8D4St773Vm+JKCYz
DfpfKf1gWUxVbijzEGTJEhc15LlKlBPuOJIPhZXeeXFnpz/O4pH/PFrqcVeVpkCp
qf50rawW4Mp30uWS3rjZXl+wwKnhIPdT3q7la0MH/JdEjaYFiPWyCXR/TQ3vanBS
/cr2GXDTWp1tO2zJ3R3id5pSCNo4yaymvGdPipxi+jgyKMGnyuWw9fW+hCxsVPYT
udqmglLSrGQQYq7/1a7hE4lRa1JXybaPsl9VcjKiKH5Wm7G7/qfxrgc64w7I0jY/
fbiK+arhQgcftSplXVEB79R7+NCssGpL4VOfnq2P4FowzKy2UeV6uPonOu9kr0Vq
8VmHG8mATjqujqRIXf58NwoXiAqCEbI1oC4zVLl3ZRdw8G+BAOHURSDvp3mKHIqM
FNgcqehbmg7vBTAae5RyA0rli8Oq75es+WPl7FbLnUBRPNhUq5IYh610hbZLe8vU
js63ILHc59BI+wA/oR5TMGCalN9tpu6XMwpdjR9LEJx0QYdKP/HbqDIo6aUe36rn
UCgvi5NMBVg8/oxwcM+KuDA4KlZNAHJK0ir/P8rd7qUNtDvqpAB4zWmvyTY6fR5g
3a/w3fWNS/6bd3Ei9ua1TwloI5axlCcLGsI8ostvCSFek/lHe5a37w8cpzJXSxv4
A519IpbN9PwmKKDRYU1rVObBTdYmo5NfSEFd1xiGyC9Czc5wpVlFzBVdAl/OAivJ
ERbuB6ZSDaDCR92ZlFDjx1txDZi15002OIRePv1yP7UCrQ3diCXI5+0wR49lhZlK
/SR2zVLr3dXaAOJgvb449JlGZUHtPzTz9PtOg3c4cU3MeNR+W3DRf5jZBZOUST5T
2F5gy9FLVmigIhO2t0QikhXzSL0cM+pw+aV3EKIjqYoGNG94z3grP7ayFNmD4LKe
AZ/B3KY0W6qiAqkDirINdj/f8TIA7zZySj1UXw1zFay+6b+X17a+mVFWTtomaCds
l+pEmnDe7S5a0+yO4igdqa0YkFeKHLNQOFw7ku4PgCfzMMH5J1RCzHxroF21J+Cs
nHcRSmdCjljJULcKGCZ89s0SQyz4CbCBT0rYCJfHVc4vnumpiFfs/4JlLC5CzbTo
E3tSf3EMHzr3pybh6+lIg28fv6qT/LNjz2PfgSStpqeK44FqUTQxyvs3UsIEg6ZQ
iTBo5c3Bmm3KwfuyguX98UWQLHjZYl20ipCc45wyP76Q66i2JIfEs+kuCjq0Bz+Q
uMn1GiHeNi8gHI3Nd7YndW1j+vc4h+xf3vkUHIyKWVkIAsB2jMrUB2cdUZbnQEV6
ZDG0ffu1pPjx+yu7KtQEFt9Q8bAoxJcUTp1tb3LIkNPEbdHWEmUHLnsbxSW5CimY
goJpqhIuDRNWHwnyj+Bn2H4k2cbm7xVJAt9BOXE8+j+zGOURzZXH0giCQWwvxAeO
ActfCDNRiXmcDTMl6JzrnOy9X9FBdK0BEfJr+hzSQasgBlrPM8uec9xMJy2HPwmP
eR7fPbEjkCpzZmrLsU7drIX0ZFT9poRmSsmFIGHN1hRhSmLpvGjkggXbo8qSgZz6
Tu5EYiFKWVPgwxPsZT5k/qCq4ZrluiyZjcsWckQ50q1PKlqSd2UWhrsbcUBFcx02
wv1N35GBYJUKlv3hCmBp4Jyj2/Yec23WQHEoBT0NERt9K/4AZ0kFIreC+ad2V5Pv
Y6Y39xg6Dmpq+w84vOHrdAe0M9DPyjwVRB5Hq8jUyRvV8cIpzx71XJOQYbZZa6YP
82MBi0eU/PjWV7hIDvQLn387ILyGFSwxIt/7WuKMQWJfXOBwz847RRR2QSn3Ricv
lx3QLUGrQV06xVv3sHKyN7DHHL0GTXtXoiuy6WN1Yq8aSCejDyqH+gkWTap9pvFu
I3kzktWHpeANcrngqHJh0ifjyD6helA6iSlKmseQAw5lxnLLkvWl1SxiJG+213pZ
LY+EWFGxWzTVzq2TpgWwfn4W4ebZvESFXdmvATH5qj2vFzbR40oq+Zghfgh8Fyu/
fRZhGnNYUFH52ImU2WdeyJLfGRqcam6kIEr981sBEYOmIULAlX+472oXogFs2yXX
qmju/L9yBlJMLM040UlG9aDifduHWW0G4azyDLvMLI6VZB8yVysGPGfIA1VqpP8j
zVg02toSZD/ImwtClQQYfkOOiIKuZluGO23Ui7uHNsvg+wNKL794dEWMWdy+fs1R
GWg+YsUuGRd5FdWAXHkFYCxRHEQmRaYrXR32TP3cUHWikkbnwcvcFWAwvj4lX1F1
3qghPmlTaa9pb0X44fIZAr9ZrrjQE6QjcyyMvkw8o4z+4HrLef9/JXw7lQWdnKbh
OvScXrdKzYJWI8P/boVuHabH2oaDfiVBTL5lOWWS2Fudv9iAmTUiEoUSagZC3xlO
n5cSiS+IdfMB2pPfatyNkGJubW686fLEcDi+VO7GaEWXeYD90o+eowGYXIrOGJA1
CpaKozVc1yvD3AAEeBHwYcuz3N/mOzlFwMEt/f1V1bJX4K1/F6GSzRFnWIq0bzrC
LVQZlrLFSVlY4fg1tOR9KmZoWjBBXvJvK3nzEQrvpfLBUt5lkgnqsGPyqQ7Irfr5
ZIvQWB/PsOfP/zgKswur+9eij3o0jaFMugiaK8OGtFfArrBXNT8crLsM2RcxoktS
abdemMowqUVHjnZ7+E9wLds6C/xMUa2HDFIGTdPSdt20OT95Zwo6NGS2eGTtPflv
/fMqPwdIL7IcmXLIRqkAlBWLK21jWsPjfsSXW6KqwjM0XL2UnON4trRO72vwKq65
5mHBsXMYAIjd1vPX5BpzU32cHPJbgsokwz61b0WRrME9ZC0bCmb406IVTU2dItIA
hbL/2hQRujn4QKE0jZzlhols6FmUw2Q62jfE7d0LqM5nbcou3pvS/gVsHurbyckd
byg85K32QxB9T5wuytRJE7NVAmfvzzxDnC0gKU+PPfi3lA2GXpe3eOAhUvnhy5PG
aJ7cOgzTsWJklsgSKqhBYzvZVsSdnAUGwaU9uT8VKtWxO8Zf0BD9yTmIP62ULGUg
SenwR6AKZZDqFZiBSgJcRssta67B4uK+fKwD4/SFG07BR6evfxVCmfKVtbTY2iCN
HVriOFYcWRbz4d1xgdvTOLzBicc8+hPUgJ1IbkWggs5huPXiq2zAd7iVCO6t2RjV
3qgoPZF9L3qFX0dEzW6TaNJN1XODejDcevW672D3Ps/2lFLZ8eD1g1eGNG/LgenW
fEyKB9Efisxyb7FG3/cAMzKztColxJyj7qNcA8Z0reyPN99afKEuwu4q9gdLmsnV
BZ5ce+SDGeufxfo+1adbyeJvC9qsdFTdcvZcGzAI8kwxaV8fnVGtBsl8EnpY288U
zhXvQ6BeSqjsxijONUTVB27ppdJvJB0JvJy0hSDHT5a5fqDm9DKOrVC0k3f7+zB3
1tmNIu7cMth1ZYjlcBCgwVrAslbDDP3OBhNQ0VmSx1d1SFxFFUoQlmu9w9SNc9XK
FJoxa80vc1nZu3mPP6aRZRkFRj2j1hE3TGL22JzseDv7c6rcxtsu+rsccB5JV2Ac
iKweRCC2DDGXjACLAoKes4CIRbmSq6i93Eim/wLQ1Fw0A1jiQAcmiqJI0RMyBKGI
/PJPa0E2zXY4WBmTf9lYBj7I6S45t7DyzDYZfwnk6NrgXoFunfzK3EjJFMtkoynT
e6X1gxDtppvqmbc/Tx/02xcwHE9ACNTniXF2GBLw2lTuYgNWVlAfruhxReT9Nt6G
ezuiwOZHnqjl1mfZU6Kj+/o+mLht33CBQkM04FcDyDUdCFOX/qMvHH/87nkMaxmq
MEzMfaqvaIsKd3agvtcialvsY6sLAQH0XTr1RMGpCxJmlQHYw1OlfB+zrjNeuFN1
bO2VWUfROGZajt0Jhpv7rDoA1m4fuOYZhpKD2jP/Xgznzco9anQhtz4sTxXfjlXC
ey+QjTKGylweyd2bKhS4l+G+F2DMm7Qt/9N+6mf18tbceEMZ3rU1D2nH3414MHQ/
sEITL2rmx/xKDWgwF9ajN4HFV7kKpZxd0fo2fUOVRR7Sn9N47cofhDhn+iieP9US
DE2NLHtjoPOFG0mFjHe6Kh9S6TDlbidfNOXU43/0O7DZiInSaUaM9RjMafQpgdep
KcpTPnXYedXDMtP+0R9ukztgL/xQLRKh1NM7FXSa3VeeW26lNmTwqMuBU//ZVnVf
pKQ/jmSR3+IJpub+pfbpm8VnT3b/FBT53NbOjkZGT6mSUEevtp0LjI5hc8Oygg0Y
EsWbfNq8ERFyM/DeQgi9sNkj2Fco++WS0kTbUvD+m98AAqCK+T9olAmQrx9KXvoL
bq5e6VZVpO0sdlwEcIQ4Rmnm7qBmMdYbIvPbIKBqUiTGFfrsZRCNnIIQFl01vp08
yluIzKS1OLwQdbCydL3gZW8nsk4Gtk5ZdBFD7tnGsab8ibsEfZa0g3EZ3kVFqHCY
gX9kexbso1674ZPaXse423M+BKgzhDKuomOjvb57g3Ms6tZuidmVIucJj0KCgVOR
qaCocg6GDKBZRqmifO7lQ1Q9dOwWQ31lNvxoJkzi9GSLwX/s7wami5icr84iSdFJ
xHCOJCO9Z+Ky8fwe0wiQgds7geFEduEpOcaAS1UunPhJuL9/Pwl9zV4x3BOScl1R
kcFg778Tt6UPVbxE7UJJB6Bh2pE8+4TO9VQTHHArqDi3YNYETV/wndaNQc8V3c1I
dasXaHV6vxWDOD+gZhW3lM+HkrX2Ayj8iNj8fyUbHwizl/5TdveZXFgoAHaWJvtO
QtZb29MUyqa7DwpHbg5qn5uf5A2dTQkzowKHh50lLYcZZ9BTmTjlm2Ohxv7+/Fh+
6VQ7p5Ez97KVBK1Ee8UKziluHiKrEQ4bY4FqIPwpGTBVZPjz8xQuK1sCWBmaRlwk
j0Lnw9W4dXWU2nFPWNrHGoQJwbVAKZgN2F2arPNtQ/t1sXDEJ1L7s65+wFxCiCTt
1EYBkQA0iQXmy+1/hi8ksWn4A6eXnpdXiPwjN9KJIqd8Qwd8n21EzcfNx0OdEZnu
VjBEsRzZBOfQDfJsszKERUelNdjoXb11B9mkpTfwakkTcc3LDH6c6VCa2WxzwD6J
hbDCbMo5mGcPtSg6+10+lf44knEKKr3yRQ+ThTJ7oBeu8URGOzocJpyyy/aEpFZb
O/rTGqiazGAGP1Ord6OoBw+9w/5VfGiyGMO8mr4xIqoqlsznnwK6cLgov8O4iUwu
m0Bl3RwgjcimeyiUmdbUGQFuyhf5OCdFVuxlP5TmTPJT7pCekx7/Xf6usUvraHpA
Y9ZEghxpbbRH+Y3MCGkWWlTgxyDF2t4fOcmFUeWZGfprNPXQbFbGztCroWnLfZlA
4sonLLILVX1zeVbCGJas55TVCheSWI1SVqNe99ytQRi/XyTNe0W6g9Llbd6TlhtM
VXC6DgRr82Dv3eX6UhZ6mBP+vJC1pj8El3Fluz+/TtWjkYmT9iqHfRTtaZqWOJO3
dsQvt/HA9e4Hg5KcmKlQWsmSH5FIspVUBTuOW74FTLTjP94XHk3cJpqUy0rPj5Pk
yzcN3IS62RSM1S0QNdgVtrFuaz50v9ZT1NrS1pGDqhUPDr1ysFpgg9FJza0s4nqj
cARMEAT57oMS4b7eqIcQh/OH0OmIuai9xSd4uLD08ntNWxQBGrAABrXp7CjMHCB8
xRbjCOeSpdtpw9x01OyluW3egPRJi6QS6jxkBXF+22FobhHIZ3ituinL4wjICXqh
H3hlZYBWt8KhYNj7pTcGrS2U4INQSivkwYwiDBZiHFUk1gMQqCoiiwWmnHSJ3hCM
dz3UGAJ+yu4/Bx+CSY9BQoeo99h2ubknwUQedf/wsp2SPmcTU417XtztjEWlv5K2
fiOdL+Zk7axBov7R2qG7ZKyOBKs8O2+1C95HBxDjTCvKXTruOGvwdBBWDP6TnwtY
K+EDJsg3P/cWS3KCyECGt1uFYqH2G1A4Wxa05OWPStT5cVmqKS+wu5GYOKtTUHAT
q/ZqODm+m/aIMwrT9b513GUiT+PmTv+Yi3QTyMI+c4bjpOMHgVkgzbgABlfiJts+
kBF2ajisBI5Rdz377FOJVgB1VmL3ig++bbDmMjNGPnPVTRVWOdhJuiGiT56PDkgv
ww3RTYngMq2ceYaB8JI3a+oo9l53DftVgzO83QWoRnaS5zNerZNXceUmWPz/qEpg
QN+5l+IhqENPMqF6tAJ2KNJtVW/+9d98PjSprsPxNd7fNC3xUwBNY9rvjPf955ln
6MDnt+FVGUmUkENgn6nH9iIMOLA6Va4irE2CeUOlxO6Amg4lFOF+S8iPfqYAg6k4
gaerdwhwE1VhzNXoTWrdzURKwsSjA4/kia6v8atG5jXFsJnZA/l7NzdwF574bZIQ
4FwPcmm/10JOrDvMTeminp2HrY96WdyaWx4jyk9n7iTR9Qt4wOjQIxKrIurNs1tF
ieQP6OK+gPJK2C6O1gSDnTCkIL+11ihx5NtzquH3viP5bH0RjL55hKvZ9X7zRvcT
m/uY8qmGvGo/YN8cXxoUd/5BZQ/vLGxD+gqj1lZUhV51hpHBtmFvd5/+tyY4Gcqr
LbozKj+MQy2oOtXFKKZDXHjt1YC2UgH0PHttci/GFlTqMA+gZgjs7NcCWMxDY9hz
T4Pcpv450DtXF5yr0VSCd1uhfCr+5+1ud3S3QLhuExlw49C8xY1HTjtxcaaUFE02
KSHSNzb8OEO8A5aliwb6r+EWRRp1X1M3pgjF+dv3CL4jEgrhNMwInHW7T7HhwvOP
Cz7PPJnl9ouryBy5J74FpK7Yg0UE7GyOGhLBfv+O1Ipm9DZG2PzyhZgZUDyDE5iZ
zEFVImBU4Ur71hLYlQX6yzYtymX7mmIkDnNjsDvacAKW8y4orOPWIWmjzsz58yBC
ur0u2UI0kvdxjkWzxR39q2utYgW/PqNqQla+IkrhmD4rLJ1zSsljitb+a9H16RDc
O8Uzj7W0P1Zctvp56kcF7dsxJ/yCupOJXORTAKJk64JRqmFRyNKDI6UpqUy1bYG1
STxP8i9PjkGaHnRWx+Nvb8MQ4qf9S+Djowy94wdPZ0XcqIOcJNs/mmi1YEzXDOuc
10S0Q6e5z15pv2eyAMl9Fjm8ACpjou9qODhAtIPmoEXG35jgKNKwYupGgZWfqL1e
3jRjjuopqjtYc7czWh68LreMJxSV65yxAhhvkEZRcdjcqUlYJ+aa0WuQwIg76tuo
zPVRpjtqwmVIEbkpusMP4Chwl4cC3omILjUh3SrpPBm7TaiKS5QIWYSuwO6SvHvU
3xepTYnqE8VsMz94B6AT8A23QfJILcmW1UYool02qlw1xF78KPJvCYkTDFskdnJ0
VgtU54bU6z8alZcaRd86imGTxv4kiiSget/EltZcq8gIAnqljttNCiWpPDx1fAFi
4rccGbgxGXvF4oIpqztaG/ZovKWIR15RDmgtsvgVmq7MCygrhYToWMd7mlRE+L6/
gArTB4itjfvN2JS+bhSyK4HgZLATlUdFJeitlPoD1LlEn60XYUyUu6Cf/POnOtJp
QlQ4SuZ1QdwxUvw5Qqjbn2eUNSI70fqILEXHRcsZnpltlG1NUvXvHJiiDnNuYhDl
Hi3f5I6cU98ahtJFPcEAyGJnZCkjejW4PTyTnvF69ON6WDxIy+Ew/mh74jJInndr
+ilSVpZXPk38mibqat52eJ+NAqYhg8H+IXd6gDn85cUeVpdhM3VGI8E5eosxbPkt
2BPRU1uiSKisBCn+R6c7XcKLIHWyC3oSefiisMZL3E4e/XAMdf0m+gZbB0FCLHIz
IDvBOhPQn7W1glrGLizc+PuXNIwn177DpOTo+eZXeZjWKO8uft4aGECvj+yFM/HZ
LFSa1wN6wRaEF4R/vfOnS/aR+y622dp/o2Q0GRywdXAdaMHaN5CtX6hh2tnVPdAw
p5NW/7wJjormdeaAHRdfpJgSJQeRKxYdBQNYauML4G+YPyRkpzarPWgWpZWVNtP1
264mves72QFFMhkFswOSCcVzgLySwQgNobLlrsoXIxyy1PDcgVyXnG4kZaRLQTYy
4Yt86KkNYgynlQyrDEfh9VDeg4hnBOU5VAw19VOGYuw+I+XOf/BkeOcDE/lW26di
nsZr3/qPu/qzhUp18o0GjA6r48fMaXoIUE/Otnx2fRUUCYMMMe+YNeJPIaeP9y6J
6Mmex1JAOfFtCsnMYZqjErf6KOGvrBjYLjdMvbQ7J1inaVf8/1W53euAr5pkPJdB
N5q5hhV9WIXNeSVJIw266kwC0MlLE3KN1ukHBT9K9U0Yli3tjq5kSVYizKM+k2sa
6RCuhuZeWGY0bUo1WZ3J068P8CaiQkv24DZRBNwDA82QKDfFBRv+ZP1UqkYFKWxd
UA6OwlFrxwj4MJUEiFsEqFDQR/F/zTVNUQu7YgW8aDKZ2Vg2RVvlJOCp0B03FH0f
4SeQV2RJHvVpYdEwJzlYhLYX+YSaMfheGhtVzhRh5lPMImSfFqEkXvZiivx+bnkp
5jqpHeJJMcMgeG6c2RE0c98TRRe7Ppai0pYBxOPNfo/ZoaaJQOgNUTxtyRt2a+hR
ioPJebPuHPjGQG7PIv9CdRR5m9F83yS5sZ9fUQVrDRHko5fQUCgnsneIjFPboeXx
ehivB0U7dtsnpti9TUCtE4ShXcEQYQGvI3ry0unKuKCPWPEznA4asnuyKS1pCsHN
VIofHX46EKeX3kBcoORpcI2U2Kc7gnTsxrYG1NLIlU63YBIC4rceKnEF4H+UwN8j
VRaAmsnWWelCaOGQGCAISRTWKuiamyI/VNgmwGUHJN71XR2KWiIO1C9peL/0NsMg
+wYCJLx54YfpbXrluxU/Oirw/pgLggqL3wnUPJfPyoqw4dl+n2w8E3dQfgzp5Rue
o8d1ORmrP7AmSgNq1sWjl2wxgOE1pqP8S6Y3Q2sNAXO1tdJOQ7JhuQ7OE5TN1Bp2
brZ6R+7oixF4QJlp/Itu8zi4H975HXIpROK+1rtnWExkfh5FcTvskXIWrsOmX8OA
818akOPhEoLjVI0FXHOzKcqQYMoZqwHycd1hiiojcji/CCEmqp2jX2S+XTXYPkDF
HCGDK2OX23o5ks7M4xZ2ZoD6PBYWVHiaWtWGNPOw/kazvXzFkvFlhxT9XNLpwgRR
j3QFHjs83+hZlLJGZtmfcE2c323SkAbi8yoD5/ZIiBrMIpO9qI3SnQ7AeXaog0t6
e9dsYxe8SyjS1y3fa6yto0GyPy5F0xzfH8BCGTvj9LyHpNQa3+lDGVycCJEP+0fM
rajT5hJPuPUff+wfWU/9hwFdOQBSrIGvqtn9hNaomO5ZR+L5wbJqKuMNyDgBZB9X
wJWQRPBxWxclX9Xvkyed/3pOnhPIUUbtULQ7OkchVGynMdOqWodMg57eQ9QzZsy1
wD3fqZsv3XEKdhC0MuHa8iuEIi3jhhaAtSzpJYrBTuPjwHdmDGE8qUit7wLwvh/e
jGTisQUJ0iLkRHuPk9BESbY9v2s++URS89HtKqiFq/qhAMKQsfpfb6qwfYg9/vpx
Q8rM5tCfx1vRALEp/CeUJhb5ZVMqi8Xyrl/a4nGYhNdrNXqVaF016Hk8qzi/VfaA
mxd0MGdDUhAyUYViNbgJEA3ThSMTqgfxYJf2mgp4h7dSM5EO/WXvoG0BZ5G18qby
a1dfJWAKvxC/DMlVFaB66ofcc5jTzhzkml68X35klwuTKb6KHgraeYElJl0t8Xpm
lwXx5PA4R8YiCIPqXbwlsWR7qTUl3qde/vN9k6HTMx1PcZcHeHuOwE/nJhVOO94J
sYYxNzp73qD6SX5qqzrD6BC+4yzb6jDPBp94jSfFH94S7f5T+sphXZUjg28dGRu2
LoH6xXE/pKrt5M2Cyo3kMXha+R7fKl5CS55fD8D3M22a5/9azXrd9s6MDYlqIHnx
5eoQMp8c5Nleqyl5Ki1RFItybleE0tmnSf63UIBP1zqy8n7KlVqyAY3hz7OONfOt
6a2hnP4wvQbymBpGUv2T+qEbzWzh54pcJlx7VrhmtEOkK2EZJAfaHzYO8aW0d+gw
l4+I3QsyCPzElXitx+6rAbBOuPc1ztXGuANxFHzrB1YFFLt520vlfWvjTvJ4ZAaR
b3syVqQcxu5QX3w0Aav5H7sLQjZb+IzshJ7phvlVtqgoqUkjyKMHx6i2f70ba1N8
MWwX+TI113xY+Bvz4F/Bka2jkv56Al4PRaUvp8nR+Sid8Pt0eMan+EhlhV2qkOEN
4pZWRJOzpGmsgYdv58l35poJ/iZJX7jOqqfevT66tMJ9XdAMJY9/gRWdmtwO1wmp
etySUfwkbTJHeKIgXnmaCLtDYmQBuP5lkev2Q7CIHqc+GqAfTAHbOuWd+ZtaMpay
FeRhifNUBSs83meWtvbRKRxwN1dqVowikerXA63jL2VQNq21TUWTaDx/S+OtcFLc
FEUXSSr/x6HT+rJ0dexEm9dZfVSuWmUja6iYUu0Rpmr+/QlRupJBWdUzC+tWmea/
MAZAa/QBdTrlRMg4xi004yEsd8qBzy/27TyawVntxXiRp+23GkJab3jRnL5ZZ6fV
GSeBBN/ROmJSgWuAKPOlb7dofHbQou4ukjh2ypbITJwPjDggYrsWrFx/I1a+yQLf
Q6mWs6mjJDz2c+QoWUIYvHCaoiv2yg6Gi6qXsPu5F7sY7U8nWHJfbKfDJCbXldLr
01hrPbIOfrs4J4DwsuqtROE/d2OjcrWt/JbiEJ+3dBZsnbeF3OvkJUuzbIqbo23I
HZ1F8FmiPtA8x97UpyTnE2+FXcJlgdlnlPVvQ9JLGZcSOrNofzH5VLXsL3knjUVp
DGYqjQ/77auSKO5VymZ0ulSzncluBybgdgBIJlAeKpQKpuerCQqOGfe2idmgzcLM
D8J2CUwgHof9tLWl6r0Bj9pWell3IqxygK5ZhZc+w1w+PlRyC4t9uJAv+KF8hf/B
A68fCLXS03jdeBoZEEcl6aHJWfTq+c3YV2/mxZDfsKSO+DioAV4elxj50CTnOmfp
Jvw2zrBuqnPfZmONnEXumRC0Gdo/jNq1LPM7vmTmud4M1yI/O5XZiOAIqpZwVjyR
L2U0EcUtZdVsuQS2pwW2RqwXn5JRLex56VZYS/zsrGQQ2ntTgyRJsQss7cbkrQ3u
vqoAJ7HWA3crOXSw3j44UmOD3UF/PyBcj2y+E/oBgGhqqDHVqLDNzA+z7y/nx8/Y
RGputgNtqt/DTU1hk/JVEK/HK9TQikCko71utUxDHbJbv71PCDJYPNMXQpeFd/q7
jIklZhxK4Bh76LYMNbxEQB8DXTA4h9vrnLU3Gho3Oxa9+OL4ggsCUgCmcwVws2fv
9ZMv1AuLhicmMKxSRePef+eVv2O860eIEilrWA86vAxVrK7WJIYIpusK8k30FM7m
NNR/cgHi+Tm4yA6odApmMP1sMdtzTLhZNXJJhs35E83DoENrUZSU0WE3ZyLHXb1s
9sxSCUlZynEG192JyRHO35c/UkXCNcmGV5GXMg6LIYeVlkvzWhbNMKcdoDdukZeH
+AY8Ewv7izmqwT21liTkeMi8bx9HROQHYMDN9i8jJ+MUHQog9j9iTz0QDUvBhD/m
sWt8ljyr2vUf53zB0BQLxmgRAImWUdkVdS9m+s9yytxJ9rLaftILUhDH9y4O2vme
bm7ekeBCrEgHcorTm/8uTs26I3uMDyot7bZxTDVlZlRb4dpoqAlQLRFYiWcz+Jwo
gda6DawuIvNuFyMGh05A7ys/ksF+IwmsGvEXbv5vo2P96lzGICnieXO83/47IRfe
+P4b090qKPR888KfGS/Nk3rdKIRcoaV1NgJ9CYvffyYihP7Lir5mS2LL9WgIeQxH
g6vLKMqI1VpY83DBqxCTrURMdKnWPJS9iw5zSz4Gf2g5uvHH99bdjlVrA1PBFNvb
tiPH5ZRYUBvDJJoaOIchChgZ8tLwThlJ2dWXKwlZ/0BqCbrx80Mm3bc3H1Fl7yif
7w4EGkosFUsBQbT9oOVeFXY98HXM7bMn3SqQgac3pag1TqVIFLRr3VQHgPDV6i7/
zQKoDWMtRVigm5YNumM8EALDgfO/A+A8BBgvqxpjm4fSZWl/b1TO24zgbcUwRtaB
VteeCCIMLHp3Bg/tDIS5MdTvZRt9bIzJEm0wXGcAQIDpsFlSQILKRT4Ee5NUzbmR
xFb7zPlqobQGI0FwQM72g1QyjOa9Ilr75+ZGBQpHDyqIh08JSSo9YbtF2QsthefQ
oIWSO1wffg5w88eUzaURtqJHdgS4YeGB/SWC/FFhtFcHUftBNYqnCRlYcziWDZsW
F4pc3I3lrrVhDKwugHLlHB98w+fUtibjZkadTIWntYX1dKimva5uwirfDHYblCrb
GJEBujUX9da05FETvm1T76cUASJDwjoK8j7MKnzFN8WV3YUsyJIJ3KsHIu1rdpC3
y14IIAoAOWCq+llELdEYDzltWoYrrihs4an9hSWkk7SSEdI7mYyV9kFwKw+ycCSN
wOTmiKCFrhLEzx0pYMYLt20sCb/hBob6y48AoGGVLrMZ/IaVMd8zSi9dExm9/84C
7bKHWDCIr351d7soXlIPKQDTn380mGLFIV3qBSA9RLSze7vwQnQm1+cvKD+ICjGz
2Ch8k5OGK/WlCSnKxfSj+kqIJOi+6l0HjNuNIcdIbSLbWmseicFf5NIvs1BfDHsp
7Iy2ReAFRYwxqsPghWHSDH3XMAcEA8qK0uFAtirmm75Kvo7qhpOgEQT+R3KUNqbz
lku4olHYtmDwg3TNYYvBydRe8bZFd3tlXIxyVmTYDvrCyVwjuYBFj2DdgIrWMrEZ
6jYm+VDmM30mgekl+pPHfDIh6qAS2ZsYfD/Bpv8v0iXRGBrsDhr3gCu2Lf0z1Dax
MeJ7KsffYGGnzylvkPvwRFqeQML98gqKsimW9hONg7AOjQHOcCoyJhf/t0wB7HbT
6j/0sjRgc6CIf3r51rGgMKnUCACjk44ub/wfBHz1oQ2aCxR2RBoSf4lG+e1OXM4J
ZsxMvfjr4bLr7dug/qnCJmJQjWxVRpF8NX6+uk1dl6Ll5lhLMx9Srbz1G0uPuj3c
`protect end_protected