netcdf YORI_VNPCLDPROP.A2014033.0000.000.2018274194737 {
dimensions:
	nx = 145 ;
	ny = 2 ;
variables:
	float Latitude(ny, nx) ;
	float Longitude(ny, nx) ;
	float Cloud_Optical_Thickness(ny, nx) ;
		Cloud_Optical_Thickness:_FillValue = -9999.f ;
	float Cloud_Effective_Radius(ny, nx) ;
		Cloud_Effective_Radius:_FillValue = -9999.f ;
	float Cloud_Top_Height(ny, nx) ;
		Cloud_Top_Height:_FillValue = -9999.f ;

	short Mask_Liquid_Water_Phase_Clouds(ny, nx) ;
	short Mask_Ice_Phase_Clouds(ny, nx) ;
	short Mask_Day(ny, nx) ;
	short Mask_Night(ny, nx) ;

// global attributes:
		string :time_coverage_start = "2014-02-02T00:00:00Z" ;

data:
	Latitude =
        58.2, 58.18715, 58.17426, 58.16127, 58.14824, 58.13515, 58.12197,
        58.10873, 58.09542, 58.08204, 58.0686, 58.05508, 58.0415, 58.02786,
        58.01413, 58.00034, 57.98645, 57.97253, 57.95851, 57.94441, 57.93025,
        57.91598, 57.90166, 57.88727, 57.8728, 57.85823, 57.84359, 57.8289,
        57.8141, 57.79922, 57.78425, 57.7692, 57.75407, 57.73885, 57.72355,
        57.70815, 57.69268, 57.67711, 57.66147, 57.6457, 57.62987, 57.61394,
        57.5979, 57.58178, 57.56554, 57.54926, 57.53284, 57.51633, 57.49973,
        57.48301, 57.46619, 57.44928, 57.43225, 57.41516, 57.39792, 57.38059,
        57.36313, 57.34558, 57.3279, 57.31013, 57.29225, 57.27425, 57.25613,
        57.23789, 57.21954, 57.20106, 57.18246, 57.16376, 57.14492, 57.12593,
        57.10683, 57.08762, 57.06826, 57.04877, 57.02915, 57.0094, 56.98952,
        56.96949, 56.94932, 56.929, 56.90854, 56.88795, 56.8672, 56.84632,
        56.82529, 56.80408, 56.78274, 56.76123, 56.73958, 56.71775, 56.69577,
        56.67362, 56.65132, 56.62882, 56.60617, 56.58336, 56.56036, 56.53717,
        56.51382, 56.49028, 56.46656, 56.44264, 56.41854, 56.39425, 56.36975,
        56.34508, 56.32018, 56.29509, 56.26978, 56.24427, 56.2205, 56.19859,
        56.17038, 56.14112, 56.11512, 56.092, 56.06533, 56.0322, 56.00462,
        55.9768, 55.94874, 55.92044, 55.89189, 55.86304, 55.83395, 55.80463,
        55.77501, 55.74509, 55.71491, 55.68441, 55.65364, 55.62259, 55.59121,
        55.55954, 55.52789, 55.49657, 55.46488, 55.43129, 55.39862, 55.36501,
        55.33157, 55.29919, 55.26945, 55.2412, 55.20166 ;
	Longitude =
        168.7603, 168.7203, 168.6802, 168.64, 168.5997, 168.5592, 168.5185,
        168.4778, 168.4369, 168.3958, 168.3546, 168.3133, 168.2719, 168.2302,
        168.1884, 168.1465, 168.1045, 168.0623, 168.0199, 167.9774, 167.9347,
        167.8919, 167.849, 167.8059, 167.7626, 167.7192, 167.6756, 167.6318,
        167.5879, 167.5438, 167.4995, 167.4551, 167.4105, 167.3658, 167.3208,
        167.2758, 167.2305, 167.1851, 167.1395, 167.0936, 167.0477, 167.0015,
        166.9551, 166.9086, 166.8619, 166.815, 166.7679, 166.7206, 166.6731,
        166.6254, 166.5776, 166.5295, 166.4813, 166.4328, 166.3842, 166.3353,
        166.2862, 166.2369, 166.1874, 166.1377, 166.0878, 166.0376, 165.9872,
        165.9367, 165.8859, 165.8348, 165.7836, 165.7321, 165.6804, 165.6284,
        165.5763, 165.5238, 165.4711, 165.4182, 165.365, 165.3116, 165.258,
        165.204, 165.1498, 165.0954, 165.0407, 164.9857, 164.9305, 164.875,
        164.8192, 164.7632, 164.7069, 164.6503, 164.5934, 164.5362, 164.4787,
        164.421, 164.3629, 164.3046, 164.2459, 164.1869, 164.1276, 164.068,
        164.0081, 163.9478, 163.8873, 163.8264, 163.7652, 163.7036, 163.6417,
        163.5795, 163.5168, 163.4539, 163.3906, 163.3317, 163.2777, 163.2081,
        163.1362, 163.0725, 163.0161, 162.9511, 162.8705, 162.8036, 162.7364,
        162.6688, 162.6008, 162.5324, 162.4635, 162.3941, 162.3244, 162.2542,
        162.1836, 162.1125, 162.0408, 161.9688, 161.8963, 161.8232, 161.7497,
        161.6765, 161.6042, 161.5313, 161.4542, 161.3795, 161.3029, 161.2269,
        161.1536, 161.0865, 161.0229, 160.9341, 160.8566 ;
	Cloud_Optical_Thickness =
        8.62, 9.86, 10.59, 11.24, 150, 15.9, 16.34, 17.44, 18.18, 150, 38.5, 150,
        47.47, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, _, _, _, _, _,
        _, _, 71.39, 29.03, _, 29.83, 22.72, 18.12, 18.08, 20.18, 33.37, _,
        18.76, 29.29, 19.94, 34.02, _, _, _, 17.56, 19.39, 42.45, _, 22.68,
        22.24, _, 20.54, _, _, 28.59, _, _, _, 38.47, 25.09, 22.05, _, _, 29.4,
        _, 23.36, 28.13, 20.84, 25.15, _, 33.34, 36.44, 27.32, 45.52, 33.91,
        30.69, 28.7, 17.71, 24.16, 17.06, 18.73, 12.37, 16.53, 17.32, 10.21, _,
        9.72, _, 2.21, 3.47, 4.47, 6.67, 8.8, 9.14, 9.51, 9.77, 9.28, 76.02,
        53.88, 39.17, 6.32, 8.23, 11.15, 11.4, 15.01, 16.83, 14.73, 16.31, 13.3,
        10.21, 15.79, 16.58, 19.82, 13.83, 14.4, _, _, _, _, _, 11.14, 150, 150,
        150, 77.99, 38.24, 17.73, _, 9.4, 16.57, 41.24, 56.43, 23.27, 16.37,
        15.93, 28.09, 25.51, 37.43, 14.05, 12.85, _, 19.4 ;
    Cloud_Effective_Radius =
        16.14, 15.58, 19.68, 22.81, 24.05, 22.59, 23.01, 15.92, 9.29, 5.5, _, _,
        _, _, _, _, _, 4.26, 6.2, _, 4.96, 6.55, 6.6, 7.01, 7.04, 5.23, _, 4.76,
        5.78, 6.18, 6.51, _, _, _, 4.02, 4.94, 5.39, _, 5.66, 6.36, _, 5.6, _, _,
        5.44, _, _, _, 4.02, 6.13, 4.22, _, _, 5.43, _, 4.82, 5.83, 5.64, 6.12,
        _, 7.4, 6.79, 11.09, 7.06, 9.86, 10.59, 11.43, 12.7, 10.28, 15.76, 16.2,
        21.93, 11.58, 12.67, 16.17, _, 12.52, _, 45.9, 46.95, 41.41, 34.32,
        31.01, 31.86, 28.67, 26.78, 26.07, 6.08, 6.52, 7.23, 32.03, 30.25, 24.88,
        27.83, 25.41, 25.47, 31.13, 31.07, 37.6, 49.18, 34.19, 35.59, 30.86,
        42.68, 36.2, _, _, _, _, _, 44.88, 4.03, 4.28, 6.5, 7.82, 8.24, 10.45, _,
        25.05, 14.66, 6.52, 4.39, 8.12, 10.79, 10.26, 7.87, 7.35, 8.07, 14.95,
        14.7, _, 13.02, 7.42, 11.84, 55.1, 10.32, 10.37, 11.34, 11.25, 9.45,
        10.95, _, _, _, _ ;
	Cloud_Top_Height =
        2791, 2762, 2832, 2841, 2970, 2948, 2860, 2805, 2791, 2566, 2779, 2786,
        2939, 3072, 2910, 2914, 3742, 5057, 3901, 3372, 4072, 3040, 2782, 2853,
        3197, 2840, 2893, 2855, 3002, 2786, 2436, 2870, 3085, 2938, 3105, 3246,
        3187, 3180, 3198, 3289, 3217, 3228, 3063, 2936, 2853, 2877, 2978, 3095,
        3250, 3153, 3018, 3429, 3447, 3334, 1888, 2042, 2205, 2304, 7451, 7399,
        7001, 7038, 7051, 7092, 7234, 7233, 6231, 5760, 5422, 6723, 7362, 7339,
        7172, 7163, 7199, 7596, 7600, 7604, 8044, 8021, 8138, 8198, 8174, 8149,
        8076, 7306, 8224, 8222, 4638, 5013, 5230, 5151, 4742, 2370, 2099, 1945,
        7143, 1944, 2495, 5935, 5863, 5628, 5404, 5205, 4316, 2047, 1907, 1872,
        2106, 2326, 2628, 4185, 4226, 6394, 4945, 4866, 4612, 4811, 4604, 4881,
        4569, 6378, 6369, 6808, 4674, 4428, 4727, 6315, 6357, 6289, 6316, 6391,
        6299, 6351, 6745, 6768, 6776, 6779, 6708, 6712, 6894, 6884, 6847, 6880,
        6877 ;
	Mask_Liquid_Water_Phase_Clouds =
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
	Mask_Ice_Phase_Clouds =
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;
 	Mask_Day =
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
        1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
		1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;
	Mask_Night =
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

}
