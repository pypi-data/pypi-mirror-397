`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
ESp8jRyPtsiY+Gb1bQiTIEv2DNBtVHPanFyrcSALM2m+T4bIiXw+0XcVKqJJtWAs
HqaHdjOUxOo99tpQyJWb0/R/MBCt+eWLa4fzUvis89UpGRQTTcb3wpq0IzlCvYXQ
YeB0kmPVj+cdtOH+8w3k1tGEQ8elc2wJnlQJigWmI0VTs5pjr/RCJG30jniK9uFI
ARuzAC/d5LO6v/qFSrI039vT7L0pxGuhYgxAFqckqjVLvIUPpbCbZR00nleVKMDe
LZiUCYgSVJcIwX5iTTh+lpIlh54mZ7g45qeAR2GLcjcr35i7+3KLdrBhPYcE47+9
b0aRvbHU6MWvYESnJ6gW6VPPovaLenHiNYX90Py13ckbst06ngVj7yIDw3AfrFv/
x4o3HHe8k5RAvyCV0l1D0Ap4yRZkMK1VXeli5PKkZfaSzfbu68C5Mf2NP+9up+2c
T5s3vZXYcnShx3UBcc3iJJHBBspyFzFfLr8PGOMeNh5Rf0SZRNPCbGI+ZmnxOFaA
m88O7LN+dDE24/6EW8IgEMUy7Cz2Ea+ONLqOzZz3tlSUTqxThh0W3/kC7gXPs+20
IhZVCypsrEusU8s3wfqv2kBDZ7zTuN+5AbIOvoRvopaeqqpEwpLHBYx2eNQ2F2Mo
jRlLBTsuxknV0GrqYhVJAFHUqefOCE3igMt7mVGw8yXvdpK3sf7y+/kojFb9ux0L
QS+aZ3Gpr3vmzk074iUZHY0pORBgpUp7D9e/mLNkcria9donjYgOz5skI3b+tVg2
kyNXbA5KHG59AtXcvfjhfa/2ZiNN5DbqFi1TvzZkIp73CmD6HxJzJQcw2nknuGKn
kYrgBAa8sJe/KTcRw1B/wAYaWN5nu1hwKjJGMW+raSLZWtHfeIuvZP4AaHnrGpU8
YxC91biFZcr70nfjVp7MUEuGCQo0Lir/ttVMzWoQT3i7ZghAes9sd9wDAjxuc4QS
3Q7PUMRerECs5YLspNCEAvBia8any3TOBQfVvgIfWNOQ4PhpNqsO+cOxeJ+NIJF6
7ab2QF4lhv79+2jIWJlUvOZqT6HDu3I0n4PwUSzWThyaG9keZqFO1oDNVooSIbXl
DKprEM6OleJ1I1ZsI+hfMi/J558mtY/ZXtiVDMg5CnetuljyuA4LXUzjTpvT/6Ht
0/60DFXmD66EDF8pLbTbOaiiAeNc32RsEJ75hxpd611GROmmPts63jOelmdX+89S
uqwLi++mTp8otuZhKdqC5BQKZNEkWoNmMwWM2AcBPUOxXOThBarkPCGXKPUrakPX
TGQNx/7jimJIuYqEbW/RUl4QA5I1Y39cy52byqLTED2GvbcdTfk7VoCfhKAKsIjf
ET3Bpr4QgtOuS1jBIytIve0URQTZziMarhZ5KO+FPjCA+S6SZbB2SaKV1E9vQwOL
WOfcpBDoum9O/ENHFujELd7SnlGTkLoco28tFqHkCxtWQvS7TfemZduTNxbOg+NW
Vr3lihTdV4VJK1s9w5tz1/HdG4ZKKgERImUqDKt9C+LAq7jTgAn0jfujUOwk8SUC
wGjobZIgWHKN9KjQCbLUQF6Zh2NXb3OuW6BikSzSr6ZuOpQHeJzAwUG7MI/0trz0
B3DFaaKtBxug0K+25GoUi4Q3LImkjA2fKJKE/EJS08Rx48yxHlMrwzyf51pe9tHR
d3+APH1BhKclbOWHYJCB9HNFXKMCYw1lbiO9sUMUi/SsfdYyCjhzIg1XU7ULLl7k
sDC5MO2rurcdfv/xXmDV9CC4Cu4t10/oiaJEV7S0Hzo6bOIVLT0BEx5sxj9eEaOt
ckmsxPj6X5Exkmpyr7r6wQItTvtZg0Yew94T2W3nupB5uZSq4Gu2vnA2gshRb99M
KSmccBb5dxgAkfHyCG5TiM72pKw/tBDtILAfftz2IR5oJPpuhv9x7PT06bJKkR5h
q9JDoR3Ofvc7Qgdcr+ZpYrt6/9H1wBcVOIugA5zQAT4v+mnABtWcP3PwK3yeBogi
aUg+7hdk/wKBZHrmqRq9gv4J6XbMu0pPfhd232yjBI6Jz98Kfa/QCd99SMUm6j5T
eKWHRjyz6BTxPEGOE9aWSBHu1SJxF6xUafHE3YeY1wxdPAFwrpDGPKtU7Dt7/QSx
orZtjuPwCp6rnguRe0d+Z892Xwseu0Fwmz4nZG4jcCXldEUZ7pu97tL8G0GN4ocK
+EOayFjX5Ql3xLmXOQrccKQwSKGKZrUkJSmMaM89X3GytO+UfRbL63uanWkJpWtj
2HXKiusLwTZmngplGYNxXKrJ9pgo4UgvdVc7IjSpauXycJsEXIGc77aBHdhhP7Wd
ck0ouQ3mfkxVoGGGeai9YHusV/tOG7b1Wnk5lfV7QcHaxnABxtyG9x52shuAiSNS
yMezjvAe63w8HORQy4OmCSM+MCXrWpCdxIbKnUKSj7G0MYGN1dvShSMuQc6y33Il
Ii46H+Gm/cSxmxHpyXgr6Msuxiy3A8wOjZLob4C+ltvnRRzLlTXUsW/0SEJoz+GS
Y/Fp+6PMdIo4vcqmYYCoHqJfqxy/XFUQkKaXZjcd7JRCzkJt8qWsHxIlyU3hEtrY
eGrPEA3JTc7qMZO/Cqz//ImNXkhdQi+J++MLuUofoR5tB7ea/1PUgJClBA/KS8qp
VM9s0CeNMaTNvETtuvg6K/GaOr8lDITaYjpGV2T8wCUPXGofGPAI48Fxrhso2ApU
GvigN8RIyi4Rn2vfqhRxTvkqzrlv+EYZC0EdiLHZthzkJ/VWP5QguigmW9opIzp5
G9sH2S56h1HnrwcF3J+hAea9G8Bx7+FantuFZu8zYD9vZXSFNaKpk3hRy+2mMIRT
ClsHHjAaQY+74IzqXX3F6ZxraNA9B19wJ8M6Z09qhKC0frzccrC/x7ptYDZcdVgT
3cW0JUxVGFhNwK8iqzj2n39S08wtgqtiTrW74UTn1FIY1sPajj4/Mtb0jjFrjDBr
du0apFY+QPxiidHvbAM5l0ba52Ud3kmuiqoKRoSvV/WW1LDYuluzj6KPnL6TlgZr
OX/wkomt9ky2n4uuSiemL575x5O8bKlt7ReLSdSXYmrJth67LDZoXadMVKIQ+4nU
DAvCiqbIhh1e0OyuxZu8FYF18UXKO6114mwsjudWVuU+WjIred97lcD772uNjwsT
JrW2E7jtIEBihtVH0Wj3M2xdc+IgJ0T8P28z2AlFOLRG2T/u0apL/AVAwIu+nXUP
XRLaEYfyxSZfFcVnvf7E/n8hhgtXBrQnKeiDJ/qIIQ7etR2r3L3HMskXKWQ8zsx7
LExRipDzUSaKx8sEBVIUIHUFKeHpqHhxH2Yq+7HMhMG66Uq30GCB79bKKPE55I8O
hvjAOiigpt0NY4bL1djg5ChxaTmSAn78INOZxZmfnAWriGMvbn1wJu9al8yo5ldk
k7u/eazcTtMDroLU3Ps2fFhT6nSesxiBgcIY68mTdSwnt/GakKSMetLHMLk6eXid
bgD+T12ew4SXaiuYw3sVLfGUhPV18WFHTeXzeo7MHpwRtmUr0GrwgmgWeV5WT3ey
FAJ1rIfSxtk8mZbu/c/jkIH1c7RkGVqVdKHAWkEM6hMNClZVCHl6CdJiARsCu33N
XYLpwa6yzUgEzhRkmQhXzGPVzMkRqNZWpeAXKJPtTJYSX7uU36W0X9zmlGffmjuz
cIb21J9uqqqTjolq02LQ8x9BZ7I3cekQiKnkHi2cJfsQVQWga6HH5SS6dNyLncxM
ubelLjV32Qjj6tgMXfVcGLJ1cA8hAcby/bTzM8XC06u8rG0+l7uY0QNUm6DWIX9k
TBJrZDTGbgFMBcGlckBIqPkSnYSETIjCKPZqdSFaY7vVh7vErM7mLfVB7uTzn+Of
gQy+5Tm2XgJjTJHOA76Ib4+UpoWvT8hElsUyDXiFbpK7WcGMvxlRv+UWSLsIUmj5
YNCuYOntQTxxdVipwQyf8gvhZDPhI+S1+kvm6NLggpAeIBmqSOHgy0BXSdqnTmT2
91tvmnlAvbSc2crZB4Ip8qUw3IzgzTzWme4xTHAvNo8Vi09ultl/VGnhnFRSPvPi
H6g/MURAVQBHcOQeL2NLjIb87CEkjmreb6JJEiL36ILuExD5ef6uLq4kUu0dCV8Q
mxlts5LUmkkeLm7uDNIW0TqMF9MP6BOZnCi8N2OrMBaF1WCzGefFbj9sARoi/0xb
yJnB5RgU+QWdAm0b2J3my/iQ2/cM0mhhrnLU11Td8ZE/SwiCyzxxFlGH8kPTueng
VyhvwJpy6PvtknVkRJ/gbuigEZxlI08Sc9FYvFdA19xp57wh7IdAcTftlQq/aOAE
1Gktbx0hq02/+fEm5Z1xzptkzb2mVwKxcEM5mjHqr3WkA/xojO+2IVZbpglhISM2
ObYxnXgwL+1+DXAawifvUCYK8W8zCzWvRdMQ1gb/95u6MzeEu+inqC8Neyoq3cGH
2+4pxT/Q8VbzkD0cnV6XZLXIYcTJNYBVicvbo/7pa8sFseObfwo9VyTmdQBBm1DN
3i6JghezlgQgUH8PQuJ0bIlD8rTxLidMxz50oe4YuLQ8n2L8x4fFhe+Pwx1ZzJZR
+/kqAfMtdc7EjktGRETCxzsABoU+c9AIqaoRUeuiLZeV0O8j5CUWym2G6mW4l/9G
LYN61kbrpAnRst2p2cXdInEoeZIfb79J1y1HvA4FgtL32HBrAq6OnhhDxZedCyZV
TFvEPTRFyIBYgYdAW/DTPumh2EO+6cDky0Fv876nDrGapka872SrovfCFi3SJqzh
BwSgG1f/cE/8/tBAcCd88frbODMP/LNVz48+U74Y6JsJxJ2oIMN+VjjHUEsJKslx
rffgHgVnHlkmZxcuy1LHT5wC4AscETrZKVtN6YWFJk4vXgku9LYMlS3lEy0GtO6T
sblnpdEjDVZbJ67817hSA9z5ZEEwOlWedbXMaUEk+VCxlOEaqJmGikQc+qYpnTmc
Rqz0s/g1uKlE6eWvWw0Uvlep8+yG67gnhznI3jlqtFGH/mZmRH2fJbBgQGt8G56k
wqH7dyzWruy5FIwLC58Y9tF17mgLrln4aiB8M7Eq1fFzPdM7P5fmmKlkEEbztDIq
ONHPqRP8HG8oV8vPQ/mS6uisyyKWyL19nJe0AozIY50Rir212PEZ8SF7zJR//fsd
7Ji9xWPvGbr+t4q94POX1kijuqdHCG2IYVGFBaFxSFUkvarx07h4kALufWIqi1UR
UI/a4lfdmCvrSqGnyJeNsKCG1sbZ2yGm4Cx7dOyL1KPu6AHRSgm+JLFTCZxDMSL+
GyUW902b3AZOlFYw3O6MAjtPfhyjsF782SaTcV2YnS4EJ31ZjkljsbfsLfK1DVPR
0sHv/5zAXoNjbc3mMMZvasUnoZ1+YFyyy98urvFxY57Qezckti1ZqaajhCCWP7hK
RW3/yyYkrnDHNpcAsUv+MRFpRcPAXgh9DkdOCp17YjBo9PKoHsM7x5rcKdWaW7lF
taAoR7E0j3bHN1J4cKtZ4oZlSURBU48gik5SIyXGB3t8/WDSMesTNxWBhtNUoXE3
BO6M28QOtJUm9jn0Rko2SWuf7Ht/1G9XSoldl6DelzIGMt36r4irvpLxwhgrDLtw
NnVWYiqY2KM1Aw9s3R+VL5/g17C7hqP2LMOVxEHwVkoxlkFS29iweoH98b/dRxLN
ZoZMzWnZP/zxT1GEUQswRD5Tk34w/dJuWHdhFlw7YDBUKY1pJSoyLiqewMWRC1vV
OEOUCFhSlvt/k6Qe5aga9uRw/GOxTlsv9N0YB8srP0zopqGnKngjLqKgZfxMOIQx
xQpf3X6s33tYO2nDF6H0XnUyjRHAE6YOsVqx2tpvp7nvCaKA47Yq8BB9VO6BU5Bj
uYjxv+sC8uizlj2Vpt5rHUSlyltQ0ks+q+kMkgI7qCsRc6DMVzzKi8UGOMeY83nO
Yt1wvIH8B8rgL67DxUWnPLcBwUC3ICD3ddgDwZur95DLibXEEBdxF3IGnLDdrmrn
VrDMAEbSt7Gd5vljbGbFpyGk83tZt0tKP960wv3Ra+Xij4gtRTpqFzwOrfVsVQIa
kkZP6RRLUeuYz3TkWTB0DGBtOcM1SPzc59SPE2Cb2PaPmUfvf9W4OJyz+8WDVBFc
3fVKE/R68EEVzF6xzj09l3BoxXLjpKyfnmaTOW48T9lVkfAxTwAvbLAMF1uR7thR
n3cXHIOSPigbC2rQzNbnQCT9uZuCMt6efrLW6cPXqSCssEk75lI8OU0SdMXA1aJW
Q2YrKYp10me9Q7iN0X5qDYKJkazT8Rkmqnil1VRhhCCPXAhGbh/kxoQxK/ConF78
h7kd4GUSgF1RugWr5yPBbEAOM/eruJ0q7/6ylR8mXsD6TCiSaaU/OSaNYdO9eSom
BMDW3DaU7GCUKVx6F5yNXMuF3HIOBwX8KZ1ke+8tJjjJdIkQEWBvtA5AmQvZvA2F
zGF8tCag2dDAarpQActVBUKZhmA3Gx3Q5xLbyvKNL7178kTw0DF0TjNBHbgE0q96
MXSEGickhn+IDMKXa4VQbfG43umFO6LFFX3eTH9EyfjVqMgmUYba4F9/Z1P3q6J0
+SlX8GbXfgeApvTKfdBqTe8kvyYuyqpmlYajuAL7+L+ec9tp+Z9hE8CFn3Yz2ybC
SJ6ImlEpLyVhqzujY12K9PqODiMp/kMKxkB2Pfe+OvBQ58cSUWLPag5vtzH1h5qU
g9jaQdjDMWqfmm3Zg4c8zzXPiXg9fdodxyx2hwUK44Y+BhOqDHg6uShFIOHdxl9R
f812dCGIOYGKJ4syEaQANB5gSBSOSMhGaWcER90onasm5OeUAEQjHnvgnOX7vy+p
OELDSPlxjKDWgFk64CZkfsA+yzClJ47YYaWv61EJBVAXDUEMaZPCxEZCaPrXPkSd
c5ETmZhKfUIiyewXDUl46aBCH+VY9AL97UN6M04T1fhB9yCOun26XSzJXbFJuqXt
gyj48kBqLIjmmbIzFdB/AEtRWa6VMfBpmVWi/nxk5PfpvEmlZfvIG/cvoeH8TnKF
7Oo278eRx0c8SgtAOZy8BsGiUMbx6PvYViQqdNgi5lCxQ+Tpbx4EC+iuBLAkob1T
oV/InzLiv68K9KSLkRpj3bvt6h3QUSPXEknFA1Xj0l6LOFDaWRcEHqN+L9YuLlTR
hCzh64Y3aP4RKRWbkPGyWDklYSXbTkQUWOwCCYTJ52o7gjB8u3WfEm6qer2SFuqo
PQ93KR78Xj4131k6CVAwwLZOj3+HgmMHATJj9EWavKzMOaXyacOzRXpLl95Z7d5h
wiDJGpf5iOziKdVyAGmHduRb9SiJf8p2qgeElkbKny24n9ofsAgR0FXjD5nYFei9
lxJwrOIMOwUmvpbUZIYM+8LxpRHaSrNUP9niHc2aVotz3byL6CFGT5i1eKRDI0g6
VHRrwdJZDqZegtIpqTwtUjm5Ms/+XTg0qiouOl0vTNbUrvu3i1WxeTyYgxTDa8kV
VBHvBXTDhkE0/J64/E1ZO+qvwY5DtTysNiF+5ue7W3kMoAaoMxlLDOAV2xxkwmQq
C3mMoiMi9gQhVIEPUQ1qAIij6JPS3NiVcn70QBwyPJzUOTJ0I0g1AFEGT6ymehr/
LL8mTeEErDXmuCBnyWeDP/ZG1cPh3kdI4dhtjT7A48fIjy/5KRirBWVo712vKG0U
HGA0mNCNoMPX1cYw8kKK7l91YonyNQV9ZC7vM93XdK55nZ0WDcT8GJH1wayF+1ZK
5Up0L3qKf9sCA4JD7kuoAk/G6mD8ZFcBr87QpvMuWRHkEB8WaI1rSni8FEKIlttO
goKHxo8gVaMEQow8eAr/tFA5uIAGq0f67hBowQq5NbEl2YVoFA+JZQvfEKuDTaDs
rRtPP1zFZBPrayFrVGzV/GqjuALvvnQRq0aBwbeXoNmPUG7rp67+AGIv7cq6uj6s
nyyymoiXlKSbi/qTXeoRFzA/hvgjYDetCA2YF7yiEBmoOVsldK6+x27ul6L6+jgx
fVm62blC6SLQNfgushvEBo32poSQDb2SJ3V3yuZzI4f/KiD/5zlBD6WqtYc5d+Yz
b5dv+B6ReDhKF/KixvJmEXNdIkYXZBZy023BWDNDNPNqaOXClTnw2y/I/0G4G8hK
x50Rpfga0Fptqm/BiZj+V0wr3sjhvuRrD/ltanoVSguB+nrAKSEbUD9Y58a0R+iv
n4fEmOh3eGtB4dmq5v3EMtn5Q5un3dtB8ychWIM1d7m6Qc80xWmvKqlmKYtf2zM2
vXn2RNhQ0oMHQGFkiYl/p/CjGJsKXfD4S7FB1dqkHDhsYmi7VY1HAP+5x9vuzTbu
`protect end_protected