`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
FzxwnjNthnS6kXdUdDdulLLNN1NMZVX/DcMBpD7PlY+gnfZ4wC9K21qAFJKAcqBq
PJIYdNU4f7x4tz/k03IVCMneY/N3Wzwe7JQ5f4m6Bx7Kqsq9+XW29h2FCUpmjkNv
j+jUhrLLwNsrOgiMQc63HcsmNiJ8Ab1GKhsRxPk8Tr04NvzkwhO+B16iZqLNKuie
MVqao2h0Kmjryp9p6gO3BnbKWFpjWHcRtUn4EQlOYY1RuaicpRJYfcfMaTSVar/g
DZhpViLicWITw2vb/3XjSZIb1c5VG/mtQV2RLPK2GfTWsce8nnhMejuVdt3APVv/
EmsTn0aFs845Y3vpwgxWAlCgEZ050Cnmq6IctGPN6ofv1BTzjbp8TRm1RJUHSXAv
MyLBPfSSYSakPD3HndczZ3JOcGnSKZEqWAvbemkiNFkAFa5+opOsMvGHTinWs5g+
Gm2cHxJDA7FD1ySFyO7ZmK2+8cUcyP2pCas8KJyhrSkWPVOM37R8szIT9xdBH+/E
O90NdRwoyymTHwHIl9dwBQjTttQKoxBqpnedWoyuqUL46G8M4D2MImbr8TSa0y7s
NF0cNa43Pr4CI1Vl4gPQjAHU/IJ/BtdzgJaet5QJJojCM9QS7mzwHaTRttk48DUL
qCPCqWm96GIvB0NMabTSKAiLCBfZMdgM+6NliarkkVAjc6gt6HqyDlPciAnAZunE
haLjUIA+1SsTZQXWUltADQdAu7EOUZqXQ+vg7EpIk0tG9jriBHXxwLdyRzYnffR8
XaNE8izfHFt9lb0BiINSTBjKoc5yion+h7lgaX6J/jrcT6VnnpVcmDtHRxotkN2y
qUL/tI1TLTga0Kxi3ny0OqIG6eq/obBDV0BFoDrEAZWOHz0v1qDSlmUZB0dWKyF8
58CYM5VnhGEVk8YT71HtEgXQWIGriEcpjkXxBz3qrJv1zvMHYTHc0NzPtNkJIal+
h4JBTzYC1Z9jeoyzEYaqthJkCdXpAtSPD50qdpTagxt0fXSxwY3XLNVTZ7qJbtep
qfPIwOcuTpyGZUvb4b8RF/4gZtf6h4W4GAmf56tx6Ed4NWtAMzvtcOCoBW1TI2WL
cxxQ83DL6+lRXiYL/f7tKKgaef50cOYB+X+pg2j4IZIL/FYbNdBC65HUX5AXuG4F
lPfCJkQ0Pj4maiA2VUUy6qBNNIcBFYnovak4JrzJE62wIpdKp5D2FPUfdva7V0tR
9dKZ6FcburHq63Sh4vdx7bDHlBECdlyg2tYaRYUBbKhw+yw+hfuwjOELaX5VPxz0
VAdYtTRu3lETlaRJizuqJo6V4/GJ4gQ/epBvML6GDm0V5lS6kXrhW30tPVqOSXfw
NnXH7EgPL6TQ5/dTyJbd389CW39oH/wQZyZerp8E1lV/7WD1PYcgtGN43HTVIN1e
Nl9rE8OtU3VbES/qLOlcvz7zo2U3Ukes86tfSQWMzW1JbKnL4xXC4BKma7fgC1vI
A9GqDVPIjTcqEiA08O8BnfJuZosYiWBEYo55fqCVgopZCX/5cbjtWI+vvpuPWeOM
JB+aC87DcEjdJbF0qSoPNnZ49x+JX2QvCDRdb3i4EayOuI1g6z8bBiJPpxQjpl9j
Eax57sWfwcalrtEVScJZAfZrH58lNjuIb9F1hQP/mdCFpSmVrKy38NU80zSEDHKK
/xxRK2Z0e1W/mcFPacdoT/UadI3edtcsRgvBBP1DIEMnkTwIbgNSU65rRCSeKInz
1HCjAsed9RQyKEsVu9ZmXrpsICa8CLJKCGHv86RvOP+Wxqw0P/nAiBmcAfrWVi48
xCVppct6DOR1lDdCrsEJ7/lMKKt4SZem3R6rUp3dsHbBDSM2TG7dkbQ+HLyYe9TT
gGkrur4v7enfoFVvN1e1/5fdb1MI3F115Y7mQbjnsA8Qp2sJ4s/jAZDR+Rcuddqk
HHsjUhHStOcpNizE4kDvGd+136yIDzQlpWwB71B4h/BiEGNf5aGnECkITAF3lr/E
JtE5zUhgoB+SNhFzWAgcslc8V3JL46TrZTkgcECtTcz8cIAh8dHEfAmP51s0nxKb
mFsIaPd8pjrOaZvNvbQjtDivjAJw5j/lLwDL95V2HAgeBeKXxe51svculy4FuR82
wCdmfTTcg+q1avshSzbnAyrXIDCIzofL/1N5CPTUGqYw//r8fx+kpDqxy9PHfp4D
BS6f1bn0PyqK/0z7YUWZQd4f/V8toSLgpzFYRs9SzW0eDRp52lc1s1Ziu8QjWXnb
wLiTj34f1HpLTvooRwQRbUoOg/+lCSUVmm5jwRnLLPYgvlG3Hx0hUxs/gtxvC3qb
e8JmReXqkYphO7i0pi1hU636SexRNIiGF/gpsUozVpgBkR95kf/4CUSX0mVoT+iN
PUihx6zpc3/ZuphVCgYBQAxTs/r9HzQqiPKIpwc2Aq+iU00hG9AyV44OMdniY9Cb
FIKalaQxweFpaUn8Q0dl3ewtg3Od7SdEDW9JAY9EkLlArAiU+keq+MLxzdU9zBkP
1xkfkbB3RXMJqCSw5tLn1bBaLwGM97RAXjq5zWvnpHs3GNPCrCLXGfpB6kbKB/mc
4XEuvdt8bNYevEh7ps1fx8B8aXxOsFLh9StJs/e8RxVXN3XNq8VVyF5N3fdiEnjD
M/8YvtyHj82/e9gjX/zdZ2zU4bRU8x1TjXURjgG0mc9d6DXXvkvjk2jQVxGavBov
NYeEyYzyH2llqurREH7Msvc6545UwQWXeJ6d2q9ZPmnpr4T/wVFQC0bY1/QQQddb
U5erTOpjK3NJNZJ53x+RxWISH2bJjjL6Ikl34PD1j9PVFz65uBX1Qa+1wsfOh0C3
BQYp4+SHI4FN0K1DuNDhd8RsJVj75/y7c9MHffxQXyuTLP3o0j7Svx+kYq4wqd6F
dHd7bWJZe8tWw7ZHPDnrS6ZD2iSWcEU8v9zXf151x/7CntepVrqWU9d1lOvsAg0r
7DcP5GiB+llpg5djXS72wlphKV8/PSP+7SEHw781ByJfr6flQM8dJXAyA8Dw0FNE
lyQhbEmX5IUBs0nrVuNRjtAihGXDu2qa/2VrF3QqCvVEI5/oeIyhVWSGspMEoclD
Cn2nLEdDkiJQj9BYq5Sea/cwA2PswViEbRxt+LQefBL4DKNeWHgoDnCMv6V4JBwT
qGr0zY7/gxnMgemeuFSsStT6nRlW5z9DmLj/c1hYfIUvPQiIMFBRFUAdbIakhrTC
dpoRI1d99zeZcafHuxphk4gJZPtWAkqyDtNHQfjIzXvgBUV73omsAquFLQV8xFF8
XS3Ea4f4KDD9OWyMpGUg235lHyI+zq3tNb4bgU2gt+g0m+ep4LfU+CMDP08vC2eA
PJrlTJpf6LM4NzNGywiaeIuk65l8VXYl+OGyw84hy9QZkDdli/C4ZO4fl8Rt6SC/
3DQvGZ1l9wUecXOM56glB2tM3ONAHoyzwzRjWSOU5ycfqkn/1HMs/Quy8WOzKnVe
e9AsE8U0mmjGGkYGn2Hqm5JMtptU4Fjy/16i9ufOq0dLm1baZvkXkik4Z1SqNyfe
yUl9QccmU//pia6vl3I0fjsAeUEsEmv3oPD4DpR6qGzKxpAIEDl419ZDXrA0isSs
sb6nqn861VjHstJaM4D6F8Pz8LN3wTErSON5um1eO1AFcl2cLMgyBBAtQzwq+4SQ
k2lJ4cLCdpXja2hkzyknvWHCAfUZK8/Gch0OWmg4uY+s0PyrU0H7eYNXK+3SOSnM
0AsHs7NUIlAa6nWIjhigohylD0qbjBhP3Eera4ku2n2nhIUdT8tN/8x4Z8T3o4aO
PIV5Cs/c5ytmD9M9QGmhPk09Pcye7VYjl/XrrcsEXPSd2fBxhtOLLcMuIGBGLTeE
BSRPMBvar/R5TqF1OPYjXgGUkV3GcuKO2VyoVpEJfL/dsixaklnYtwqQDwCU4rGs
KmSXa+nj4ylgpnlH3Q/HPY9ZZPYeraxkXrgOj6OM544xhaLKBgOepf0OnhtdcGPi
RzATiIhGoVsES4HUmnH4Ew/g49SdYQOf8tzPtzaLlkxup2b57lktvTJP5hgbjCUe
h1R2dsVFT9FwBZjd4bnfmtMMYoxUG7lAZ664OPZUohRgVjh+0v7eP5OCf6lgNydh
KoG6u7hck8pNMDhn6wMO4zEKSw4+wgIBTI1vsjB17kY+maKGIDun3YVv5kX2/6RZ
btkS9Rj3qVvg5fE9aCZ3qT6H6ITJlShBMDz8bAA1mLxfyUkzem9Fd22B6zVqFsoi
bccohiDSOli3rzmowJQQoEd1d6d7qo/vwQ6nnZBtIhH6menGYv87lgo9T7WKswAF
lERQuCGszASZAk8gNjiJUAT/bMyS6Zfy2uFmYz8XYhSgVvVDx1YMej7/rJ23Ue1o
mKkqP+y3HG8nL382Mh13nteaPuiCT5SqwS8WZVKZSas0PPMa2M+EW800j6qEDRd3
WTxCN2Ghq+0XGQ0do6vkpAOa+9Ctx+Jt0lynyoHOfuvrJVq/grtleAO9M3nsLr4n
5DysSFKKuffTp21YxT0JvC59xZrokFwemP4mCDN/uUOLwidccG2RvVOxBkkFFmgf
J4GXYsxltbZ/U0dAAl7aF4neHuBxY9yty79mtr28oYiTjUi8qKwY43qoZz0zljp+
DaLrHB48FO0QLzE3lb787WW/PvO9XNMA/ZoR7QnSePnmcb6Eg/SoWwWyS5QH5gIf
Lufk0NTK/rWShJrO8LHiNEVmAkXhNZV8//36on9PDcev/UTitNMRBLu8VTW0vqn9
kSJR+2k6SjQ5vGkjeqUT/xbtOeg7MhgQjxMi+J2bEkwJY4zdIPCLr+FGpeIyOQVR
txu7r+/MhhMB6xoKaVYZcWt6abykgoCt+8q3UtL/R0nLonY2SQGuTG99pNVbMkgV
kd1bGSCtGYhnM6Y+OBzjqihDSWSIeW4lPHqthZT22a1OBY83rkCvA2k1pe6dJL3A
be0pVKonPz4d0BbZQC+Sh4cmDXPb6oVQaz8NqCnqJkFTSHhePOpB2TRcuO+I97hY
rovuzU4BXtMDHtP7z8LvYEQhrzlfTW9ghy03oi6qLerh9Nk8i3EG3QWYAp0EEIM5
t6LiwWaTDp1sPlliQGurklZ55gCuMWK3eYfC57sQ3z/9wkJYVg8yj1do2ebJg/v8
Uwd/AbYygzp/ZzcgWZexdk3UxCAfz2uoy2MemSiVFOpXfPvYLO6IyXidHcwMYPrs
q+MfpAEAQNcWPIi5X0xI4Mj5fnAz6V8aVxXfP+Gsd8Jlg5Z1LuKX328/VoawkTyl
0Md8IVFpANs/z48xXLDrbdD5rGAI6BCziwKarUQcidg3bjcbE+1RBtT260yadbcD
Uw1vxl/W6DQ3ynS99k/ZRYYTb15uL3AWSebkFYQ4/KrKl6d2RslfMM1XWMXFFetA
V8UBBaNAI86WJ5S9jk6T1vxpIpVCj1YdhCVQgSBAl612ueQIJ/pELFAuLBtgxWBK
msuY74e+Oq/Ab94HMnHkL1M3HGK5a54cfnOr0Wmpu3vONtyM8I3nRM3zrgmvCztj
ph0/emMnopcmp22BRzSlVt/qcK17GuGZScHVoiF2cCk/1YL3JOB0GxfXblG3RH6A
YCyn2qUFWqam8Rm+3fdIF7moeKxLj4Oe3TnoYr2Kzf26aDpbiRuR2Zdk2KT0TOxl
/34vOkPgJWmg/h2b078jhun21Uy0AE8LYCe3SeLxfO4muwxMIkUzn3ONg0Sy6rMg
CUhenJjUPJaZuwENYxUAi/rE/n0RADmOCU657v/AQE0+FyORGlJb+jReNi/7Mqfv
ETlLrhkh71mvdJoaMalvepI0+jQS4x8/hOWyWbckqcg8M6yNIih/iVjG9iZQL97T
7SRsy1s3DD57um/QD/rZCGsxfbVT6Or9Q87hUt81N9JlTjqMYl7689mIwjh7wPi8
PYjmUld41z2EnVNsC9Xs/mN6GKS1CpmeOY4Kxs9/gZSmGQCI1ZATHRT2Cu48tVqR
oq2iIAf0sJNLsb8rLK+hgN76goQ2h0F0Sa4S2VsQadEarCLmn/2FuUiB3fJLP49h
T5l070g58lEFPiWXccm2bXBKp0tnQLqb/AFZ/Lbr2YTI0mTGW6ZAoXGXjLe6fK4C
W04hcB7grPm6m45h+yQDsHnuwgtlGtvmqLZmYuCbUgmUpNTjhFEI/ROJLZyyH/WG
34ohb/kDKFvB6oBj8AWCclRNqPqctpkNPGsST+xl674wyCkuuD+Dj2eSbH9BLiuQ
p0zpF15V5LWwkFfy3pquIdBRWH+wF9qojuV/MWo1OQyfvUyXpXAWjnmMSBFySx+2
uSzx7v4rpnas9uiv035VRCeJbxzcfPazSSIWQTfeqSzmVSn5FJkYRIPCAIybCnp2
zylcNrjp+yfiud94ESbRruKTLzgZKH+Uk4Vbd+bzuzrjSeFfBFfzZaTuPWMcPtix
rKysnpbCcIl6bxGD+fahvcmyB7/0xS8gK6BXtq2JI0WrD8UjIgGCCbusmsbqIoG8
/g2nke20N+fysS4LtDYfOwvErN44gRY5nwDTzSxKG0rAkmUyx3zPKzQwRZ0TYUa0
5la7UUMKzwZBtc/tFSRsrNSzs9Lq2BnhbS9HMx8fWiK8a6j3smvONiD0UToRkFHS
Sj9pJZRT49TS6gaBbCHdz9hwcU/L68+aDlSMQGopxqwFjhOEdnA1Hh02g4ta2IRE
Mjj3e55E+Rs7VdraeeIkdyCGjUkyOAek1P0hNbJXsdlv72930qkAhktQeEPrWWVN
pNfgUdKobFeQdiromED9j+n5krSKMq0BleMrET1+4tkgPLQY0J+rkm62zmjzJxn3
c5nuOHK6CZOkckDM8Nrojl3YLRKEwR7Z/tN6W4nqidSGh9pc9P7nMr0gpcnL8fkQ
cFzI4on9Ca4uyVrN71kYi2CBJb0Lgk66VXZfCXk9+PPTj6pXSHk9cyDwDawKc4IE
kQCVRyMg1bQDfDDr0uui2C4g4Q+mV1GoaVL9s26YtGIk4O1WRvsfAsy/0+v+cNYH
f4Jrhj5pRqNu8LBVLlCHfuLBk7eQkL2bX4VLN0ksD19kN8yfIQCr5xdWl+/7QDh+
ScU5rMzHJ0+T/33U/3gxuTka25f7k+2LZK5o2XVqjfhFB3KVsaKiX4RXMGFyd6vE
frBMX1ROItNdWwq4xNkw8mld6soGFeWydQPMLwf6rdMwkGQ8wPoCsJ0Rq6gx9cJ9
H8O+8mwqKeW3ftV4nDtS7XuoUMt2aoUQ6J9UHe3xgxZiI8kT4iM8NbBM5jV8gtOQ
UUpctEi2wRZw3KwJWIFj/P7eyk2x+2EGfrm10pHrypsKJ9yBHs1AO6uqlwU4wlPp
XnYUZ1iSMabwRq8qBpoKi+5avxnbZt8ciVQ42X9BX3B8LuI/WRfnTWhUwxuhl2Nz
PHij9ibGnKPdLfUngiKS0eaaiVY6EUU0W0GHGrsV5auZt2R/jnWuIJMfR+6Si8J6
20X0qrqaIhgUS4l23e7LlFfwPmnXXYhDJocJXVM1OPj0ZeMJtjJRMjuxxTVln0kH
rcavOH73f+u7FyQn/+VZpKviUZp4dqQ/8QB7X7PzyVq1q1+IvjM3TjADPdGOZfyh
Xc18p0LbHZJBPCpY4Hhk2M/RSEOsMmP4McYhDyYnE4JOpMI3w6a7lyMVf2wROACd
p9jqzSpZ3eZLZGaufwJ9tqhf6qh7xUKudAGyjGPlU3GZfNKATSgUY2gG/6chtI6h
b0ZwMPDUuSrGEsOU8RYbHn981UmXqiZpmApEj78K1bGouV2nPjRV36vNs4MCPTG6
ie4BeE94/m/2c8a+B7zDxRLDSyWkATrJxcaGegx46Q783TMP0OO/Whc0xtbaEFaQ
CKIy9Wqb571I4K+gsU3uyShAvJ39LNMBU0Y1y93nqBMJWxjRO6/2D/zKK5Bgp5dY
t1qHdcKQWi2yJjNsabxzrR2Mot4/VK9haFnHkpXE7+9BWoJjoSaECU973fwPdtBN
s1E/whsIXnRJxG89GdyNGelZGhBs/v88Ktn2z3nNt3rN5LKrlxUNznM5tbOkbO8F
iTgAm8oUFx+KvprnPBBaqGN5oOGZSxQIKZbnPP1E6TL7cHQV6S+D+pz251ia2E7h
FXgGeHkDjkJax2+6jImB7fERmMK2PWE+kE6NiOjZLIDYb33fo3ld2cVnGYcR2NS+
fvUiwDPSurxcb5dHUWi48JBBpxjrHLZVHPrB5KmKror/S6Qcgqke3GRhwoROzPjx
JBGtZgrCFaYRONXs8LAe24MRtJruXbsy4QB2TJJ5jbWvwKK0p65JsfjbFtjTz8zE
bBYScd7Wy28NazZJSSUG9xrbdY+vm7UyjEAXTnVlkVs5o6WUBEKTwlCS2TtcKovw
qFAzoe64CbuA9GWSSlQK5wWLnn4lpFOrRuDJItN/+W8mr1Q1WUADyNmqT8SX2qE7
7FBzs6p9Y2YYLOvhhnVhf2wHNwhBkAJMAwO1ehHuO94kz7Z1pKlWJ8Jtje4yP1mR
3BT7BGv/kFYHqkvfAGnvS2O5hTdAEtTTTvB/GryvY9NKPGRGozCXcSXCmL8PZt1f
0suZ0jq/JGO1raw3Ji9ryoApQvqqjHYEF4U5hsRBW9ucIWbvP4AGZxUI8P0Pc/Bv
VsTGjvZg0mViWKer7GSCCwk9dW0i4p1HDte3EFoVWOegU2CpVyWb3vbE3CUbchYa
0f02WyGl6kosbz6CQSL4bDi7OqQXktxupM9HWn9Kn8T8ER/SrCMjBTrdc9y3Wvbp
C0nHI5TaeG/D6dOq72mD+xYj9S0NTo/FpMbHwAZP+350ptSyNfUjtLBnSpMtEW/w
hSBbH0f+dn1hZ4A9iCqbjrmeebAsh09/a95Bt7/ajQeKAu8uinKzcKLQCki9PAAp
bkNvANVjsralcpqkIPFZoVuDWHp07cZThfkZS1X9KVkth0MDlpwNiN8ZD1kfnRaQ
o+Eyr0E6WR9mSmzeFyauyzKxoVEcuTef9lQz7WOrW6Z+RFgWibsUksX6vG8TLk6C
z3YcedxkaTeR/znBQ8ocyziS6HkSFtYj8kZeAY1pndrU2DSNiVZuECSPQ+NWYrqu
GoppH0QH9PoslMKNqVp5WHh/Mpg40/Zs9vh29Rmy1qsdgNA9Vzob3fTDcI7djTWI
44xYGjeqT5QoHnVnvwkm0GO5qQHu+LjY2zaCayeVyr7wNwg4GVtZGAYCsLcAgE/2
1rLIvomERvh9EnwrmvEcP8FCGh+ckLt1n0xApC1aY64BgEWcdaZU9cFmI/Kb5pZW
OYrFXWN37wmXfk8fiFHvranDv7pU9XzhYeRDqYsEkmWU8Jl2YY2eyglAK6IpqgHN
VzAGTuXTo3rHKtVowrSy1PfbCmKyVBNgG/aTEbGtof8PzUaMxpFQ5qTPVL9sd8ZJ
ULpwmnKPl0Jz0dF/+06Vt58b9uB7OraRSUZ7EpJwh+BvYAPH/2i9oTlBsIIkNR1r
atKBp+/dDuKczu0EfY4na265vjFAJebOZZMnCoqsY22kKL0Bs6h23ouEi0XfYumL
sDGrdn9/DmoM5iJiJ+UVVDfQKW/MEMyYEWgifV8uSNaZsLpuOHfhWoi+P+cPksqR
CEIVIkHw/sh9+PkRg0tI4ZOE4ffeoS4HUlBiiPwm6jtlNU0S+SgkRBRZCeGZf3DC
OFhDVOh+qhZbiKKgdSClHh51zK8EhDP1sDpg+LMyTtvYowYvpFYjvzppgU2lmfTc
ikfT2oJFETMFunFb6N79J6yHlcRp8TMA9epZu+PZPJz41mxeb7yooj16S3lz/Tr1
II7ny56Pxnp/l5X95UMNUTUFAlbgyDtX+2dr7GwNG5iK5TZQsHpXi8XKHI2IgrMV
BaR6t7kdOthIW1rnse703msxjYuXZc/wX3qwfVaS+J5qEOuJtwwVoyxmQE3syc+1
Z9ycRc0otqeY65syC67+3mLzhqYrBJoKQavJZEop2OIniu9CtnPIJerLdRafNS3A
3URHzlpMhzsT2cd5vIol1mY5Uk2lfmiQWzFojAD71wsfXkrmsNCY/FaiupCpLVcV
8zeAi3Rt6BDgKD3JWZHFDaeNBS4QHOeV1KmrJBNb/qq/XK0CG+1aHvkzFc3rtUF9
iOdLlEnU7kO4hHJ+7uYI9AQINj5AFNBvSVXzhfkaOrlguFJEst/qLNjytYwvf0wm
f2h63aWcWE48oEsSAwDzE7TbhdiimYo+z6OKyujul8UBW02CnsVHLmf0FibXZwXa
sTYSA050nZwMTr0f2ukgIErZIOK298ptBfVp35rNBeS1l+v6XETS4/lYymdZ6oz2
OBwCGRByaOgxTC3YYErE6bPU7FJD+/cvDs4kDlINEj1UU8z/OOHDdJ9cvx5iXdv+
ZEL5ooxF5Lp4wGlkjAAf1bc8oDqZYpnmUcJDBUpWqq/UxzfySgwRRBAsewr7T/fD
FnPnu1C/v3pctu8RVdkcEK1bN0bhndgRBPl2UbEiRdkUpmwt+P4EFqY2BsyNqwf1
hy1wcZohfLdZts4kuypQUIuRttsisEviY544lA5gHpQpQRllzEocBS52C4Uvfh7B
aTxcoHDQIJJf9EzRggUD0tHvbY36ZxVofk/dD2jzJRrkUC9dDoPQPR5V0BcOV/5x
/VopVZ73UBQ2WH8lTXjqqt09TyC1T6vj6eEAjVx2CzugxSVMyLUrS6wAA8K2+2Hi
ORUYYWyoZjdcrWlykoEjF/v6zXFhVAqOMNaDNJ/P3Afb9G0vlmltHRTlBDtIkGU3
ZRM4C4020p0rRmu4751GYKYFl7dEezTwP8zJhkPFxLBbH88kIfClzdvIpLuYHfeA
/ub1N7+krixRc2Y8eoQxeXkWfICra6cvY4s2EtPVE3BX/mCyPeEJjf/qlU1uG6eb
Y4spMBZqDzOqyuReRiAoArCevMtYjbilcNgof1g8HJzba3TdJNiJ9QsjeF2SzWH0
1I1HSzrfTCBfSCTvnupXysPyEZNMsGI76jh3HjuXx0FqOcVsa4gp4yid9AJ0GjSZ
s7OEoNaXPum7LxKF2CfFYb7zeBvAPhg3i0obaz6xa+sAVdyNiZ2eW6wMHI5+Io7S
K/ClVb01hKA3aJWRsxscDbmnWNfA/6vCLTh5FHuJH6WiAOdfdcBWt+lREOBuOPei
EDXHeq7OgAhm2I5/7ng9aphhme39p/6AzXuzJLbmi3WbYbZ2a/MaOdGGveGCiSrl
tnbhqkLqrdrJvn9R7wR8CnoORxxQZ16PPzwzDvAfU7lYFxRmhNNIX78VA9ODLqMV
1uCPiUSCR8f+z/TVXVskMjICqUf13FKdFFdj/fcRICT2zZ5ciEjOtThsnBagUlnd
Infeh7O5w9MwANlmcuxA+7a4Vvx9QObE1YHLviD0WWco2Qr9/Sdf2ZYkVt5sjni1
VkrcsOS9EzEIrBEdnCZM+5ZzxETHNq4HUGjkq//+zyoenV7DjMPaioCDnfyHKBeD
HI9b7CAKGdX0lYPWNXd1oHzuyj6kYhPsdhoKEfm4pwSeLuXInnmHRtShQxbFuZnE
9EX7ESAMDfTlQ3CRvKWPH5iZ2pJIhbjhOxRIgCIqu3W3j6M9+8lAU7YxUTNBGtZp
M0fG6a7V7XXrFAHTWrlulyYaOMQZdOF9Wu/y13UlxwZ9IPozClUKZiYenl12q3sy
+VhxlvZGeQnobqaBn5Wd5lsTqGw/wGkxPqOhDpO/4yWbivhWlyruVeIlrG4fDU/F
4s7l8dtHKlYU7wbpoPGav8F5Qju/I/sJSxjOCHzx/hIarLlCM93kxwk+NUwSOyYc
XhygVFaz6mU2fRG4+rr0fwag7+ReuC+BJLNzVADiIoX+hPhecoFy0RODoXOp+0fX
MGSpkkFUbvdoiROTG7iN7XhH6MAxOF8+EgtW2kKFzxQZODq1vTzNAk2fAfKGmj8w
4jybvM4BPTE0SPKDZ1BjtIo/d+1iMbxJ0F46OHI0YV/INfDLyR57FuP2HCdW748d
ghp3wWneVrhwClgxleYAG+qC0EBaitdkktf2Tqxta1r3s5PiTqSZdtAm70p2mQAe
gJY2QbGeOPSmF9uRpZbloxAvF2a7ph+pcJZT8YwDW6UeGHP/5Jvo0TP69hprTaNV
Jpq/aXoCLSS0V/G7ycrt7zbg1Or54bc+YGbdFhP72pnBziq3491Y3QM5C8bJJReH
BRNwIJgJuvs9xmbHpjvMW8SKccltWVnd2CCYFJfs8jkHwCEevjYFez5ewZ5pRoaU
9BQPcQjnv5HjMbllvqxVrbJHajrh1I4mq1dYxnDnDbzcITFBD9PVUTFDy2JBaoEN
2+UMNjWqz/CZat+TNVGQHA9Z6pp5BLVtAyBl1DeaLNWdHGcpHftMto6vsc3y6Ppt
YniQvSntt5zBKr8WNWYH9OjNgRXwalDhHTkAyGfbZL9Cb7t9fXJ7Q9bhlHx3YCit
h6MP1+KUAlPBcxw/xRhGVBzTlSZyNgLy6bnKFHo/2DCAsQvyI21JlT+y3dGPualG
ASHzqerm+S1/3EFPe+Xsh2qoM/b2yCP9rPNAlYmb+Ia9MmvubtZvuRwRViI9usuK
95xCDeTerPHsTQkilJBiMtzQuLUj6g/PUlnKIpQmt+K1/QO1PzGzCzKVu1K15RGm
+u9V6uNMT7jhptoCYCbYp56JJ8YNsQNK81vsZ7SRKjV6xqY8MjzS6yDkeZgX4lUb
Blm8igZ7/4eRSGzMKNRe4ED0usq7Myh722xllAYTuEm7wgQ9b7W79aebeP5tHshU
l69XVmHd/dgafYnMzX0Q8YkL8lYDRLDr/sSussc4H3U5jgH2mtevKMurbezKNfXJ
sMGYcaOE7lb0eUM+T7WfpzjRCWvVJDrNyrkUSpYnJfu/gu0GHNnT95FZnSD854G1
Or+0YkLljTbKzYb6tB80xKKtvgc7szc5/1hiPD+901HvWopd45AM9+/5kNR1uQRV
ahVTAYIhNVw8RnP0/W4T6NzRjvBqmmlsgPBqvYQGo43tCczpOl74IfdVoJpjU9gT
hdE3kBU8I3SXF/weJ0/JBvcue9muZBVqs968TZ5Dr6fh6Ho7RNgGo19Gc4YHnRTF
+WK9fTJcTUTCJPC2tdZ9P2R0cDooDrhZV3hhh1BKD8PBFzrudSZeURt599qlmLns
J9JKSN55UOIm8nYiEPkBnL13iW2QSr02D/Zv1EzEpJCHoz1wVpVZimavO9erLNjm
lvEBxPMsMTW9IiQWS0XWWkcGbOA+2v+v7NxvylRTnS1blR2bkSLPHSkEDb/deueg
ekELH0LF9Lgk/EdQOoc0dqfUJiGnamrPghIUHGXJmVHB9yAJ6jYE62lZYPV57bdi
O5PEYERwXOEzrBwTpKLpk64xaQKLGRDZeev5h5jY3T0BX6c4O7+FF4f4n8ydRkq5
EsWXODMYucbYqdpPn6rxv5IhqNasHZb/3z+fOJOLhTM4A/nuRZ+YhUV6VamsEawl
lU9lYJK4pZlPw6jQ+D0bzYzGKc/CcKSlCFBnmTHJ4SRAoejHoSz86wwMMvO7aUxL
1tEP8Vnc1l6DHLahFkiAqwgzapa9TiKNDCN152D6MTUykC66rdRRQ2ZCDn0xKwjc
kULBKlVZDnF0oGsm13jH+rlHTNF0kxw1gkkgyH3MyZO0wLITtWymGIU5mXhDnqiD
315EoTFwwPIH0JgZDqTnG2BdYgmYn9gf3t0MNjEr161EMesbdAGzC4rHAVUi4rmL
rUlacx5mm4zRoD4O9ueiZGDtGdgLqIKBEWHb9fYYhNQ3qlyCg80E7TAKjIZa4mK0
6kYUJGe2e9OMpDf+PG4LsFDuhT6cShWa+Jj6CLRn6lZREnMpSH4v7ag/a7lUd91/
rCVWU9jC0nRpVzF4Jyfdv/NE6BuE5v625KoxRpXq83m24le1BtwK6kDytI8BIjDX
xmQevNhHXz61JOinxO2NYztOs0dH9iKpx1u2POQyHYKfgg5b8lSCK+v/XoYOZpOb
MBc2GErwg+adCRorvm3whJr0lhJuq/c1rqeX6HYYSlbHQVn4Y/eEg4lCSF7TkXJ6
NWhGFCePK7gGx2Uvj/uupPdIJqmwjmzhcSO6bfneHEXLt8pHHplKkfdA2c+eoTH6
8EOD1nASXi4dPyqmKp7wRgEaDvEiCfEmOXxqPzohoC0tw/Yfme6wjnp8bBpwnu0J
1UPyvx7uf3uT64vmgjbN8QKNNx28vJR40cVDlHBChvOEzdUF3zYXiCWNY/d3AtVG
hssVOi8WJ1mHUDaNlgKpViWlxYNEPko+HOBUwbke2eKRh2ByaHob6xWEXW0esyr3
lZ3HRp9qOKblW/InEtUVG/tpGaAJe6+hibqmTcfxupOpI/lYJH0QzT98nRGan0eN
ckCEOJ4WB9kgOaj5Z9kkzlFhY5wvKMG/hJ+Sl+W84zXHPvVjO/BhJ4PnJih3j0DT
AIw7AU5fiXXeWQg89bFke/HeFnuCboPsLZ4J7w2Oox8jQHgsDhww/gUrG/Y0qTa4
d55PDKybgPEdeUSXzgh12pyM5Yw3YP/BRfDDWAVHCzMn1w2VTBjLdQVrgb/ceHpU
p4Z3Vq6oJhzvQ5N+fpePzCNf5iCOgDVdVJTqAKEf4nDWj+4IdM5m/safhhO1gi5q
Z7Jd7MYVcbW4tEzQiQHCJvVT4+AitTvLUUoHINOoQPwdb085WWKTFwdULGrsX8zB
zrjSe8+RQsG5Q/ACHJEy5ZpyRsLqi/M69Fe2bRy/ni1+F4ZSgm9801OVc3G6znCR
ycZ11WDV7Jo5TYvTBQtn9Dr4EBTCuANc9iiSulySuHJqwRKXUvvuW/wyoArhJJT/
Bk+jvZ3j0DCQ3pNFCbMluLp3vVgoCCZc/8lYGeMwU9bVLxdt/fTSixMlgESwnwYp
XUW/yRO33bMqo3Cfse4LfCnXBr3JX1avR31fN5ZnRAZ/qrAkjWKu56W/V+emTZnA
KV3VZifWo7qbAAi0OYAF81W1v/6CYo7J2O4S+y4lGxmUVv66zbo+CORpnK2m4w3o
MzxzPHyCsXV3VatsQAorGqEeiy+Xv50scFxO2GEA07fC4ccagXDuE9bkHflZLuJT
uqPlRs/WlCbvV61de00P4oGORBRjs1hihK0glviIyBbBQqjbL7IeRcHRGQ73wobU
lUlksupfks7c4m8x4sYmW0GVuRqFwvxaulwPu2uRVrAjBg0ZL3oAkIIZZJQUUpfB
2mOBtSajOw4XKBMyIOpcVMM2CsynQ9gZKzHE3YZm3vODoWIygw15EcYOg+86G5uY
TojwhtSC3bOfIN4dYkg6TLVA3rrm1roE9OpeidzVpBpuYm2+SEXgaGFYj4pQ8mFB
JJSVdZFtBE16pgnOqVrcOXHm7DFlhNrQDSV59GqDXp/F28fpK37257ak0uWfFkvO
x4ol2UvSUkjtRFwNrPWilR7/I+OZhbKDlbzmjtEcgqvOh7YVZYjbz+4a6TUFrq3I
UqnxpO9mMqf8XDZVgk1Ahj7lrIsiXDrZfrdkDH0JvhU4zgq5gfzNOB2QKcqwVEVN
/Cl0TESiVmn4RKN4yxd/xwxArRxyOeAolW9FIC58X44gNq8zOJAgN6f5UiXRw/FV
yZpdC2rV50VGncGVoyFTijZlMSFnoUxw6/xssRVpYcSyQloNcDw97JQhQp0GH2lC
3L77RK2o8E+WjqaYmc1cV5CPBmI0vdmzuW+MZrfUX98vILQVB6870gPctl/YIZPo
AZ1ARuhZ3fqlVKs50rqJmppBn1yWgj4ElnoFZaiytYIP4VI7JMO3bti7dE6UAfYv
+PLljMzeHk/PPVBejy4/8X/5AsqfFMun6DPZHL0fR87LMBO1UIzGeS8cLljVQF4P
845XQRVtf4ApJIbj9949eIvRz903zoIbDdSAyQz7HZbG8KkNL139E6WMD+/N2GLr
DQ8bruFVTe4wl96UdR6O79hqzxJImZMRnuo80zDGy7XP/AFqn5fENpyAf8cO0PJi
EqBqTMEQ0glBhkLCqzoKQZmSqssh4zQ5qfxMktHUF/4s6znKWjFlrpZ08Mst7mD2
rVD6SS2BYfacfmqUxIGG+pl0sbMHzV581177CXClZnNSpCMgvLnCXYgmaBKx2aez
nx2WaAkUQAIeVUft+FRVP36WO2H+PPbi4fCtPnvjLG2+0z1AAfBEUMWZlJLmndr9
il39Db4mTwawbY5pW6UAzB1yTR3tAwYGmdanUM0L7HvO3CsEcArrsp7H48A+FpE9
5NhOzyMUmTNDYktfkIl93R1SnkHIu8F8I8kKaEavRsr5mNRjHNBaTzJgp4OcNpjt
8fjj6eHFZQubo1vYBd/LYbaANg5a9iZlGRkZ5EVKCKvSidAfj+KhK7C6GgNwy/O9
0qpC2WftuJcwJX6egcQTy92e2TQQuEdBPox0xWowOo5gLRbf/4JLll5N7vW5D/VS
q0Xo+oNSgaYXTzmuH4Gw5HYErt6si8u93iowC9YU0UQXGy1ZG/aVM/EUvo0rzpDR
iOO9AKKdUB+oYXrEUw0hoE+EuohEQZqW41wA22TiM2kT7WJJXxZOoK3ALAA+FHMW
Kk1ay6ih3+H7xYJJPkrMGd6R5c24S66niGRk69454SIjkfVo7MVBdbu7DXLGBQhq
Zmx8Jrfrx2O0sM885mwEJ2fQ4yFGuPeTQDPTfEOBOmOnYaCjRJ1NeUiJJ9j48MmD
EBTAWhABo8/pCW8iPA65kjh9b+jA3v4k5BsOieYWTGMAyrdqPCTBqBjpBa0ehVKl
4zu+XJkBVu9mFeB8UQRxPy9PWnwjZISfhd5olT/YuXczhhR71E9VCsHvMaF6E2oQ
Q4z8jTcgLA20xJCmz0DYEOXiOv36ta2UHkWAZflq5Qzg24j/G+6iDX8qShSNUbjC
+M1/DdmLmd4PK+QJE+XYUcvxGFJtnpP9OsTbCxuYtA4ZyBu9604ZLQtPWe/jgGia
z5kxNJhiW4nJVLzE1M3JsPd0m9ndn90a0Cb52z9+gSMFzqztv+kTfJQq6188SgfO
ebUgq9UCkR3T3tzD7aKQdZff3G1WW8hsu31ukN0H9MIzKHd9YGENegQ8ZBSWJcop
Ee0JxyeFz9+eYLlyTRIpuGAKu/2fSdVjAehloIWWUPcFGcvdg70lSzX07hasUk9F
LxQ2w9QWkfZ/TA+kEpApj3pRnwrPYkgojcwYaFlbCaXtlqNj75Fl7AdtHb2wnhXi
4kssbX+ys96Tlurm2LZBZx0mhn6ay6luwS0Bf2pB0MWXRXNVmT85/+IQeKOG6DsM
uNERgnO3DNxfXrEnP8MM4ziJbiOaP4+8vgrNCFKSDEN9V2Jzp0nJT7/+OoSsfP6a
JHQXz6C1iZrD0jxfr1WMAtUxzL8l9CDKlrjOLQmxTJV6fWc7KR4DfVT2DgmOx2kJ
iaAK9UZ+x0yGLZS4DyBVoVzuSu6IuzchGh/lEtR1gwgzIFPipUs2Y+G7Fn7zMFUM
7IMAg9rZSWmlyAkOmbcBByUQVeMUWhaR9QRl4dWu3A3wuzytrZDwhgrb0OAYNb5M
yYvj4ffiIxcU8uGETxbKh2jqKsxjuFH5FlGrhpXK9BtK91g5nsETCBJwPXfgmC7P
1Pw1NTkE7JaMwJwrDN7CO+ZvDbNZzqyNmpaX6qB2K+ObTf4oBBBBtk46wM4X63ZP
VWxB83zcHA8g35wtHYOky7uk+eogY/wTllSKyP7n+nOzIXrwWqCioFy9GgKxQ5Iu
8WsgQT1WbOkX1MHpO7yzbwdQ4su1ZpNIndeknNRUl4Gz+Ye6PmTjL6xj8pBg3Nc1
5AsDuQi8VeHyhuUzttcKn+9IVohxs6wKfDqc/HCB7s4GJppGG2AYmvtzSYIro2GU
5npFvbOpN7aZAa7zrQ+QnLJ1nV3l28dGunyqEBZBWnRya/cN4V2HHbfTWKpqyPAr
Zdrzu5kIEe7fAy6fHK9CUCM3A++jfT9nKGoeycn/ReEjqx9QYNhflR+IAa7LPeiD
YGw3pgIjpFAEr8wgq6edLGIFij7jpeKXVCjwoqb7gyZqHYUBjI9jKU+VXsE07sse
f40sZzETrCMuok6MiAjjcpioCoWq/G0Sr5xMlYRhkuFgwhpRnRguJWfrWW2AJA4p
QgXjCAnY9V81654CGCqHf1wkBzmV8kRrkhkvHgwNQP0njF2XOp45Z7IuGNZjJGe3
yehc8fgHXj1OKoCU4pW/LNB2HJHaLrtvFtZmwTcb8c2ctD8MbLLB/3BfU4olCaxH
SXWtyOPSL9rUlC6z6Htye0HNGQw3ZLd652UArHWNuiS+m/Yc0jVcsiyOaO6EvPL+
T/zNS2zM8bbAq95K3VoNWM2fElJdDWheotP1kUyJ4RtTJxfVSBi9qXuDJsKegnQW
Tt2M61MVjhU+n8LsBAe0bm1MTwP7KpFB0exoyY6xXhNPN0byEK9TRK5cZ1oeUvUe
s1PaEU+uqJDzj9J1fwQ77sPIDZ8H3ciAE9/ruTiDvKt6xVqJIwsgSD7nOMJb64xz
ue9J8USxyGiuiN4SEXLzq0N6MHNk4r//uj9zSgSObf1KQA9Ou3RF55pzjrr1THF9
kXXCqz76mZQr9PoM6sODDADN1D0LPmgnucPVJVonflKZheQwCYTyRF2Vdv4DE2Vo
mvN5Z2KhW4FPhxgAO26GjLwiIfvPJGQxkz2A/ED1O0nvs7KYK4PA1qTGcEqWY6Sa
ygxJ9W3bsbkzzWk9lyghkjsFxd67ZdV6Qty5Qjn/Hg+oV53y5leiQ0Syj+/yeHuR
w7qT0RjYWqhPS8mJKG+t2CXmP3OD1ED5BzrwX8Yu/sQlRfZIbrjjfvHkvFpzPsFO
a/MCjHnUS7kmaRwAKA4wCB0klWgdtxgWb+xQBHL2NBOfRC6TyGUYcB35KYQyhV7d
Ypv0/tufdtGcPB5ylqfgXhmMpR+BBle1F+ZZyXGjlADk3KALWzmuIPsZs3mVSGwp
w67mxAMgnPRGwDtNG4JF/F/rAMBciu0TM5LD730EoJosyoKpu9Gt/Euudq3tOfcn
D8SlYtalhJDKEo4sxwGCX9c1Dc2vXaTXtJIqCOoiSl20aTk8RezymWaOEeZa8pOA
LPs9sMtp079FRI2gQFXUP1ghtC34t3frtQaC4mfbuzBRtRqqoXJQhHE13rFB8oZU
hs7g9hLBdlkxAxqJ+hucxF23BramC7/IrDl9TefRrBO60PuTQR1TOOPZlaoIKNu9
KacoSfvf4/M/hOg+27HnKBeZAQKhgq5UK9fSXiAOXuaMhrwjHWxU0Ktl5NDUkda8
4KngWiZXW+KjggqmEiMZfGk6CLdm+UYuBsPS+5OS596xru4NTlorlwVoKaOt8djv
YPFvy4+SuFo5kgZcus8uK/4VZUN8cyDwNbNxp7W9m7+iKMLK4arlAijpUeRRyP+o
7ozgBJxHCInW20qfZFnbZDlPqU+LZ56pRbJxjcppX6mBxH5+3nuLQhf+wwzizQYv
mDvH3qqDSHvRSk0IH7V9N4b58zwHmhmB//O+4vlCkqx7f0XMeQmCcEvoLPa2Wcw+
6YZ+s9IE+C1mr8H6y4QRQIDd9dBcf9NEdW0KgUvnEtQLv9mTOC9j3p2CgQeznX5L
w252XUSj3AmyDRDsdlb8kw0ckfb2DNyWg/ILyEyccv14RZPaE9aWvW7bcjNvcg1Z
ukYmvCGNsKbacsvrG3UKWw+CnzGMuyKpkxOxW3fkyFZwFjibe9HJGIHW1nHh/jq5
XmZPmNDL8+YYWPcfvMH3CcchgvUQCazJANhhoCanMUPC/JM8gjzcBeFzfEQOBg0q
9eK3kbDSHk4oIstisoBz7kRtzhxV0UL+Ew4qbUMKqROO03PekNj9KaHtaChCyRko
RNsGuXFC4ntZsqgwFsqBZeQZPZ4KKBmRvSLBIgYDS2RSbMAh2Zn11Ykd54QjZ1Uf
euKmSXCSetXy7C+82AKhGg4NtlBqNtfkdgZ8XNt1rxkPn4BOZlYn6ai+LJHM99PT
zVDj3+GDYNbL5B6I791UP6JP78SnNERSPwdYE5qoH9LidO3Vcp8G0mECnr5aSLI0
xwEWfoR3e43/llSsoa4VMihIl9ecrHLZTCXny8IgLmJzm5Lft7bI2tkftRukuu/H
eXNmXohPZS3CE8zz5WMZWstufRzW+iV/ajxxKjU0e5aMqNfjIcx1IhDYbN1S6X3S
tyB2MxaVi8tPEhdwdeuiXGy8EsrYegtaLJf/j+MG2XT4DlA0oPw4xafFaaURwke5
v/fNc03L/92Dc8VO2oK6L58iHWN3xWW0P/0z294OldwKTRwuUZhCpZmeOf8GHe1n
4uTM+xTGC/NG8PHHbeE2DPv4aVyQSkEhIJF2d3T83Fx+GLjWCp4YxeyJpRiYziJ9
q8EzTSZKiCWBowUKOP2sQYaSJ4svZbhaTaKCLfS/hmQHnXn88hC0vEF6GAOM8NNy
Oi5tRiKlDsAvHiautqGUe/8zBggU4dH87GYwwQX1Ej0bIcVJpkAvwk95bTXJ/zxL
uA3g5ZlNB8Awhg2KelUaq6en8YVEIJsUkBkukegwW6kWIEbVxKjsvEIOczxvfQHs
eKT6RP9yvLSbFqSs/qAQisSUFBn5WOiMR0Ku/cNkK0nwFjtEMHgMOLNRMSPXVUuU
p5no0iizwDJFg1HHdprYHDPjkjYIT3DvS2n+mvNhKBx6pXiI63Wy/U2DbpSZk8ET
wbus3EoGhEiUt1esBkNHW6oqbHUWwkXvKrtYINvjoXOTezgJ+voRDZD1pVm85OCX
2cDFTIsDtnPR2/dSP486GuQatxyxIdrLjxtTWC9UokSpdVz3yYnfA2wZb4aVgiPZ
YWvvpIaifx0nlntLWKpfS5l0pq8G55p0Ad2gZ8nUQT91bmL7hoe2fpI+nD6XNj2Q
mUIRM7zIpHc9VNAoMTyQfYa954xwKIkiGXB1S2kHsxBzfKVE3uGFIhQWARKQWCwi
Nkle1xYmXWeH4p0b4KPpEwOS1/Glhh5WQWEFWShDIiEl5Ji+n9ZHFZ73ec9HTALb
H8Z/4iCL/Hs3jrJD8GnrkjxfeE3xxo5Xme1aeIjp1JYlPql5xe0LwMe4oWcs5Duz
OihAnXhKO30yU7BSRcO8DH8Io1ADigIaGWI8AE1E89IPGKAWu1hZNuCT5yL/htjJ
F8q18bluvDGhtA+MZg1AS+7X9TeF9VBNj6maiqgU6GHAPah285MlHseXXp7BGcKC
h7vdYPQ4JWzJudLMvetWD7KEni/MHBErPPPzQw8Lg47F0N2WuqkoAgkU6TBvYAv/
h48uyDWqwganI3/T7dqUBe7f8NhmRWjLPtKualfWr2Bk+OZ8tLCPIBGQjV0p7mPy
DIJB3ReXJG1dJz1RsO3iMr2yBT8XKqEQGFO6+9W6nsbtPOCwx1jmygu7V/8imkLj
9T355hypQMBxk/Y2dFoDqvWwHXJlpheGdH037Zkf+mCtTbtBdc4vaLGvxqjt0/1Z
jGjrsr0eNabiA2GE0IDjxEn9NUMJrCrqlChIoZ14BC5gR8epNIxyo1rRRw0/Xsh8
G9huy62BVtfd8xBMD5tUG7GXj1MaXSesN9a4c/DI1kpGZMHbwrgO4nyTl08VjzUQ
aUqAL49hOCU4ur7NjzloWfBjrYWK4Sq00I6az6/XQO0QZvOUDfq3MBC5xquoxipW
NiOBtYTNbgKGlIMkdIAMAe0Ft5QP/U0DLjuvxv/YMXV36SnCOlMRTSRljBtfWvlS
+P2QySq17iZko1IkRq4sLXjJOdszdopr3PWXtYOs3c4BuyXc1lzDATT6ge12ReEj
wlGiPHU2Q73Y+pC5FqEGqgZuMiMc5XJutyt9HNOzT0hAS8kExgtUF5j/GawOP4VA
H5fV91u1F8I3AY2WmMqvGHixLquQLpIuEJNfie+vVCPAxauRtpMSDG/1a98rgXXw
F5f0b9FPsyH/aXlGIN7D1Hve/+MmsJc19Yxm+gvCCuJPnpZJnlHyOoUrxbQsrIFu
3dii88LQBVGA4RIb6L55QaQq95fNCgYVEEzs5c+sN0Ab9NtgIOjP4CaCflHIN8i4
b/5/FN7JJPNOd827w6c0MrxrVkAJKszDN0gL0ERGfZeicYFFd3Dd9aQ8x8Y8cDy9
4Lr/el13WJngu4uvLDQtduP6EwdY2GMjWNzMx/I4hH8w3p1LoFZBiK0fAJlHAbv6
wMZQSFKUspEVKqFyEJcKOURoxHOLyu7wxTBCh7SQdSFwctdf4P7i2C0kOQxid1eS
1szjTveS4Ahjevdgdzz1HDNzGdNGq9TdBSJAIpCG0T3wDzBV26nEjyxItU7AHsNZ
Api/hY4sD2wBffnBLsVt/Dy49HV32U0m8YoKAXqwoR5MgGcrRh2PlXjGx6dudkIK
HNo0nRtATpKN3I/JY3Lh+KBPS2aUCdE+oGN55nPIIumhBdxf488BpMwB2CrYhjL5
sKc2GdOqo7xdVCJu0eY655Iw8ZafRKftb4MEQ6luAsIfKnhjwt4fyg8eCwKBnP8a
AMlwxtFsb/DpH411dHPVNsbrzA9lTiNhP9U/cN/LXS1PPoahS5gTvON0WzU3kKUP
uAcOf/Xx8O0wS7gERVYjVBR4RH3d4/bJidAVSHOb2zYLrZ551TAHuWOORvxkuXt3
iIVLcdLuWJD8IvZ9ZYKLkdrn+oXf9+thM27xG+T4u0gy5QRSZSf8fRzyjAzeEZw+
fpjY6lqOHRBx7rjNu2ry8fiJyHsxa3scazyvETz/5Yr7chDrS+wqNhb/TNUlqIZJ
TbAcsuJBR8CGFRJqOxVCIhDazvoOBLLOs8mUBz0S4thW2AlsuTiDO8YVWhN1T8+Q
gtU4+KJ9GQuzRILssgmHtPWwUEki5B5ZBPum0P3swD7Yga9iIJH2kY9jZMU5bBvW
8b4JmdNgrhpkLbrjD8WZZ3SDxniCdceM53YUBG5tKGSEH3ILvUIcR23mW0KoztI8
ZRXJGFaj6NklIeeey+imhKm0jpC4fn/RX0BIdvgAw+IGEzeFXh6rMpctHQQ2Puj3
eRxcgRbhF1feTiiayqkQU54qe78BVaM5iWt88dRyROWhGQNUdArkVSjd1xazkT0s
TYUhXvWxiMuulSrL2FLLH8soK5BDza7UHNn0W5jJTJiFQ/zI8+SuOs9LqzZlfvnC
w7plYDghR5b1c8fwR67875AzVhwxW0+XHGzKmczZb5QnX9gypbDvPVrA2I9p/+8q
im6Og+5WV2Vpss71C/8+bh9mLxrHbVauyMFCtLMNccr1VlWHN1l/eHmk1wkMG6Y4
MPpbESAaVyRgPMt7zB/u40/NNJ8VdDLUwTw216X9/7jM+L2GRBBz3CVQmkrSAgq9
ko1zzdf3LTURoIpTIsv9DvkEtGEByrCNDDLMQuyLtq0ekwkq3sENlJz4kULoKNej
byI0LTXjB5i5WRmkdVn8f0cmMV87k/sUT5N+/KzCWtwuQPnwZ+Rr5IvW7yR/QIjI
altA5X9lEq69KsHTnrYJYdRuvC9SLqMaNkSxp6AvFYoobIYBmpUpqsOIIMbsYACm
nPbnnZ8knpThiSPu1p6xA6PESkWU95JxLU36s/NXPEwLcMqzuNCUS824kZurZ5wi
OMtw7Z9LW2tfkF6lHeipEyIeJTUpLHk1Q9aoVlcUEGqHYOfG6O/KxF1H0SJ+rAM7
IzTRd/sB/hGFDjM/MkR10Y8KHWipmUOUL8O+cVBVPsf49cm0xlRSNm9evqdyrcGK
S9Bm/ItwQDOjeh/KZhWTtJ7EJdP6Xc34gPw+90w80cTTENYsMt5TTbH0TsYAysm3
DCmACGOMkyhn7GZU5xIase510wQ5z9T7mnL5EajON+iJ5rJ3re6tSenc7E3AZZnE
pKL0eEOxC33aGQswHeJSsZ2IfEiUZ0IX/KYEwv0jkbklXJGxqqiEUu5hZoXymPeY
pHyPEmKtuUbiSL9mAwi72P7kFSZRpfiYUm2Hxv1kCoMPUYedwMErnj/fj2R9jhPy
5fV41HIQFvZxg1NLsQhczkKODSUiDrJA6OyW51Msf/CHDEpCCSHLI6PhOPTHmU9j
RjycjZM+64T9higWobbaZ7LuTjmK/Kph9eTkniJMcygtocbjtFoXRSHcp0v7wOD7
T8Se3oB2pd61drZtqvHyPHYwA+kTFjp6qw4FSOZxcpz5GsFmWqAK8YerBftmg3Z0
t9ZOd6QeqGlkemPMHbFCNHuSfkxHnjfgw1Rn36B9PE/QeRFIjnNncdaVtbRkSoUR
8rhxB0EC35HRcMKm9GhHGNlqCBK5Uz+vUvczY5TdcqXqBJeDSc5IpzqQTqg9UV09
VGRZe9a0ciBuNs8vVOFwKuzHk/Ymd0yUI9jbpyMWe8SCpQ6L9vygFqurPpWNq2MF
aFmj0Xa2FSA5P68SXIF7mV1JHrw87pWf1CBDVsHtloFerDe5Gaj8IidSXEK7vYjY
0RMzvQTogyRrpDLT1Ycdx2j6noFM5yfBPfsOr5SMFF0vTDq7+igbUB282puxoUjG
JoKBT5PAgL7rB6fHcAGlI10Ia7RaioXrEgLSOgnTdzkt+qE43MKKXq7cDzrzAG9f
DT4CDfF8XGXoGrJYSqimTKYGwxjYl5eY0zqSXA66CjBp38thI0EraknCOsh64WL6
joja5+E0Ao210QpGc5NhYldSHeOIGEWzo+sO389SyBYo6vNGXNHBGZabQOeNZXab
hUc7Z6c48Ay/nd96jI2kpkE6TtfsMXUx8KYtLO9b9kti2UHEIZh6I3sqWQw59bZC
sPR+Sg23IAdyWeyUPTF6jk4zFSQIho+0gdSTERLK80DbPT3kg4HI5Cqrm7gJosSd
X0W5DWDjyGxR8CZWxZa7n3ISq1wEHGYjLEnyCoAdY2Z4LDNi1TwetfPUkXTLhMxZ
ockuR+KozrzfZ9x5z2IpVLxfZNppnU701/4dtzBhGxdKmnTdG9s4JnAhRReG50cM
0DTLYfs23RyxV8yDLGgczFYig78Er1+4fk8aHlvdM/F8PIMAsXDfyxnRIn9CHdVX
2jLRxqlt6te6gFwE9gkF+DOONdfCbzCNxUWiOhhJwElEXV+wnQHXsJMy2kDcX8I0
D7qLzC8aGDg0ZK0zJbN8hB/6KGUIxUqYQtxBwxPXuQ6hnz4sLSsbAgVPgLjyd++h
7/Q4I/v5/oYTjdFcv8Wz3B8XmSUp4nEHb2b4AjWhG45fdbtWbOAYZ4SSS2lTZ/QZ
KetmeHsomAkSS0RF/O+f11YGSkJ07mi+Ka373eTPGQPtegDxrcrX5pgFfQoJ+jz8
obvCwZ1bCT+b7nIaTcE78IZhoGmjAu8ZxL0te9GGV8nah4QyCm9g02vfqmXHkKKD
/wK8P/hX/rs8k9Y2Clhif0MQD2WQ8z52uYi2iLCl1k3EMar1EyfPQEWmO+zidP6T
AnNWZ6VP8G78O65Tzeu+NH0R4TXHaoC5+cyIelYLNKd1YKvbQhMEtK2GLwg5gyhq
uKRy/9g8HRrEMsRmXrj133xOWGHjAXorRhVN29HTJqUncHQLK74dLjTlaR04IyFX
lm2KOJZRG3V1FBBQHED8Dxff61ekn9xA3nrdNGKHVkLlWkVX9AH/C4PLl1V1rpax
ZwLkim4YC1VFOa21+9tQU3FMPnYS9f88WfGo/pYDV7pjsYRQI6oYowc9nee+UT5D
lPr/LcMjWiZv406UoR+Jwbjv09VwPLdKgfWPUG4sS8tqZQ4a/mMtO3irtdX3cAeY
IlzkvoYEl7BFES8CWWx2w0A+J/4Oknji9j3UVjO3Nmmje58CtP9jVd+4Nek0Hh8E
1wU8lNc3fpqDG6B28VsuhVArDBUc5CzNfv3c7mEW+uTpBJbM9wfCCQ1a5u/zcjtm
CsI+QE9n4KpFVfUK6lPZUQ0aqsra3Js7ucf4QXvDurM9+ALA82B/sP7g+4dLFrDo
yN8l8sjmTcS6kCGnTfw+s25I7g2pAWdjaRuOmoXmxWVkKhuBawf4hTgToEa/gy+f
rd9mTDd/piG3tGJAIC75MdKmEVgT7ulvExZ1Vjvib2DQvyH5MegGGkTHnMkOcxPX
9UFK9C9x/JrYj/azq286dTPowfHIMWp36ng1MTW7ewRisy+AuFQOuG8TwppTjZvg
XtHKjP/3RJ0IjJmxaBqiQBwjoD9dpkxkqlqmY7Ot0Pvj0eU0GrLWPkA3siBojrfy
gC7uRVCric4m/kGEgV6WSH/3c7aEl0OCbvLr+YLkyQrEJoge+IIbRw8gEBm95nAA
aFoD24OEVfnVXRCKreYR0FEnEZDOPauFgFd7hx7DvP+xQJrvKicp53OlrRieOKsG
K7uz9q4T0Qk3UgkpyqADL0rbYGgovVWODWg/qMNLrrtf6eCT/i24MPcPscCB2Q2l
pE4grb/pBmUNWY7fdfljT/7fwKd12uudd8tBTkkEVopd/n1gGCDYaAcYsosPHN1V
VjGeSHcALbULlQOaWZ54GP3OHHnaudPMr3NRDpiRuE6dLWeWRwVJgkma4NAO9JGP
P3sLAh60/RdlCPa03uTqpCB2PC4VLQLrJ2XJKbVKnjWzQZQXfL4didS4gU//S7tK
9fqt8zA0EU2TOvGoYcozzjr2LmWfxjbIu2m1DoNesq22+jnY6ftfIR1YH/J35h//
NYba3HyRI2tO/mfpu14nIRYS3YXovoj9joT0wnoP3NBa4u9SXQdZaPa+whpS4sDF
X8IimHB2je7DcWem+Usfw92YDg/OrmXZMjqIzGJpLAOI7QotGSeAtQJyLKYXbLwN
x74XlKMNwhbH4I+V6EWOrApvby0ujLa+glvAqq1KTEhPuxt0Ex6KRAj+cW9/gNX/
N7VP+5iAnPLrlLYaH8fKrwaaRRLaXmCNMs+iqJlnFNDa87XHIqPv2qqrR33Lop5W
JSStujz5sKGF9PBgn/YI5KrrKNr4pkvqDaOTGqrftV2twCmVOY2aBHMfRekzrwL6
hFNvj+q/jLvmUoJv59GMWd2v/XBNYPjgZR1tH3BRU2VWQ3o+c5T3n9wA5ru8S0Ni
+qdOhK9NxUTfVEX5hiy5CVlqfa6KMFFtkCYgSIEwCQhDI7rre4KgIwFef8mHuxRM
NqcItkCBYhuyO3jJgMPA6eGZZZM/IbHNkKgwoMX2K9AJh7MZzx82ETtd336H9sdw
1g6aVv90f979KNHhRiJXueOWhEV3DHZQ5wAwxEwRjXekRhCw6zHIFwPzvRatdI8e
0HQmYsQtZwG/ngFh3JW6Zaprxqym9WhTALJ2e41pM05Tm+2+7avDUE3Y5x6rt1DG
PDuN4vuampBgbTGjWEweSP7EMe933+c2sP1jgJrKXcmxo5rCr1hdkWu4gnoSFThs
Yl6j1ln5CV3RWza9+B2gGIwRhvuJdNxH4J7A1fXUiacyNzMeWeEgliPAeZNSxso8
qoi2ZqdBDdlItNbvF3Eb7OQOHqhTr/X8wHBnDoYvPvBJbUTWffen0scdWmmT6RGH
shilhyERILOBJI+2vuyqYA1ItuglZQmj1kBNEviQUbqij3GbBp/Hrj3VEJOw26XF
uwafgg32r6UUNPHn1oPtJ8k91tyV6TWM6zX2W3FozvA4Wez9NxzdRcd2Haew1KWa
ZkMdehwbySVEuXCFI6HtU68bHhTPxD4p0Icw/yzQ5HvteuiyKwqXlR53ZmUvAO2e
j0klerb3QAplabx8WwS62olDuy/0NR/xga89zqMV9hyvFj0dububeQxFbY/6SV/5
sAD7Pwu+Kj6G4Anbs7t2ZWrn53Oi47Ib6c1r05Irx2HknhmTeRm573oR5iVQBpdB
WFQixGEfBF1uqh80glbDwY8l+i3NZ1OMvdiv1qqnesQ8MLlWArEk7Eauj0QgKCW+
J1YQeMZIg2rrGGMsoAyFCSTIy+Ox+Jch9MxkWAz8bHfl8JqueieHUBPNDAFTi27F
S81WW5L73uUSZXbC8RGkfLJK+qvx2TJYIlDrbvOX8NXZk1Re9xz6FdKkbTtTQTK8
48Z9tH2g4XtORwDgp/uGstwys7MgjPsNZUOyHb/fuLeUacL9AXJX3wlZc35E9HGE
VZuLkRHFrn0x9lYdUt0M1CfIoYZpl+h0TsAnCY6suF6nENc33tqwu19Sv1uqn7v9
RnSWBYXL3gY3BFNXwlKI8Lxvk6m7SFYyKKVFBTIGnlgDjTCAYqnjEmduv2j270ff
v7waMkWHAi+I4jyol6IKaWzeQDvf8DBUxEtvaZPNJJdQErMi/b7+mxAzzuNrhVlB
ahDPaapk62cKF5ZEjtUgGW8V41ISy1DWQXIvaAZ7ZKti0uamF3yVhKy4H56XZt7D
01u3g2A0UaZdb1STQORX3x9jcss53xtiJDFplduKiVUwoZwQOTWuaRTZ5MLCUqHG
v+BOnHDMHUQNuEoL8fXGEztp+9GugJLwBQegBve3JzRE3huS/rA3Nr/rgZOnzof/
3mS62VsR3RgiSWXG/NOPxclonL8cl+jbL2gSXi5LkstzQ039hr5xwnFWBUWXZnRj
Pmxlc7HnQPhRSvANp+Vb+cXp3IqfVPb1l1pZz1N/8sIFpxQIOeo4AJwT7P2JJbO8
Q5iifRgpURCVMGA3aG08kFCrrnEG/DpfKJWZF7m2EJrIpWozqwy3H+mbzLXdEC67
eQ84Fs2hq9/7eQ52D15HpUWnzsyKYNUX/QqPaXlXVuNz0axthyF+qr8t5yXOt4pG
IxSIqTcx2lOeqZfFJMIHU5xTx/AEFlyM31ewGaekLf5ipmpC7tpRtJFVYzibH9no
ANidDbHUvmgb/zDNRTsYxUmJrjrxxkznRIaf85uMnRQiQEAYYCShIWL/zg4ebhFI
qTLvtGQ1XdXlKqmm/aspBO83H0C+NO9W2ONPi00krZZhWhfE5ZNBkbedk+oQCNGg
R4NEiFkLdPm8TlcxBabCVCOedaTG1Tfj/WQl2sW3eZm5ZfLaKiPEpLOHsMUyE6C7
XcPUUQsnZQYgqd1HvUP49uEZFfcqhqJoyXBs35eLCcj3wEVtkGRFmz4sYzr2286E
3RzmHjRKPrtSxFaiuwf2JoKpwE2meP20o/oQAYc4P9Z0odk4qi2yvEmF1zA+sKYg
L6v8h8PIRo/rG9hD/X5+ZDvizLjSXVa02Tl3OgnLj20VSv3AVraCkKJ+fcOmT6Eu
YRu8JdJkc5WSYdfczlfyeLgZEqsAHKGL0n31wHHB3+G+E9zetJBlwZsCDK0HfwNy
W/VUs1AzXmdsiAEZn4GtpXydr7ZlMSLSlLAoJXB3eNsCZZ9uP0UDnVdQIAjgLiWA
FXw/8NMwBiQIrraQ22GxIfcPdQPQvtlRpR3O3dSt+by0iyhJvpT847wI/P/3t/TE
+Vl3vYEWAOsH0IJn7jWwwhcm8x2SZC69Xp4ECcYqR4k1nn5VDyGeVNXGlLsxnQze
qlaUzdutufsh4KnqnrvUpn4qQkiKp7/X9JOXGZnX/hG9ABJA8Mxb51GW5iTCP9j4
xmGO1XBjS1z8/bLCD9s+kEmbsOfxH+irNoFkUXZRH+KUg0C/6zBfzufwGgF0qTuf
vyjI6DV7doQeGioW9H8IqkhMbbXRdII0EmfyOYBRtalqXusO0fW6sg4B7Mt7elSY
nmaK9gBh4bJodQbHr+CIWaZM1KLi8mf/ROlL2f//ti//o0Uy0Wo8RateJBXE0gnd
0okE4MWAuhPM2Cj5kl1lVF4DUk3SASI0qr1PKGT7KYRNpwKHeYXqVp40pEBLO1gV
CaxMA0rJYXQTYSRVW9+qpwhbGDkBh/NUqWsC9W60pL0qQMRCdc+OknQpYmk6iZy2
diUYxpSLotfzAMUoO7XyjnnrpjcZWissa+e6mdW/WbIfkRQsMHy3CGH9kvjsOF2J
R3qgJ+Ks/sQ4wzOriuVL7qU6Da8Rt/4vOE2tzF0jf4rx1XbuAleOhSgFlZCgUAXS
QYbBOIO+j2ma0OdeARl9SSOw/LBsUwuZ1I433CVIr8NmMz+k7GEmxjXhMJLPtjVW
K/qIDqCBpKMElR1S1+d9UeSRvDXBDkIpoFqgHF/DeJvMI1qukU6wqhSTQi7/mMbY
ZOfeoBiyDcXOFueKS/HtXbeJTAK+G+1de73m03DABbsfz/qpBGpOsODX0A7k8oYR
wplMOC4ZDwHzO6zkZKTgo4F//h4XT3+4txWqY/CBhAqgNtv+uKPkm3DCnc1IEcsO
fqF6A6MWHyqY0VIIbn82rlgnsJk1LwG/rOsIqHo9h35aOCrkBtx9776qo8Jh91Wi
y3bbbaxM/+AgHNtcAb9vB+zwOtF+xgj+QuLFhVoJbJ2idm6wcdLRFcf4iVEVoPD1
RUnteuBLFwdoBlnLp/9TB6MRFr5ECPK5rDNzKGs1hwlzpU9ylbEaNskRYS4fqNNQ
3KNGRIcFp6Q8UKDdB4LUy1h2UDMN8jBvareGdCizUgHULrgWLg97pmqqtIAUzzsL
ZDEUBJ3VvxOispDn3nPTGspLecHq7QYAPOtySNOSacU2idkaQogo7KdrIfDp91jP
lUfdEn+dPu2t6TT3BYUa9aPNM0Gkh3mTUyYeCkciEL9kMtXQgJJN/4lWXCFRFhk9
8WZBNLKnzzJQcSukvE80EpNS9CM9Bw4Yc23sEf1dRoMvZhzu93yQxOu1UPi4tX1h
euuP1pp25me6JvjCugSjniMdjZI9/UkWAVrHNi+2UZ6v3mSi+yTcEwYb89Mzn+22
b6W0hGjn+BOtYT6wB0NkLSYaDYnXI7b+uBOkP3tNZfNh2cFAHMUBuTxVtrz5cu2j
TLjzd+xefBd1K3PCKW1rHo/0r/E+ZB5F0t5uzXuVAms6uXOiMS7QMghjzab75/IG
Trtv6s/vobj3r5q2oCAbComZerEW+SPxfk9gUSJYXJNaZ6wBfqWQRbprm4UoFgcw
znbK0QKhkgrWPLE1Yg0cQTfiA/j/0YAJSQ7hbSUrz5W6B700oJOEaoj47yQotYwz
OBx40UnDyMh7cnlKLL72MERy0sIAYYIhuALVoRryQI5Cr9KYzwJT5pBzwDRvoCSp
piUQbBc3LpwuilS50JFbKlzdlk2VWTyd/H13YDXALmq/Rc7dkPz+io4YBEtMFvSa
NuVB3a5SytfVC6c1jnuGepe+NiyB991tq1Od6QbjXIfmnHo93uftygbGKIzl9rZG
24ViL4NOYRjFH+Hf2TIKCBDV6SSfQBayffn/Lx+a1Cvsxv/4a/7GTktX81GYhk0d
XBhcDPmNpbht+YztKKRUcm4yUKK/tnM64IA3RYCD4pvG4o3gh1TwWTr+XAVeLrGq
tHa6UVbCFF7rb2uywp/KSLrY39CZd51LSswevUEQQWO4u5xIxeDCDihVBmRfpVFk
gWh2vmlbS4jk550v8tjIyZNb8T2tvT9pOtg5O7Q3cSAygeOLb2aKHAzZ6UH+XhXJ
5sfTM6bNfkSeAKvqNrMoRDwEBJPh1/LK0hrcMlq6PFqudYxgATZeF2h470TQCvMi
BmMQHvBF1Y/QF53FRCmCei3c2Qkm7TifbCMaToOPcbcUx49LyVsWqniJ8Ympttzk
i1ymGXQYlscohgWpMd/a1uoFWzew5yLCMGyj3kjX97dQ00JpyoVPWhAWrbG3V01C
EjPq9alzLczza6Uj8HeyTqNgZhcKBSp6W+JyPZf/AryCsSDgceJJb8Ti7c50pUVk
KQuxPtw+NKuyT+iFRT9qbtSBzOc6h8wy655vu2SqxDk98NGK9devHqIkesI3QYlw
2J024taiwCxvdnCshFmClG2w6IO6Sy1yQzis6iHi6Bj/AqvMSRc0Kl4fjwPulW0V
6hSqIMTIAX98hrHqTUS6deqwCGQXAko71+Uj0cEZWfRJfqoX6nSTfi7SaVzcu0kO
F56FITV2keR6+rm8UEauhGVPxPTnr9Eqx+PletrBDQvrE28vhkyv5yf7Tvt/mYWp
0kC9ZPwOLp+Hz0DojrIld0YtvuNn3OgGC/XfyxYARnIUOdzogxZz6efCZsbZX2Jg
I4L2OXlMrt7iYjYxio38Oqd81BbomHqA6ph3Ft3CBq1iTz/AeI0dTaHI18Tvdklo
VM7cp3ks3JzOqNrG4ISrj54k40PMaL9DCHLIjlvEGhfuiRwCVWnayZ4JEZdRX5cE
u91ZcoEx5EOIBC9Gsf9FPEueyWwCmWSaSrnPCWwVDDedGOHJvk5L4ki/7GzSKPGX
hYws7qL9NyABQbyBTTMrRtfxVEHTBSwUj4NZENgcAfKni6ijFHls5g2aiC4S6kAR
5Jjo4aJe33RgpTnquLiNAjU8s3ecNhitGwy/sL1WF+Tngrga4q0nkJEk/lIDv9fa
VHnjxiACuDD0AwEOWDutJ3dayOdRWyAKkEDufpLss4e4uexlHZhMQRE0ah5XT88O
cgB8SNiLiyIn1m2RexVeaP69CYb1OpF/thumTH2Ub+YVl2sGoKB4VrWnFFnt4gyf
0EcLZpK7KWi1egcF4CIuejCO0Zw7sBXYzV70DGmZMuW5bOIwsYvqASIDX3EpI6Lx
w2uDOsDgPtmtffMm2GwbseN7FW+5gRHtZN6Xf3a4/1cpzzUZ+0pphAPjtZ1ZVaZl
FefjFk3wVbq1vl0CtmAvZ2WDgrlRfrYH1dIc4DjaTW09JBfpk4RzcGR7lOpv5C0u
Wg+sTMGRlZUA4qn5K0wPRts67iOAOyrSfXkxwziSsooOWwEQTM5+lMoL1K5d8YqW
WSbG5xRU8HYmAb5h8a5y3BlQTruUUolX19DnAuKTBZKuBNdXlYvZHiCcJTwvA/hK
Tx8iv+XOvYc4dBA98ovmTd+XdByNWS4H27I1CXpz8mhHkCrVRdkAHp/0fUyhN74p
ppAS7bZQHXgV4r6vMW7ZIqsJuPg6QKoL3A4eQtJ6lmwaZrOTfr97JvD38ZYh7mWy
2iWPImuPUI4NBEurvW16hVuRfJkrOXd9pCTAo21dr0sRbZInZ6khiOA5XxT2DR5T
6CxJj1S0TmWUs3Qgygc+EAHCSk/i4MB/MH6tC9dSElIJ/g7Cseci+7jHjWVJbXR3
9FjQ92/gAOMsqe4uoYpYvsyFj6/kUR65Rmv95bVXdllvfR64zbq9WZLWUXobYFn9
mNkb/rnjrxQsCFlPAM8z/63CU0qx79ic8ulKlDcrLisRO87sN/xv5nQwKLd4ndZD
4Kvs9sktoBywOmdJP1y7GaPyo+6qWkB1yTqKhDo/A5arh2fIbAgAF47ZYXL/RD8R
/QHa6L5BNhXp7RtIJLgx6q8EwtRHlEMH24fFz+85vP7lVCrBZs7WoIdK1MBdt7cl
oFKOMPwS5hV4cZqAvQLeWJZU+GOt6FEEdEj6uSQ/d1y3xLTe/thUWfR1KCkTKSyg
GiwpdZwOQQEZcRPPl6QDug9Odw0DfGoQNrqpGq0rola366PO6jUHWTCYtmGX/tmQ
NHH7BOI8KDdweALA+ua1iPekU3kgBFwDQpTypOqlJsz4K/xpMx51AR7Xf/jA5Lmq
ObidGE+n8W4yNDti7WN/rRKlk77bg1eLZYiyGFh/XH99m5WntnL+F8llqwR2Dn0E
7h14Il7L6mLGiabXMMGfkR7ThQ7nNHWaQqBCMDlyniaGXA4jikskG/mT+scW6TqD
3Seua+OX7GhopolbZVm815xYKAdhX0z976Cd4xpNzvjhRkp7fYgijV3D3Fn+wgT+
tgpFdpufdLmTAxFa17fcGG4lkHL2Mj+SzFN5GbaW3++A9L9sjFMOFiizFupBOa5T
5j3PUxSG4nZyfZ2QbeaJhxUod4SgzRCFpr/PDpwuzZ/5qR0Wi7imUcTKgCORZNsI
e3/SztHRn1m0ICEZuYi3XFpvMbzX/qX+Jc4HK+VrCG/L0YicpA3/oTz15y6ep2pY
pd8xhqIh3nz/IyubzzP9xMiLzSvgsvL1A3a2jjCW9lfJk4i1qqoj7gn4keOSfEpP
OwNuyS2KYcvDto8wBci4uvikSw7yWHnAig4eHjNId6D8Xuw4e/0gf4VOsoIN7W/H
4ZOFakQ1ii/pXPIQDEaQTpPT40bLHBtXWoksj4bDwFq7G1n53eEZm3nLNiv7ZZ06
99pRktd5XG+gkD2okMA46iqhws0/E+paFV/1k8OCvtwkYP5koxRS66XIhhEyabKT
WSaRHp2J3O8bkLast2284AtI1QDV8Gc86/f9IHZH8eud3OaC6WwXyjJSkaGaVkBh
VClZSpXCGvI+2X4bRHrxuzx7hLjnVu2EX8Elxt6OkglSFAq7eJQF6J3Aa9Eks0yU
5j9rUtXPh6faIC6DilMvWCXZ9S+lX+bz0hKRfyBlzrnPJhcqy2pxBlrBVP+2QdPO
V5WSouDP6H0Wp3u5qwoWS4N3Ua4GPcNv5uu99mi6uUGhDSqUiLLDwp2MvCQ8DPIx
QUr3vKsuLB0R3lK5FCp0c47sTIuOvNmJOn/iX9aCDq+Bw7dJjLP+cON0EkZuj6H4
1plckrRHY0mPNmdmIxaQOUDcSgMk6gd2brW+//p0eNLle9f36pRa5bvqiMX4zOsu
eUZ7NVrxzEbJ+FjfoqZTxqwQsWyrcTE8Fg3qN1JoPf9NPCS0d2I2LqgfUytGUd2Z
NSClgJZ0xc2ssCIMly2/J2HU29q2zTb7Nyb0glTjgzLY6B13QuWKWCToaa1R/QgV
rburWfs3kHWwweTOWGZfTT4NLZJXr1spN5gKFC8WxHRFgACoLI5C4gBSDZ7y7DMO
jkN+IVU2TbKi1tk2Jiw4JLJUNYLMvnX/LH7mb1AoDghiv1SEYtQ85eP6mlQ+MnsT
Ffj9fuxpRjPOAK4l1NeT3G/vkaEl3XwEHA06dFtYowmtxXxmO7Gum/MLj7JWOQ7N
HqxcmXlyzmpLQWjYmEBpGEKRb4c66IYzL7wv1lP28g00wC7Q9+N91dwmivYKDLsp
xeNmltmcSoz+i+/K2z5qRRI/ak7w7bdy6RL0YoUL7a2lkb3ihqtMO3lZ7Ggmkjq7
UjU+p3Ko3i87qYKpvtxMBjr9JdFFO3uDQZxJjxs0ytem5zs/VsjnAUe6/Ysrqi0+
ZvHpAPLXfUdzncktPIoyg3AHTqe5BM/ozYIiCmX5/G36uj/PsBtRuTvs+FRuh6Og
lbm4Cf3VIeX2lZn6PTH/JyqgL6Wxi/VXBBGUgjt0Bolv2UuifPStro6UyGyNcV3Q
Ge5zVLcfxEnme4CfVdj5g1kEjHUHT3hqj4eSYTfMkOVJ0lLwpl26geuaVbPVqbnB
LoO57FASWLvjNnOYjSO/rTADEWGeZDrMMC81NP7HTDqumaGciazGZJZvdJ7rOTvL
2YzTZqc0vmSFtK3TvhzsOjRR3TrUcokp2PQAYjzw5fzbk/BwzkAe+F94jAVifO+M
pH4ToIg3q80FgEs7TwRlCqYQjZ7tiBBXYj1krAjJ6Dhps+6A7HRrIxPRSVfwGc26
c6OKO/xDf2yTDcxsF4sL4VTqAG9FbaLPngO15t37X3DZN6LPjUUsuS9qZTBT0/zG
FYltsY6UwpYEqJblUBmD0WJvesbdJM7dxaNGg6CqBkh1wLIglJb1SHun3nOVXweP
srZQ7hygHspqHDTEvtK/CzQI6FV3r4oVOqFeYzndYZoVvFNGFRZpisoe1U9C9KcA
v1MlAWkZhzfGA4+moZF6ZXSamfVt58mls0TM6RYsq3H8L/KyhwgqP/1wgXmRioyc
DARRVbBNdrA5+sE+PxgIbQRPHIH1Zxy1ADKe1p/ZiKUZJsGE9U43AFCfPXLRAVbc
3w4T/vxBIJY2GafOcU5l1XkkuL+ukBvDMUWg0KIeWLb93i+ce6sCDrvb+Psxyk+c
emBaUHwjkB5/3eX2i2doQu9E30jh/q4HNLoTJjMTq5ACwrga0Hi4YZPPnq7h/0KM
w1vBiuSYa1Dhap3KhvKISnQBYc0k1z7S3BzjHp5oGpja7l/BRdRjkUJ0qKPwewBj
PNHkwrdqAIec7OMMXXEm2BTaBnjvIMLmiioaKrLBE7k5FVGAUI2AoejiXx6yua8q
nwVv3krtWVN6smudz2a1m3Q1aQRkh0soWPty09b2LF7xb7QD4KB+ee5BdTBwg9F4
tTUn8wA60zkUIM/8TFQcbt2P1wh5mOpX7x1pODu8g5Ur7Lrx8fuEkuy3XSksQPS9
t30vgws/tTXHQOK1CaFVMxZ6ADIX4WmNorI0msoEEmGe+49hXE3hvl2kamHV+9iG
xn9JeBepdyawC4ow82HuCqXGAM1Xu1koMir4S/pwT9Lw9ZbSK5PSGSVH76byEMnG
bxoTgIZIbzL1jUrmiNELY45bUNguyvwZC69o+NdPlgHPCOgLigZ1eH7YPP2nuSSX
4iyfgY+nZ3yg+OEBa8QaxKOz0uD7AEKnU4uv+0QiwoKDbXjnpFY01UOoHYmJMeMS
+Y9rLJ2Zgf7iXYBUA+lPJ2yyeBtMHDklP5M39QKijh2lmJpveg4QSAWY5M1BbOsW
5RVO54k5Zi6PVt/je+LGkL8U+F8ynlqdrna+Ovj/qKoteF+uIz+plE5aUezG2IVC
23gDukzYVw66IW6wYDnMPWBW2P1JFleALVW9S5GBonF5fR5kMdqsKnexnqf5v9x7
5V8R5JRGrXyg+ZVFyig1mFA9X4D02JR/b58y5C3K73WbQB3zQgpZz9EM8J9qB/A1
w7PRp3OcQxKO0bK9h+wfWpiNpLUegz3k+cgFHObe+5yUPpZYV9ne3aaNNQW8w8T4
HB43cgG2m0FsNyCPOuwnWG1z9y7SPsaaWPo+KAdflebda/ZE0oYbUESD8LcJz14d
Kp7elCODFPkYCI3dE8DkOLr//n9wO+F3e5HtWyL1l+hZkxWdSUl30xIgBeBHsCsR
H2Nyu4Hv6llW+dK9RGkEu/D55/YNSd1DygBClsP41FiicEoxTuNAYLETs9hQ4su/
kOiRmr+qZT260sjOd+1eEQ31nRFtGaM7gn0S542jfjNMox79reMD+JogHATEedZ3
YEDJaJRPVu4h501X0E+PEitkAIFTCRU/quL3wMGAkCE+sr73BWWhMpotmJw/Sqrd
AzeTSr5zRtAdLsdMH9n09EZNaGFRYxiKqDOHqD+XoLcU9wBTPMn3enKntE8eH0rD
o+51jA0hxLddr8SqjRcIkhUmPdFe/CpyMhRN4aTdBdkMbi5a+86GGvj63awf4dRI
ASTpbJqQp5YhRLMujTvqFLBc3f2hCsZSJ+GqecYdnGKdY26MPTF/XSovOkjJcbYf
8vLVgj2MQXpMsv2XV2Y1Fys5EKvJqDn7BjY1c1hqo7ujXtQdDlpwl40yK+Jxs+ws
qySEPOE3701+oSPdW1gprjdCy71kdudYFAfpDEilLjyP1BEdaIHeM7UXw4UV4daC
/4rh3hDjNCHRUqpS2cPoHfYuZohxu8/bNNTiFUiTP0tg3TqUcQ5+9gYa85ZDfQnp
R2HNxq5SI+12FTW5cP1tBfqSk3cAe6NfmzLFWHLAVHei0+16M75D2buS6ZZpEqOl
gzNBfLDI7xCXC/f0qc+jerDqSvmdCFfEsn3zkmmEZYjlwW4KHa6RJosZng1zFc8p
HKZPudfF/xxD5kt5DIlTa2DMxvepsPvGH3mWmwwUqq3rff08akcmrewXxxy7CHFT
OtuGEV9e1ZRbFmm0DkL8FzLHC2bjzEkN/rBGkYGvg1KOjfTPFRTOKy/ju6RCzTbo
WeLB+0Utz1TLtomxS1UuyUtXGnKK81mMd93l+LZ6aS2Z4Ysa9lAIQkTdp5bO/0mb
/reAEYaQcRiwjlgeG7/+EraLLtC+R8kF13qcLhb9vq+zBYyeUFzl3k0celjvXvqA
INupMfvg/g86sTANeW1kNVDSTuvef1zS3vz/wtRGXj9Ao0JgcSFd/3jx/CPn/Bdx
viv+FvN7MlKPtFeJjJzpm0BMvPmrdzQJYi6/ySeb5OIhLmgXEXGGIrhBZwyFgb9V
qOf3VyCioXqn3w8qJk1U6FsSYw239Ki4CluGJ/Ovl0Gzc1huNwQ5v/qfHG8babzK
pSet0U6qd6J/Z7WJxUsCqgHs6TQiXrtWFiXq9srR+UYGxugUau9rIUHWckNz6wEt
cvKMQWiIY1ed6KnKs35WkLhST8x54TfixC2ocN1uChgYfwICRDqX+xb53L0CO3Lm
ZvzG4244A8CrCWruMrzOhQuTycIKUD0qecV3ecjk9qgAFB3snfCL4nS6L+ABIAw+
zISJIx+18F4IhD4WePxW+7tWZSF9whF6D8ughMZ7yBKqbLh8+yOgnfecNf7kcDku
tXlbr3aCaxeLNd/f3uJq1WMbg55vw8gudI6Z5VwK9rBE7Bbnc3kyDySzsmZRgCVq
nD0DcC9/IyznXkJN8NhN8XFrL423ZYfSw48H+snVxLOvSDKeYKXB+5nMST3ePbRl
yKnKSnyLCyNA4sIBUgOfL/7ntBOtnMpSxX2vG5B0Ha9xV3mRGsXncN05ZjLqP1Zx
aBQdsfjN+at/r3/uFlVhimSw/NFK92ftcNvqG1ZwGV5N9cgacOE4i3MJJU2TZlnW
Zh3uhQxsbEXd/JOhiIR015UGLlQ30K3UIhResezyvGQLB7wMdDaQ21gtQ2tYNaRN
dE+e7G7U5OvZs+aetNQDh7ec/7WJ5d9P0DuDOZUCTUHv8nAqrJ43CopoVM3SkGPE
xnUpSpu0tKc36q3iKxm8jCrhb6Z5n4yuLI0XIJ6D6BTELJVZLl/FYbz2JA6BRJa4
D9S87FomY1ry+PTBoLwdOIiCoLAUGM0DlC+Q8LcJCtClH5Lem1+MUJXNGBqkv0O8
ZIt4NelWa6g84ow03jItXXsLujZvXKfGLm3Gye1JORus0X4VTkCt7V5HrmFO+sZA
If3qIweYZcIpDy/A4IoBeBr/50n/3hTVYUSIkaQRcQi0Ct4vMz3rq6wkffpWIQWX
GuY50O2z0DGS6KdQq6OsYY7ov+osxNdBTAUrVC6mNFNSF8byja9hKA6EfFTgnQTY
Dvyp7wAgHdCVXc/l31QcyWzBNLMR9B7CbDdMO/8dZpJVOXvAB43oXSQSD7LDfJcu
v2W/3I0j4IOJ97C9epQJubOokcXISdAMKiuzhvGAPMVtuW+kW2gAhvfO0ACIWnbN
XnGGa1EhGu9PjV/SfHy3DktS0DhpRzAdqmWlsFIOsy/Y/bPPIF2P6uF5s1rgP2Sf
TdmbLtMCqWYYQhuxPPLYfCj+1ieg1Vr/wGsvkJBktWD6RtIHGL9JsLwhP3fUP3ug
F//H7PSwcQHx4Si5F3ShrmOmNjRQuTxsmI2iM4tt34jkzAHmUeMQoT1A+P7LYVFA
7XbeHGZPkdB7iDZcUQu6BZpaC1HOYyOw+8lnvOX8+1CyM8y6+5BLYzRBDAg1MOPW
lP1XaBOEuJ65qFWpHNw47wbkKDPssXbgQn30rGo591gh3XlesRsBHvhw+bmjuWka
T/P/cCtJ7ufaJGLLh6A+d4Cfec4khmfkZb25+xKll029P2+y3Os9a47kL9vRKR6O
zr1lI8bJxgXHCJQm/EAdftKZx/un/bfcCS6ywh0vwvMF0KSHOGR9ZnX24Hst/Cf6
2F6OTEsJg5SPOLNmgvrL4AhMlEcYtMm/TbqM7/O1G13RJQCFq5ObsCFmTN7pErKH
Efqi9lQg+P4w3Q6TqkkNRln9ihT75rv6sNH/ltIiU2+4nAn5jHGcEZs0hlq/gALq
WfgmSvt6w5Uyc4vOol4sdJYN/3LbYDKk+KwxW1kJNGf6mF9PeCKW0AgG5wVG7gjp
Ko9oc4rBnpB1ttL5xx5ndM3qW1nwlmwtTGDof6RkUE4i17Fwqlee5xQvly+4ztTw
6v8et44eSQhO/vmTzBj1YMes0+H2GfZwzmeeLx5CBEzhLNyuvW2FaEy6R+nmGk6G
+oG/QdcjYSTCVZw/LQHe3E6J3ZTIhbQE8B6JoQinl7pCeIAcm3QcTWcLrBYuGgEI
GqXNDOI9tDVrex1L3+hbOmCiTkHqA0dl6k+b6ZfR8mXyLv8tA21yWLyFHRAACLzA
tSVh6OJlklG/75o4T+obfV9ym/YI3VSLQVVyiJD3TnMi2wAcTVWhoYRUFEeCLh7r
M9vsv9orM9Vdvs2sk9DkBawGvezGr9uXVrQIA6NFOHXlX+4f2RLxiR5CRmwaSoAo
Tk6uXqBWIIFS5kORa/4qxqCh+Jat4HBj9sz4AND44eICNpfev2cps01W3Znpbp8m
yXrP2Fnx6ZLcIlBIWgozZ01L+3St4sk/92+WwHEzndIaFACip+LuBh1ocLZ9J/iG
mljTT9M3Lh8V//w/RhFpk6qM5hdyDHxUnULdhdMvk9VrjY9oI/mpjF18j0xwkwIl
+DVeuwdauxi5HyQzGVBnwKdBmonB6M0FQMZ5lhaNYmxg2QqNnvv58btz7ORtcVRs
BKmcF+4X4kYuOqqML5cGW1XVttU0Nvgu3dlkVjG+hpCR/5RbkB2nKn1B33HLrg3L
SH3gekloNIxV3eI5ArCHxFkGQFsu7taAtagFyE0MOiX43iLJwp0wriyCoxY91inN
CglFj7wX4s10Xf4eRa0vd02P4IzwtA2vdp+zunTl2mamIIoMpLKhT73U3E/P+zgJ
xrXxn5QLn7VMVQb2dVseS4V71KL+yYjKzR3ELD1OeJFGPlaBqvY/njfV1Pnc0JAD
jfMzzwIWJnYciOcQ/ovXrg/N2djJpFH8wtdzkb9/5vV9vQsGOgFiOs6Dxgz/cSs+
a+cREaLDHwGabaLSkPtZSlJ0TP9Zxw7WT2D8rZ6RLsrOncTIWnVtGlEdXgdfYyPo
QaMUnqO8Rsn6I2r2muOaVK3/IabfRoaxnGSzw5LiEzWojt1yPRRAQsrjNwdfZKik
KTyhFazb5t5Eye+TpnK5ZxE0+ga+jOAv2kxIvHwvWL+P3r2CuefOMtAw0sWexPzJ
a+nFN/+538sMAh6V8rwwe2sQFXLEj2LBh0CKmBkjmi0H/pSIleiztph6Uzmmv3Og
wj7zDRmPsiY0XHhToM0XcSYH3AJFgKeZYcv23U7MK5rKdy9NZf7zl8+MtKNYoZAs
jK89wEb3j94KKVdhUyUKTGoeszjyLXzNlV/ygfZg3nIwqzxblWg+UtAHUEfMphGi
VB3R4w2O/8JR4K82qE9OSwb71eNzlxa1NGAQcFG9h/B3Hnl4HSJg1qu7OQ8sNfqN
qM285aQwSBlFaLQcY2gvS9VDgsqmfV/myYLuYEHRfl6y4CKgypSXzY2sahCUpoNu
xSSKPrx6rA5oEyr+0bqSioaC4BH/nB2gDrfefewVAvNrjiBKbWN6htxmrF4Hxmu0
dNcvTpO2pZVpQW3Cgz/SIhVeMGe5tegdDo6w5+rB7fzxs87YfvwoixnSzkYGe+sY
DXLJmpgPv1TzJwPNmK4tc4snApffhQ7jUMnKHwRY6gOXVdTZKNp6vnhZp8uUQD5H
EEhjcbwZc9Kl+T3wXjgmD6kh5uZ+oBxB7HJhxk3Gwtoo5Q7OKCoRGIgmFXqhvRVo
thrThUyX7it2PZC2qodb7ekqkySltL7+QNWwSjmfyrwKdOAtO9Stgtfk01k9yChP
VchTaByXK6eZ16/ziVwmMYZZ2WoNsX0Ux9elknLoA/lx3nRi46/oiQl9vmm4YafS
eXGgkVNF+GpgOOeoa+FvZ0Dn3B2c6cKEHoaaks+FmvQsKwi0TgMiR4IMaevJ9Dj1
cpbvh8ziej4D9Dg7QaPKuqNt8ZyN0qHeas9DrfR6VfHw/MM26yDxxriZXUCzHQOj
5tdF4l5VmmZHwexYGf0Yp09ey2nDcIK5iSB5RjN7XqQKTU5tkgx16LdAuCVUW49u
tvzQkUdL6orUDg3eZ5XLj6JlY0xdfaz9kgPI5v1fWFzEkWSiN8mlE3Dwj5fydJFB
oEbVBPbWpKm/JvXyOeL3YwwEn7iNYXukRFp7mV5hMJufhc0+iTFxoYMpBzMh50db
S/phcLFsQUiy2A5P/nAbcxhf4SYJH2bGce85StlsQ4wsLHPzvBLPi6ADvazJR0ZM
ZZb1LaTjrXQDAmSuhrfFmi28apZRues+7dyKR2Uf6AoPGWyZNgCIbg/vnYxf+fX9
mjHXESV3ME2Bo2E52OhDaAPbAuC2C7c0ArStH/dx1MWSKXrzehArIhYOpBrdQIPT
NxJWazP6AQSTVx3c9EjrbahhF9d9hRzJnrBrtfsth3R7e+LiwCaSlk2FSBoMLEy6
mvFhLhvXkQ/Ydxi5ev/Rzz+xlnWhspprbrzypKRJ/5qAWflpilrNBO4xY5eQ/hUl
1PefyU4w1NMV3uvuWXgIW3OLD8/xONih2R3McJOOAF5OkZXBJoZaZDvF6nbdpFdp
gj0fp7vtntg6CpI21okyeEVe958sVZg/dqRONHcSZwdEjACeCv37UOLxMBxXq2ox
2XP5yC70d/DWwr8TQnYW+jAr+tWnSWtqGKJrDuEAia5eVfyaN+BYEDaQmvT6Xh2t
3QetFFU1m2Z3Qf82MCIR5LW8qLOm6Vsdxr8KT9Ylgqm2U/gBUdDLzEKj8bGo3wEK
E6rdpkR4jiPh0ahW+XxVIizqeO5/jhAitKEu2YkfcUcrppiReqPeLyP7JIMl0s2h
/nPkegQFhzhmu3XoqIm5B3reASdQPLyQ/ribcTVRHKXxecctNJCrk654HNQns4er
TgUh9E50WbnZO63obJA2UkcXdTUYtWdgX60W55Mnn5iUU5HshQkkMRHraQ06XNiK
PxdiAKe9NtVnT+QgcmXBMHcjMsXKTcEOmw/JSbVlVRPZnnN4R4TX5I6Mv/GEy/cN
BI795KemesKurD/+RuzPcXZh53YG8nQajzqWrGFdhcuHCseYBts+FO4StbQBfuoC
jOajnqB/avu1bV/JU+lLetDqdf6VYqhCRyjza1dvNy8wtwpAfqjfupBWKlR3rgqh
aAnaCJFUnnoFcGRDVIDJbbbOfo0UTVf5FFVtAZtU26LthgJ5rUyYgkTwpshZXurS
anJ/6D9jwzpoLshNGkXV2j69Q2MVo9JtRHtEPRyns6ZR/SD9iS86mUW2GbuZr9ce
EdPAg3CTk8Aesy6cd6zlptLdpKhRljqo3kiVWwAWoHwbR62XZT5nQJSGcJdqGs+m
NXVTEXNKYGtcizseqZEbQHW1rcxcn8hsMB/mhXXfXF9I4STjA/P4D0F0rMlabmmf
wZg+W5EYmJ14qhdEGcmzP2/lK2nAhY51PLU+HwXZfnzBGvUzs7Ao9xcDmIG0rChj
0ve9a3Qzv2TGL+L2pVHIAkt9vgT/SY8wXJVj/LtVVrmTuNEsQYGzjQjBreiJDLOs
k280JHQxzwNBXKM1dN6EPS3UkKk+rfLSJWo1lBBsJrqsHkfFA5mHcFpNd1+TdVQc
z4FGRSTexa1cnXd29fhlI9X9zTIGvUj0a9ZdLMFaeLVIEo6lXFCKYr61e6+pApmy
MfA29rXP8U8xe3zDjQYpYhmcK/7y/Vq2TTssEEkjPrw8jOG74owc3uEjrsOwUIE/
ptJ/JdetRNmU8VY/KFigYxiX/iZvqPkZlT1FKoUBOtUFnSLXLI+B54afrk6FC0qz
8l+o8Brt1BKykS4XP6u7lu8IL87DkR1aS9oochHmJuRpywz13XwXc3QmnV/7QkWU
x0vzqgfhjWdvjLA2qIoqdNA4mVcNm8YlydC5Ok72uJvCNXHIgXR4j5OpurcLModz
qkONTqGeX7ozHnb2EJyCT1AFH9ZS7AyZxz6Xth4iny0w2I4CxndCetmx/XNwf147
MgdAqCVVgAX7tbH9+JydpxN5L/QnOifoF6FKFCC0tufvO3tT2ClUNcNfuqj6IpQP
5DY+wlGfhFEBB1FTHQ5k/uKW95DKhdAO7fQ57iDmRVtENPtgnMl9YVOTmBitFBBa
T5+EBdvrs1O/CsTKlx+/4OMlrepcCxTGBIeN6GPbAvYNliOjLkHBlilWeLyq3FYr
h05V5KADEyI0PDVMDYbRlDPh2N/J5DWWyj/m+VYB7qJ+T+dnqavXomsK1OTKuIi6
HTx3cBWDrhE0iqFJU8cP2H61eXCesNtfrozpcOwrrT29FIS7meMBdKjKE+iPM24r
jp/8RqOwGyACQYVlRzdlx4KjkrHie6OhMLvEfEVrUPQmrNhTWjWH/99P2jjNspAV
CsRq+jrOj+98WTMiFguiMBMSQOZI9x6AUb9sk3TOW4HpNUSQK9t15lN3wm11+EtI
DJjDbNfK+r04RazIfyZlmx8WctD6s90KPWEVbaLNCSNG3uoqg83oH4AOnH/rVyJJ
6FrKB65pq9Qob4D5lQHsUnQZIsVnTqWypbirDwCG3iMq5mY8m0OyNe3VARe6xWsM
PLq43xtPOTduxGtBoeq6qjclh7Yw0488jK416IVwAbm6FwktWnyEAVvqMJTEo9Ly
TeJg6dAj+A9pucQGZlgihUg2eCd4NTEVvRAP4V10UlmZPn5hvhlb7X/dWDGKvrvd
hRcSw1N1RhnntxW8CGhWF/gfSzRNxzLP+daAPS3v2wrG0AwYtWjv5rRElTcJtTp0
XbhFBIPhH+NOvn1Bf4+Q+jkTDVgCzO2e1CPmVUTo76Cwi8JV437h6lSW0goC40qG
w4j++Vi281i87TbVQde8+pLr98aRcbi4oUjpnrhIIyQcbTLAG6VlrZ/Juz/fp2Oe
9h6dePuIqNB49HpSuRWuDRZSnydGwb9+surTLjpedLeo0m9a7eR9YPP+PK1e/MIt
Waj+QNs351EUww94f+SwR54kYfar3nzTwTCTX5fWG0il+DDNLlP6mRxfY1Mz7Ref
qfOQ0osqQDQYpd2tvNaOLd1ouPrJvQSOn5NIE3PbDRb79E3uJBgouwSqPYpBWOCu
bxL/zlNoxSLwkC7kipfmOOfftAgCncHZjTcuKNdTIByvX6Rv9+XzUlDHMZQ5q+9S
gSwSMMC8Kf1VQh2klXSsExDe9jhHnoJcOszNihi9NFoao1VUpAAyji0kekuIu5M9
d3Pv7ZPeSoz9G+VTNfvdiri28V3wuuITDHg6bQ+oMkQDj+gbmY80cqyTbLAC4nud
tJ8/QJcoK6buXxExvY8f6YXh3MIOGHNJ451q2fjD2DJQDMTupkikYV++j1rGNDE8
ZhFrrXVkl91kZyF//DYMC9u7zHx81Y2zWDYY29ExK70eUYIZmgUe5SZPlp4iuDkJ
kyIZyEWm6koZ5qSj4ZLHvdmqzjlLVNpboELQi+cIeDnaNl0awl5XDdUtXiWkUNhA
y4TrD+AlkmfQhdnaQFCMjjCv2MaVEELL7PdQNRC/ciKIso/n1sdblZ+nW3+3C2Y9
8FmT8A8wBHwBB7DnKtlgmEgGP+NckK25HTnrvhXXwKzU4zqY3ckQ+1vYmVFFq3KR
HhzzICqJJcHSn69oaqrJIEpS/TP9hoLJFPlK0OfWQghHWF81EHChl4GSCLwVwOgQ
kTmeE5juId/lfK9s5aR/p7WeEk8HidbQey+dBRjXKlc28ULBKeN464m5/SC9LXTm
CWZTj3lT1mMy0H5DKRpApNCefjsRh0Bd5M1ECk18QzTKCvUT1M4yGtORWyQA7t1t
6ZPqPMPjbZwGyx1gtXJhT17cEpMrQaOlKjFVF3O4RTv9qHZC4nhKeLmEtnyqg1Vx
YXsIXeo4B5i1QAvO2JhyVa+2DXXkY3yMwX9RlLApkgxYLlM585EHQOow1U43ztaH
eg8EK6OeIV0OiJii22NMQMfz+/3+D8bAhVoafYR7yiVypyXSqlwd0FtWEWbc9E8n
hjgCYcMCkxD4TWPyzcFqanw9y8XlDkJb+pIE3zRE5k504biFeCGOOh6eUrhpfyPC
0Jh7R9udM9IZGYZ45RG1sRHQvlj18NlYrn+ZPl1km5UheZOY1OVQWho6JDYOIrlC
10a4zzXdUSApFWOoGSewCc/srl8NOsj0ZCYPB6jaw+89lgVFtPcmj8XqkokIK2r9
dcreIC8di1OVALdnQheT81CdsAEesXWFGC4NFrrykRNgioWIhsaQ/bMCKy/4dLol
B6mAnMl7vrOuJJLotpVE/w1tQGsYJKtfjfMAmnAXAQrrmhl14lSSrZ9dVvRJxJOe
JOdZ7mdbCa9w0ijwkc2b3JjkvcD5ma1TYYai1hHnfLvRSw5Urx6FsU0WgHAL/IGp
JGQCOV0PuaifZl3gNj55nVbWzV5mZSvqx12KB/+41ZKgttRxRObQbfB25USgcHtA
l+TpdU6PdRKFAmpMzMgmlWRg3UZ1XD+7IDMEeENwxNPhOJiEJiaXW16SfBxH9K7C
vusDBFkPjAc8VtmKk1aOMpXr/FCQERI09XGO0/+DCwZ3W66wsizdETKUcdC8WBxM
ySHYeiWCTPLmX4QpMABSMdLRX9d0TRnunRTuSADBdHfnk0dvbOpdmi0QycEZDsIQ
YbagqghVi50Ywp29jkgj5aASBNrNExcgOdvpRDDYm9J6WdmhptZVQ7ql3R7IQ12C
LeJjxU+gk+76vOciMPPVPTOjfTkI9qTegkfTAmmNwVplUoJPDdtCEYqumkVu1A29
4HtR36+PlCgyJpAHwi8zI9I79iR9OIbKY4kTWAsGK90ixaJ88roqpwmlqqrOWSy2
dPPVFzRsVcXdbcgmznozJoQjqhT5St09mFOkNo4kXm/8yQd8q4udqyoh9Du5JlhK
eVy+F4rTJMehw00xg5n67ww9IdMXjkBlj8V9KNScwBoDqz4XXblQYR0UEWihY/SE
nbFunWpvxDjt0i5MX3QNd+MtcBUnsCyNbfuL+28mh/J6YBhQbdTuDW2puWzQbKUf
LotddFSufqHCR4NgmrpDWrqbQ/XthOLf3W38NPz3mD9LkXuX8m/AvxXL8iHy6FrH
oPDLVhvdnCFisesFOAonAQjtrl+X88vBgPd5kcInorpQyln+RcG13iPANmsF73LL
qV9nwR4/6bxOwFOmJCVa9Iqbd54JADjs7/X/vWp3xLxIy3CzzaoRnrRZtNrscfWV
VpqeAKS1+iUo/gT4AvNFw4dcQMUkx17/fmUHDzMjQsBLRSVzhgJr3mtghkZeRV4e
xaQGW81Lgc8fSg3TUMB5WmeI2BEOzsfWKir3xU0zDoIJkTtBtrOioXLcNZfNer+l
d39mjl3kUVsJM6W6vNuT4knAHZBch63XeIMrpJe2fDWCmkpapDMnz667z0KSYD18
lJyzprnB7D+IXDLd1pzOEbClvD4kUy6GBo//mlgBbjPybiqcHJhy1MKrukbP0ARW
i5hRE+41rfawdRbB1kYtWFiK2DmrsOg4pACzz4tTWGnqOJzlr3Ss8E2fplfFi0+8
S9OObUtXDWx+jO/pZzsOYuPMygxNobBej43NIQR1r005gN3zHIXtSvM+dbN4SwX4
h+guDLfL1Wffh/YnRGE7znaN2fTw6qAb/7EPyai8RoXnlkPm1TLr4cZPIL2veMYW
vS3TjUYtWvaWr6P2EZX/G53ADFRvAIopUBKAZLbwTvxZcVGV2xQSjOtKmcc8qnD0
Nsdl0kQK5mSg8r3KHLJj7VkiYoaGaOuWo+m/QCOngVIwaxUj0hWJsvtdhosAeMud
R2AT1Kvj529z2PZUzcsqQE8oaLsCHY8my2O+DnqyL2NPVd5H0wKGKe9v7sHU/kNW
QvGZ+Sy2waEMz1hepluRRKZNyXPotwM4MX7CD4BHE7R1KcxLT62pmpocdpD2CWbW
v9DiwCusxpu2DI/W/YnMDwO219ZHovCv5JCMz6X2HxRuY8WlbpzyV9j0oAhreDSN
8Yc4bRyHsAHS7wgNeMv/7/FIOr1Q2euw6q4Q8QM+cSAQBDdY+UOV/eudv87Y/c/M
/6IJTYQ6jwQlFoekX5/QPGR21sjc+rc/u9nuHxs54O7dSX2PIzEZ980dHs81Upxt
GXE8XhWfr82YvlpV9sXLWRdvuUU2XGq3GM/xEQmz7y2Se6sprOCUyDGEfRQbR3ty
SKq8Br1fuH/tZm5bmv2oqyvlv7P56MTyyNln6yj5gWn6xBwf5wxUiBO92DvhrEz8
frKOcWn7O+6+vlnX9LyXTei8g86xOaApblVaItVyRFVB+ndf0vc+4/oYMPLcZo3j
cVXRJQx97Jstf0Zre3iNZaHI5HS3w8jSXBY+fSX0z7S0FE6Tq4WgvCPKgjt8VvNP
13OCWJKIvLydaXTj0PWqrEv45+RsglME0YHWPSxdEcJTvFgq8dVtQErqbzHe25xi
lFyMihyHd5HPHEwCPKz9dgjYuYd2F4nrzOpzl9HAAWvWr9yX1x6SIrzdP58CXmkw
KBDT15b1e93xJ1lw68xb2quPeVSbF4Fa0TVjBTwso37CwMrmPq6UKwEw6STpRPeS
gFNCt6sriGXAJdsxKTHjlCrC+G3NER8wljh/kz+oZT/p2RH74tipsjhRCf6cRTHD
3Opdd0bSiWFyIKiGEcGYuLu30w8yw4Q6lu1ild3ANap2ccCJLBAFWlJ/x1uzswQT
pDToi13RzET8wxcvz1OnN5lVUZIavbQhR4LYjbd4Xz9VtlLrpBk/QJjUyeQxNrne
haRCerKaUmb70or1e5Q5sSfvDSPiqrULdWaIT43e7GfFEjfh5+gz5+nP5hdSGDis
/R0B0GzcVXmQVop2rO86poi4ioHAOkR7ykvCQonRf24aJP+z6Ta0eZJ7JQRXsYeE
cFZgIA8ROzh4XAkghOAChIe2cUIfpEdBz8FiH45HZZ4bEpmiAB3cXb+jJxQORSHu
TlpJ+UU5Cfl42PJpubF5IFJdupP2rpi3aEr1QYyWJyqN/S3zcdyM/AOIMiFXsGgE
sEeeXrMNqSJ151aEpk4Qeo8oqvyjkM1SJIByJyygo125+ggHaF9F3/EmkqIGWhv6
vlo+8Qj5OmjKGvbEnZVG3FvlQ0FkR0mbNvZzWLT7ciUrh2wFo0BvGXFExsSbcHKt
ny0tuJGugsLhCkm+rJMi4ydMDbeNBFNwGqpFMIJOri492mNTggcxeNb+QqdJbnsn
ocsV9IPtUZ4Fl84CouEdd4CnqWXtMgz47yMR1JJ21f4gaujju+WyO4qX2w8z6e5s
PHD92ClO9u4m+T8D/+XeBlz3C1S5flPC2FaEwqoAQGNWPRt9iBBVu1LgOLhMweig
r92XS41Rl6eKAFkXaCSq8VY5l+rHSfDeQ0ar1LbtYUuOpebEo8uJAj95IqSopA5h
TXlb0SIqmg0Yrjx8YhYMfEXN+wPwC3BalPlC+UkSPKWuFG7NIGS0M0hA2lpd+bqd
BRXsY+fHve+KhzDn5ZGKS70k6uvKrpv7ji3Iy/pBKxnbz9G7s0jVUN85tAddWM0U
w8I9s3rL4xwj+3rsPLFA0aSddIZgkBabY/PuVA4RHUAqcmJ7GfWz5UkisCQ9Zu3I
h7y51vEVXl8n1edXiNVr4kifTa7HxwU6Gd3ooAbjHIgSJP19gpScAiQs8BG9QWsL
kBJqekL+J4jkWlmP1q/2aFdOro7OSnT6KxGDyytbnhyYWOtIN8Iio9DdBQZenbz8
zK2Xp/hs7cmP3FaOJlWXdKFc6BZ6wWKKZq/SVaIIKDFcnC+OLNdcyKx/gPj/pjru
j+jiEepC3pQiUuMMnY8UytN2fh5PzVJxl3DqnhycldHxkWpPIrHP2Y6FqNAXycS/
Vac2kmcTgJy9IeY91x/8ORIHbW5XpxaFFTL1uQkhGe1fqNyp9pWAp38sD6/fZo+P
pb0t+Eihq+hnmXuuKa7tYlEcIeS5ZOLjMeXZzYl5kCFbrTD88XgfFRLbtsKvnYgS
EzNmXUrS10faebr8+uxC7hvyavX+3/zFaRQB0eQ/F3W+sxYKtsY4q7TuUptAvyMK
QwDzpf4lNXGxh/lsBJN0usERIh/m3SYHa/ku9KqvoADw+1gKJ2m8uowr0qhUbxJa
QrJ7oRHq3ZVvYjrEv8r3aDSAW+NGYwo5L3N8LgDIRhJ3P6MXSlqu0DdMHj7ONnld
rFuRgrPlMe2TIEFIhTR18kgNAtcrP2GEzuOAoOOzWfzR4O4sFEa1I/G/q6n6l8pi
4RFO+fMamIku/zziFRKQWJCKfPdJsWaSZazKUAlqlodV9SwpPdMAIE3HjFZ4HJiO
wylE57HtMwZjFG/31Wrxm/ClcYWBTLMsafw0ZmwoXXJxQ+MBazYKGcaVUKpQ9Wdc
oR7727keWtkZKbTDKSIh5mF4TO7XVlVScFYWl9EuzOgURiQA1GW4FAwdhmBjaZau
VoA6knvNQAZayDUXj0jg7iooGnGLWqcbzVoqUByJNrRdpc+gKAmKCIaYIMYgXumF
L1arFceWv8kN2ZTuAQI64cR4EP3brpbu+4KRur5o4lB4evqfbz7IdqLV1YXpcNEG
MwI3ljT9sTRVhOVWzYGJHXPx27TvxinUEC87BXK7lRQJ65GX4kgV3BuDuyOz+6hI
R13bRo0FSm0eWN4cOdfahDSKoTWnt+Ah62uDr3DDI2IqAUFNyRsaO1/i1UOesG+L
z/1H82fx4JjbuU2rqUX74xXBr319Pg05IEouVSER2ZtCyXjmOR0oZJv3fZSp6NTq
F51RbFuyxiLEy7xip8BIR9kcu4cAs7Pd3CO3nxgJnA5cCxeVucxmlYzDRVCrl7Nf
kdVAuGtxYfEnthn2zwrVR5zOy5FYHNlMj+w6WKAeGcOmJvkzqiD6I+/1Kxr3nRk8
xasml/Rz1AMBlm4WHjbrARSvfdKS1nOHT9LrB4GnkN3pGCFu/4ldMkVFp0bWVFvH
//0JhGJCr9onFbawCbzX6bm509GITw+9OgtjlGR6v/ebmfcDDAFIn2B3r9NYPlRt
z/RZpxImMI1S0DZp1XeAVtt16wpFx1MluyIYx4kbf2eRZ3eGUjKc9LdPJdO6V8dc
gsxJaBf9ifsK5vcCYhw/0KbMnJw+4BHQce8KipXkS6TdBDAxfuV+g/w765tKNnxu
2hGM0fj0QnhN8a2X5pOnQMMlwbn+poUT0+RUYpJLO8AEJj2ap8IlU0GIq/w2fypU
7ZNjAxXr4CVPa5RgZgziQ95dRXP5wQq3M3pQ/DyN72HgzgflLB1apNpMwOyPpxDd
WMD0rOxmODF7VFe/WAjF3LT7DQ5WJ85hN7YQcydBFj1tGUfZj1+KuVCWHPsZs1/0
Fh7aesLL75vvhJf+NTVKIY454aANR8HRcp1USGRf5uvNP5RJPhYW9zI/0G8tC97V
x+6N3tRHvy5+QkqJLa3TVsBxJ+f9xXvK1rvf0PmQ7q+VLn7OzmOdVtBfFPQ0ntPq
g8yTaZJvfXP/ndP3G0FV3JsY1CYQdcMAWG75Ct47iL8zs/yuaFSECkormH5WoCfm
0dnq7GUi/MnGjacCNe4u/SRc0l+jMBxpqSgjZqP6dgVruoL+vRSeRzAn3cfOe34G
rcd532GgRoewO+ZaexWoQtMZfOXWwSqyyC7RK+BW57fjDCjZySHeBwpawnj99U6y
NWNkGMIEHK+hzTTMq8v27khUn0JE/ms0G60X5s+X9ZWB4IonPcV8a0u8DS5IbBFf
943El+H4tJWOUh0KqxGYCz7zxhzJb69L2F17fJBjShseXwHXofh/ghL2U/6oX12e
AQfFykdvD5x8JtH6i0el9auaDXRFy93HDnpdzMtlyLcRiTAi7YxxW2Xuj+YINBEC
2MALpd+mr2OhTg4hBIizc4Ib8Eco9X84ECnUS1oa4tieFIejL/bTLdPsbwHpfjuO
+JhQhKKstE5CSvyMg+blnnIKWy2E72shBYkjwe7KCSEf6/1FPHe4xJGYfTv/JkPn
+PDgL7cPLwrFW82FkA+unX8QTiszCA9i89ZgtGR6reDfA3Bc1zG+cu5DOsSDeJr7
MvmQTaXuGwpr7INOxM+l0CIod19TkXWsN9NmHXoduKJSB/8kl6DxfwBGvYOQ5C7i
I3zFUSzuDYFUBasVSWAJv+Zyf7rgenLQf8cQBUkMPs8OlIQhkWjwubabX6R7XvNt
8JH/VecQe3beTfFBK8lFewGl/0ZpkZ3ycfXDf9XOoM7IS+9tpRwn+syJWy8z1SFr
b4+ct2FQ0fr0AVhaGQ3pixiSGyqg86qk+qlnzE/dmOnCLJlkAs2/pSxxTVwHSmDn
835YKbCF0aCFpwCtK0wKw7SVN4qs1QDQOM+3iFZ8uJXsoiW12gBe84z2x8A46JF2
O+3Foha8hO2sOXKI4jNWJpk16sOahvfgW4XEJxHKWXxWv2tJzzrz9NlI8//Y2puC
zm6JR8Ny+FDZoV2tdn6lfTcRRUwfa+7Js29R/2TOgGubo/p9zZiqtRc6pvZWj23K
0+oSxn6XMulyoykBilZ6VCBxbVfi//8HyfPSo5b1SJ3CUoQmpHOpy5pTE6DHdgaJ
0+U7z9Ku54Sv85aNEJ57ardojFXC9ipEGAFlkXkHK7SIH95a707noJADByMU8deY
gR2DYpyV7RE/Xn2dUOlZl2ov4IOvHiCO6iYVgXjBh2QkSXk18ENh/KgeIdsd4aTE
N569JwHHuQYuTvDymTXFtFjFqpPNoQYN49SMwDB8ubI1wfFHfjX9Dx6zw2nYfnIo
8sx3rU2ckycX78+nFoOEyuvh2qPJ+OSVQv6bz+X6EPm2L8hrXhzvizNChYHRAKSK
YBIB0Q567z8qyMR05wKvK5U8kAZygnd1CgicI+e8ppuuMzBPVRKSb3m0i0aCO2nY
ea/q6NRSfSs5F1WBFDpiZ0QZ/asUrsob15Eoj4uORv9bo81pksyW8dkumeE5TAVg
8BJX1XS6mKxKZ1zB9RKDvMMQcW26za57TC8EmAAOEjUQXTuzk30Siv9Hj2DC+8N+
khfL1hDiAmf5L1634QlyC/W7f8qtQHtYoD1GpRGI5GV+NmI43sMnjUrQ5T29z7nW
BeUrz5DsrhxSGiED6rsNDp45sScX4EGueLD8mMt9KIUXVTIDB/b+06gZDlOTkiLl
RPGpuWG9L3w0sTaNjl1nw6KdJmtimEYGlk8AW/qRxWt6a8TOlVOhq5OvhlLyyzlm
a6W+xDXKRsB5O/QOP4rZkBq4fIWygeXV82VKdipAW+z2FQLviC3w7cFeNSXxsJtl
ZrjmnNB3HH3Dev4RGrcNteiP9zRg+jpqoqBTQb8ee9G9K/UXU7Zzv+X7V1AYG+8Z
bSLCaE79HKQ+36ZHF7J7sdyAhG/rWbV2/SGmhnjImW3t5WUKMPu7gvNWfEp9xD5B
ZIWe18Ny/2uwedG9NsgbJf8q9q7DWNYfuXPrH54xWSE0b4sjC9FUFGVmQilCYQ95
HXYsBVeI2LYBvUN1Ev+G5WAQncQeD6bLuChmBd/IWggHz29dy0XmdUd1x/pTX+in
L+mj8tYRNRk+rDRxI/ww9lUcQyHEkTx3LNyObSoKg1zE+WuUQulKim2ndMyUdmMf
+6sXdn2cXe9wCkMPSP2AMKxVXagM/TwbyBvqX9W5qSGQBVpcI2Rbkhf5QnTYTIBh
MJvrLoAqAyGz+7ieqtmSHGGqsrDSBdZqlmldSU6aXktEar8X9o+bvZjO5OkY8Nnz
GcQ8v82TfMs0uHJk0ci30S1DagGXhkpNOt7PbM+x8TQDhVAwQ/8ajlMLsVtYMlBk
sZEofx5x72ZjfO6ultDQKTOS0gYVHO/TRxfwOTGZh+tnO4WdP0smgbuWCp5cXP1K
x515f8q9dSij9kx+9eK0S9UPDUxwurlz1qrynetDzA1v5Y9DpomDjl52Vm1KByMA
IINNdUZcFb8mbmkfJ9s9I9KzkhRzuW9nDEArWYit82WIwryDG4oqHkK9EAS1AA4P
ZcR9OZKslUwcVrFOdC6TOI4rOpk7f26VTgoFGEYCLn58t6sIwhaSnhYfNLrwYCpX
attqpjPGbozUjO5KF7ligUPtDeLXGb0mjCIM8eHi6L+zF3M2hnHCrJ3GMBV2Qrm4
hlZNNzIhtbx82468iSdR2bX+vlLo/7/3piIYfLHJ1M9K3zxruBXgCb07k0qPSIFI
MfGaz4VaPQmPvewTBu4WqNsrBIdvStHN3+xEOFRH60Rvg3SjtlTCUc0p8FmgkqYU
FJBTEUabWOOHVjBdbeMdqv9JngYxA0arwPcusYK5AYU8TaLHBVUTAqyUMAbVnDq+
p6klQlDeDe9Is2loADkUcgpe54rqny1ZOGJcytvnYfdqk2Wv40rz/VwXapxSI7bP
hwh0HscRvN4MdP64Z8x0Plmyao8hmDUbz2JECeUXd+bw380K8andmhTCr3RlWwpJ
3fcPsmGq+RPXJbXrjQAXIhvhgkNL1dP0aDBsLnaQh+znNGGHpOFB0c665F2vohS3
uIUYdgsF+uRqeXZAJ+9a5pq1+8xo6IH1TBT1ufuM2OAT3kmvVY1nCxQegcpxYDPi
JAxzUByQx65aucwk5ZZB8anHr3URuagE4111PwfogSuYbF0iMoe7eqY/MbS7vY06
sFReDa8nCQun9m+jY7MwkNMTmfWVcQCiOd6a1w9MX7FUeCC7ig+cCubBxAaG6fkh
3qODSSTAKWX8Rz+z5bPeK/NP7Suh2ZnOVNCHFkUaBhjGfsug3YtQgfeRJX+B6cqi
wRLo89Vhm3HlGqGdUAXlk6Kv3o1Gendmaj31dmtVBB3pr115ofL1bHXc95Lq+asp
NsPzENiALVh1ouRAWBnhmmo7+QUDkYoQkDSPmeVi9wn35VjsGrcIQ3QTbMecOhk3
hfqrF8dVnChRO6YN/4mfMr+V46qn0GC6VqlYBZ1XWvJF9aySfN/8C1KJbPyldD/m
mGOeTGLKRTw8PezwggJ4m2uRGxBXeCtUUabGqU58Ui6Ii1fbJqSQlUPeknJX9Wom
MoL6TIaw75GD6Dg1eBJf/jErvBYncirbRkzB/u99J+JeAS6UfohVB0C6+QBl0tbc
jnjYCs6fQacu0xPNqZW9dn4RlT3MpTW6hl3KMOjTZNDBbtNPgEThXf0okFlUMtMf
mWE74vj1Q0BzEH6DgyLnSRQ2iqI/Nwdn9hjateb4ADDij7V/oVbBFfXtTcF7m/TP
f1PeTOSBL0OZg+2CjPX2rwU/1U92T24JCTZrXvwldDYQ+LfLybamwkZQcaJSSqey
i0tZ5OoqBSRBJOpkcUkCg8B3Z9hQoBZkSEaDNo44XoPaNQqcUbbjhwrhqY4qcs5u
ZESgnH0eWqi8FBuNf8pbXD1Ryis95uo2XsJrcYlbTniDacWOBeZi3w66g5+RQvX3
osL7kACCGY4flA4Vur23ndRRZa6uv7XXOmBt9vQaN8W5Zane8YtoUevwhcIK0zOO
0wX4OCkzP6sAyw57mAgOGvKujAnN5kKBOFKLu19cbcwndJSw7/EiLRKSHGWH2Xqt
r8LLifGUpTPha8i0OQOAxBx8Lp9QxC0TTqGKexr05OiRBtnBnEtpgTqpeAcxDPCX
q408N2XPHg8KcN+ppwXbN4WBLaL/VJijJ7ivRizS1aUTe/vNvzmidzUIr5+iv+jH
bBp3p904XZnhFqZMQH3ScjFjeF6zILCqkCKUzbqq7+jL3dpOg1Zi/Nz9yGAt8AO9
q+UR22txRXrE9vDBoavDBu7+NKazX/kFW+/eVTNGyg210rczClwQt4piOJtDNjeY
lf6Bq+mY0Qw9IsxPRj7Ew7s8navx5WyealwiC7GboNxFhqB3wij7gxnP5az4864i
H3FNX116vgeNQQQMsGlmqNr8hOMmfpS4Fb9vR00nZ/vAmvlVrG+sgEqVLGrA0Th+
sU5Ag+c8bckwkHZjUJONoJUobHVAwdrPmE4VtWiS6hIj4nunu1QCWg7lX71+9eXg
5biMCqJOluGHWIIXdqtrGI/7Jz+mkrCwEq6FR5g65e6mMmR25WF2HJ0Qm5zvFfhO
ozvLI1v0QfTm+p7n62cP3r4/5PC1W+GhyURQQOelbQjOIAIuQIP0mUNiH8MPSfq0
BocmtT8Mxot5hFEFAdEGs2TpH3CbjbJQpIvuvVFznm5TI5pofXLNgn+aWLHTvhr0
Bx5aY6zumMTniRP26TVWdM6KN7l1SiOM26XBar//H+wYVEB1puedxPJ+gzNc3jEO
U+P5N6aLUM1pQa6l45WPqd4uioR7fuJWeKKz0Yy2cUU4lNefWau6aRnMLzPL3b4J
nb7aUuKzdvl9wYrIyp24tknqxzup2Wa8h1p2JXYWdrcrY8yoKVbt9gndquWx1oW5
otiPiAHcXnv6YOpWWd3KQLcI/SZWNFmB+fZ3zSQzbcpgdzocKK1nwEZQpMg9tHWJ
UX3Z/+52mORzBydGM7rqF/vD7qiewF9zaIQlsDZcOskF7lf5Zmnbh7H6zHPIhdWe
vZ5lAvdoq8q6WGGK6PQZh2VyJMBLEzJr4e214iyhmTvSrYFw/T8DHn646AK7JKD9
O5ZxnPTs6F4CWria0gm5VMkirtnTFnx99JiNl8FEWWsPaJEFH+6s1rVdcK1vEBPj
7exQpHBRFwG0pPLAeAqKAo7aSfVlQT6cv3Wn6IRmxyeVD1pGaQs/vbEk7WCESPKA
7KgfgwwKVaMTCqUA0z2XN71ZLuQpWqlhn7aeFABGIdcfmdtbetl1biMykXAFd7Fo
toNhUGh8GRqUuxaWk4bZx72T6YP75B+Mp6DhwPE0x19XLuPynXukFwDSP2ohcSrL
bGkp/GFSkXBotXWIhb2HVnFas9Ny8v3M4ET6F121UeFbNR29sZ7C1h0wFy0OqDOt
o1neEi8RsMUQ3XyZup+uxlh+MeUfHI325Sx5+rdTY+SpvEgtrOhpyVGrJANao2iB
UbsC577aQMp+YINqucl9u4KeeOZCLQ6YM80REkH+wjQt/qLS/gniLZOffLxHLjsW
xAIPZqlwiawotgPKpZmrlg1Q8nbCpZ8LuogmyjTDXJDjnmSXszoULLC/iGOqVu+N
T4NBplHnInhEPy+Bm9Czoiif9RANnjNhAS0YjMNREVoU1hEueqssRgL+4La8D9hf
Q2C+2cJsp4maO67fv8sCxxDinI3fGSixUM09QPs2tR8zYjI6MlqDmA7skzqxqAOV
Q5LrT2HmWnut69zA4mdFNCUdh7KLsvxgKWdMjrRutP45mtvR8fuRQa+3F/cWKkkg
sCghhOakik/DbDmnTWgbd0uvOMGHHHivPtNWU1PKvzzWmVgexzLrbITP2EN4YO0Q
pDMLzTvhHHWMg2JU3NJAiscQvHlPQc+hSSLhR/v/jLIQLnS6Uw5rCjjUrWRmAdK1
ZicZPwb8yP0jpqFC5wRl9cYoVO6yEq3FlXslBolI0Op2nP4u6V0wxzcYRBipaLIw
ds4f3rbBVsj+StdnVzCxiV0KgRnWd4V1dmAU8eFYYofS2LHmXrHWaoAYAKcdSWwl
WvxFloKHuyb8OLeLw49dYlDHCDhBzvcuUpDWEk6r1BHnl4bZh/ajZpj89u7IJVva
b2GXOf+JfLO7fZZ1CXoKT44afMK3B1G7DZAT4q8Uf6aOiAbcIEv+2bQICZIEXOrn
vUSYdnltHSUjGg4tJ00mKYWOxpNY6ZOCG3HRW4Mqn0E6vWg3he2AAqtqha9ZQCje
lgYZTcIs8G3MCOa37vwEGjAVcc4wE0Y9LBroHQGhhFRRnNPSNOAqozvliJ1DfJyG
X2V/eEBqmXCeAxheT0tavPEox47wG7j5j/ackX8NeG2HIWTYVw0FlOIBa4vB2RK+
vfPJ3NUsm4anRMbv0Fl08RUqZqaVL4JwMljl2MeFcvxTuGj8NK/Fla1421g5EqZz
VzV/rGXzo2QW77+mKizmircKWrRP2owPZd7DPG34jyW9NCKG1icjjILA/JP0cuiM
9I7rfeNfBGJBuV938MCkVD7T5618hF2IDF588XdgzJEmC8WrSNdg6wdUf9ZDfZgA
RIVIjoFd/+8jqz2Nndn1rB0OztHHKRGDJmaTav/RNIuFln6tiuJCPy8T6LffoWXA
p4Pz/VBmSepZR0eXql0TrXF+irxEAOFfu+hXbiiUVUAcf/M78voaGv48ed0ACpOu
8xPKCUye0ByqmWhEh4eS8QC+VdRNOaxbrKBvXbj5Flaiplu1l/oNjmPFOSnGvx8N
Q2iRKCt3sUJZxM2KyPqziO2SwwFokrDjxa77dDm88odSgjTrbfRNmIPOA6OwxUqG
nBomdiFwJ4c7/7wg705moYuG3ob4umyLWZ6bplLKVbQrLfHPDLPa8k2vDOjYbscR
M+vVlBiH5M8VHySUx1SR8bZ+9B0X9xJCimsutWg9vny7ZNmnas8SFF1SPt2h0HXM
GBtug4IQwx9Q847MEnn3SBCUiUoid9hNZAcxw3PoEowF1zHAfPTTM0OOWabD94hv
UZ7OsY9r0KGferxyUFHvDEIh3pq97Bn5J1XILFd3xhujLTOu1X/GXCbeZnoydf/d
qBFVDz9WWke2a5LMvjuk09NRcpXShQu/j6S5Bghb0Hw3BGsklPO1V1/qGAqEvWWV
8IukgNy3TYEwmYGwG3WFvpgY7WXHO3JA30LADd6UA6fNkXwnH9H19rgpf0BCebVx
623sDWsv+uzzIorfoMpiJOX/Bp5Y89Zu6oVIYUwQxEYQRzJli7LhS7WgzIVZCrMt
+avWEJL4TILUQbC2I0FWtSyWAQdAcvP1ybrC36NY6/Kr9Q7kzsEeYLqcXcKwT0fH
VXG3PBGcuhoHq0WTQb8TD9VtvV+dP98G9VRg7LQybi0Ny/HlsQPCZozaoDNa5z1z
1myFLqtXIxYtnNKOn6yWkO7L2U/LEv0Uyi+XNsesR8bUKC4ZBKOn8N4/3s55EW9L
4iCvpX0PdgDapP27Yd2UxHsTRyZ+nLU7kcJuGr9mLRWAJ/TFOE0xqi/pic3s/Xiz
QiZ8JdzD2JCx9695U2YQreqPdwwOFFHG+Xmc1kTbL6woPuQtS0mLCE/J6Bp6E5m1
m7sO6s+UhpnnDq/CxRTnecGHvSDysO2EQRzHEwJFgowuFAZVI3k6EedfB/qlqGGF
bIYmiaeqRw4x83Y6haRdT+2yC1XTRYgf4GYNnGNB4LkRnlnKVdbpPlXWNqOlHcAQ
iK7A+WhYBrYDrCpvWaOqMt5RCKRNOUI761FEB8M4QKrzIgNa6QVrDcjOfcuVCawF
yb+OfXBNl3imACqfBEunv6cPjqu2aBmO9wvq0YEuQyrA0FFokx0n7KuwrwZLdEkp
drLHLQZrBif6LSK6qszAiB50di21/jyOIPAOe0Ii2GbwWXFCYbKxdiJKWAVDCmXV
jDof/Ar+owfD/iGoYbRhR3gS9fOkZyEElQV+/IhjwlEPFwGtAC9H7wZOhGtz6srx
odjAo5JP126NO7J/QXfzQsh15e9r55nGAF/UFS8Jjnq5LMRMfbWMQh4ihhs0xO8R
lepnJTF48Udte6zpSwvqsCBk6dze2Np0QJkS0MBXR8R3JLj05eJK1aLNfT+k18rs
tJtfJ9YYS6R8m0PkU+dcB22/ivq8FlBtzjRwZojMaIUsV8uu4yL7yO7P9aKgRj+p
PlurrAsA8IlXVmkiM9GLJyLStfBGiNGNCaC3KjcAaofn2BmFGG1oK0Kgq6Kj7DVH
roy5kfwQtdpRzh30sl6T0+e8ibomnt6u9pLN2G7vLaGakaVC7qZHTbl8fW5ISMpv
7BUSTI71o4mnr904ZkSm7LUG5xo8YmNG9r+LnEhp/RqxXOnhtP1lPc94PJbfzK7G
BmqqmQ/0eV59xwiUuT62CDufy+JiL1pyEwyPvPeRLWNWve6YkjpSU39FN0ahexKq
luW38l3LDi+rolbHmcCg58XlfxT3Scgk+TAmkzLbs2skohgGD4GFtX4VeDrHVZNa
qokwThjo72jBH/KrG8s05uOkSBM/hBvYcdqOyDSsjHF/QJTjMUqGZlY/Z4uEWw9R
AqSKyA4uV1GZZF18flpgAqsiIArrzPCgdasFeENWRetklZcmgVXx4g96D7RRDb6l
SQcqGUS9coOI3WrXrjraxn/7QBxqB2zseMIOpMmogLfPgQBW91unuip3rnGW7Dif
CWrmbPV0gSHxoLCtLBONJE0m2iEPoNg/s1wR54zbrn9tA09pSncEW6Joowl7dUZF
6enOYnaRUpUEri+HXrFK2yywEjiRfVgivDuV1mbCCqJ3h6Pjeny4UAu2OP0X3b+s
HOaP4vPoLchp5FujNHPfKvxSYjXg8aVSKUTSgRUUFYMuOIQx6C6gUCQMmHJrDfib
QHLT0lqXCZwnDw4D+vTw2XoJg6rUSI4Ql3EkQQyPfgS5o2omQezfBDLjzW0lmf4M
D2FqMvLruWnXrxUD18TWtIgOBgWDrKzj8CBai8c6YEzhwUtUffw/iQfN77GywwYz
TtbK9gTc67wQEu4fG1qatRJCuIVcnaoT0RlTb6QckETlxIJHeGU0ZV6JScspqdDc
7LCia9+E5HBy78UrOAH3OZvwOg5s5LlHF/sJclU36gqY6VZGS5lthk6rc26oor1K
REApHQ8Ucze21SBWoJBUMUuRpGTLzaC2NIqtUxfMQmgOfHImscAcqNwbUiX/jp6a
7VQIQBIby1je4H9ZWfWnAtJb6zAc8H6f6gB6lAt1LzzGvuluUPoSKQjdFpv+PYo9
F03JWbaee0cCLQVeilNU9bt4CWWbs7/LdWmuMymVjMUnzVKY0bnqfFPBT6rYitnX
MSdBgDuNrwd6p4iwlFeSkTOBHL2Gfh1YtuJfWt/cFMtkSmU9X2RPtucve6Et+0Z8
2IoW7lUs5grtEy7F2I88mpACVSbeRmZkGwpRSBKvMUDs2CmPdLmBD8Lmd/2rShJ8
y81hop+vWE6LKimrsEhUXpHjC9/YsSnWtMqWQIjMsFdoD2WTkTmy+fUKwZIJWrIP
f34f77tLaWKmovAhZ7OXAxeQvlgocSvWpvNzqGlZ7fglVOAqqyzvvuT6I/QvwFJ5
lItsktJzctZx7c3nGIlSq/FluAsKagwNAAoLHCz25QR+LcchevJ80lAG/d7vA5jc
9VzuJlwnsEiLgKq8jQB2UYiTLBzJSk5RfHDEj7PC3qpY4Y1DRY/bvqutZ9N9IsTf
D1tN10fa05Q4HHAkKKncmwDsXGKfQ7B/nX+iVe4CfpS2OHo9pGAE8lyxqTCMBFwz
m9ZTkL99Tt+Ik89LdycRxtyqyz58nNTvzJ2SmhitPPEyG8vK5D71bjhUQjW3XtIm
DSqgm1aRqXzBbynt5H+ABMj6GR0JltrT+qz1uH0sRskQMUAax3MzO5qz7Nr79sHt
3Hp2yLmPhMtIwR5W7SYmYn5TQ9tV+Z0N84FSn+kiVmlMTjps7xMwexsrL+WJPKn9
LkiJTUc9rXMuThRMNSEq6xYS/7DBW1Mta8PqyhpXXyjgiID3vRpC2wY+EO+ZIema
gtVvXUpHj7FGysYOclAPzNA3OxotA5INq6rSISK23vw7z6y4DeY6eN9NJK5ugrW+
Jj46yUHvW8wk8C0y1076cl9bBGUDQFhAfrN92fmWSh9Kt1xwUzS4dGcrEcoGQUBW
mLWnvblc1HX9qdf6elXcuqYrIrYxRPn4HEE3Z+43OzkNcHE7P392vkQh+Y1Uu9hf
QAapfbQcl6mNh+fmf4x+DBcjaY4e28w+2XM8D7M1mlETsJHzlwFxmea40c3SwHNY
WQaztfU6hBNSKHVzCm8TKitNK05n0lf1rW2oVRct+48N4mRU+24c/evhnd/7/YbR
2BlMDZg003abnHghEKpf44NaRLS9LU2bzw1wPUyJF2JWJ0feghkXG//XIQTLSYau
wdHCisrTzSSOeTOpV5QYB+N/5oKuN/dcwEF3pbpTmjMkJ6rgWGTDpwwb2Ns2pqGj
MK+brHGicx7EIzeW3CSnOxbW0VxaQmCsYJ1CB/JV7av8rqzjMV+O8GTOmGh9a3/j
J+MRSRLcXCz5JRJU8+MbZdkZ6MwxX+FRUNwOQiyxVMs8R90aycLBOsAJq/0lv//D
UouMJ9WyCeERugRbdvCn2cmBCRV0rOktlze4397tGOYuiVACyJjMmiLPEJ2SMKbT
RBylKu7IPF3qROdit87HmTo5ued7AXSQEkU8gf/K2jWLhHOKq0bp1F4bhP9Hxh35
sFndqi7QuKn1OXVZ0GODdxBmx+s6DaB+0SASnkNpYiFusOWTbaGSTpRJpfMiJ+bt
xRohoPM36x6EdzM9llxv2VCgpHLrmhEYLKmHA8r9IbwJo88Lp4Dwigh/A7F0Jbt/
DzFQZaQcbPGWCTlNn6TPlDSBAFugDCf6kk7pvmtwgRUIPFgzDW1x17ALwNcP/jD5
KzByLEvkq0omPesx7tzCNeaF++b4Gr4ah22cFjCgGQBbh3xfB4tvDHo0tmg0PfQA
2wyO+6220ChjoaYVvFW/pOYCvpnHDQmthVJEI/KU3Uj+ez6uFVP8nxz6ja8ncGpl
As17fv9FRSZjle+909hxCYF5QbNrI9Q4FlDoJ5qi0zEdEvXhLOxgAoHJ2d6QIGsX
aAPBh8DnSqsDNwTje+2jTZHkgqxJfII8RzQ3WoeuX8vPTff0cVI15eVIm6e7fGm8
jIhhlUHTXw7oN+mxeAgFsxD+DhWBsWXmFAlQj/+hqimgZnMR/R/1dnrUCqohKX3g
9NKIHrftsKuUB6sg1HTxMjkOHWINCQX3BWbGPMNij37e6BOzxkyiMXp7yV8l2Osp
N/81KRwLgUjKVR5qZ2WLIWtyvQ72S2cv9Mv2kDVDYQkQ+vpeCJqKiYDQYUre0Y7X
shPng+nnxIwflgb4CdhmYkahS58KXJfeuX6FKl5Ao1YMSTI1fk1qNAQd5W72dq8Q
8MOc6rmH9D2422iSxYiqp8+0WIrq0IqHBYtZjUVMdnxF+cOoDQ+EyYd8ZY6KD9c8
YkHIAvByEwtFsEYuwAkj/bV5JAFHFub2Kh5gmRm3aTg7ODw08Ft5/IhvMKoR6qRW
7izDcK1PI7yw8NEHVHCX5LMTkqCLPqTdJx/FDBCBujvZ1ke35vYyrC5632qJ32xr
dU3AMK7F3lEaB78H6NnZotwLWFuOjifIsu3jKLqmr5aDR53idQf/lHvQgcSOX3+I
23LA857A6MDetqIoD9fOyKlOZeullmyy5gz+glNBtq8jmv1D6TXYPWDoqSScRQPE
LXcNW+YdpXAYApjAIRkarDrGiP41YUHQ4qMchA4ipFtnTKfsJ+iTJ/tYziOIKwpt
Rerb9/DgNCDwF4KTK7WEd8PAxVX8gDv56cG0CrUenjiMAHN4uzsPWPNeIz/bTEOg
4iuCwNXDRd0sYE62NzXm2tcGGdvoYb5rgjXbZbOihCJmdLvIwOIYVx+NP2UySu2Q
pccZks6RamzT+g0Z3vbjbHEHYMo/wG3UwVJ+2o4aijAP4xNV5Yi26WT83CaHdmyA
f+b2V9PqDTVkzi3+Kk82ibvo+yXvsjEzISZc9tl0mF4GhRYAntKUHljTC8u70Jrw
zpcEDTgsI9W9HbZ41BW+OhqX4domnCQT4XsqwlX42fa+ZIbIVi0QsVSsJUkKwMZQ
vjj7kHTBVY6cEPm2/6YSy4cufgWWDqve4rOdjAuMM/ZIwIjDRB0xSeCZRGGwTGEu
pR1eV4EwIYhZKDrxgAJzsfF86Az3yu/1EIk6f67JbzCeEuR1L9gcXyKCyYfckFtc
jSJYo3+QLBkAtk8sMuHYFXIs6f+KhRilGKmxUkHIIEcKcyqEgVi1poVInJMkNV3B
zn+w4TNe7uybFpHAXhRK2vXoSUKp+2vHxo5rWalSA6kqRohpXr9NAp8glGeAQk26
ScrTKI+Nnjiu0kWFndG7VZyX7v+CmI8pJ5NuwXjbYHU2D6UyDrBPIYTHWqLQz+XT
AV93+h2uE9cT0FxMLv6tMec4MxfXTA1EKc9QDQdcv26pS7INjItKZvHkN0+3GFko
1KAxzuDqCr6vispSutCNlVLfH/9rVz18zlBk/n490sp+KfIUuSZ5C/Ix6NWgAFqp
8b7Iu2aSlxBOdIrcpM6bnd6tFVxZgtdJ4aCdCCP2Tb2MxM+MB9YO0CjpYHpzDG/S
BWrm2ke2Olb6fgRhz1Be98GVsfU4nBndeWTuwyhAhdLDwro5QCqj+HGI0PEvVDE/
ipnc+Rg2kwf/FJEFKjtgtY8o8H3Z3MyMsUCcuFBZhr9q96+3JNfyH6InlFJ8rM/S
kzxAxuThNNP0NgUHh0XkiQLi0bZcZV6tgnLgMivhTOyDnOLJqUCghar8YiwKN7y1
4i8mIhxYIKxgprhp1JJgotbF0NMrqF9KhKp+mn/gQqA+K0Ni66J6TakX/JQCIDfS
uEz4zfkrZBPaCXYPfKDnraFSjegPFlrTTR6VcFrSUufWWDrDJRZ/s1qggXNqjDcr
gNtxTXD64t8BmN9YJCOY3aeSxvSNgzN+C31ziuD7sCHjlF4i8XDe7FApFZhh0448
ulzT+up+Hn1dpqnp+PrvG5l6CRcvvLfuELNqL09ifaJsDqlOEc2csfFhfz6bQaIY
g/J//cKkxbdQeDGImREHTLmMejABCSHU9Z9OJSTSOTQG9HyimolF8xoQsw+7OmzU
JD6WfBm6px5goBxBeoWyK/S0hufpoGbS9GltdPVIBKAjjKnho0KMplnzn4QYb4nt
ej/ieder3fkH98zmQqFiUGeQxiBeKKZgaIORvwF/1uiD6vWtn2Z4GEcRmbKO0BzL
DjUE7CIwLM0SFEGeiAvxCb566vlcgyqeyqD2PSxpbQtGAicXIrVgumTMduNgeYiL
XDy3XZXavhYpmofrt9J9McKiYpGa0xAFf6Ju4YSlGeXERNP+g9J0NOZReR0m+Z7K
GNAnAsXdtBSmhXdqYWlJf/jkaGmJBJ/EEpWwclwDyLlGgP0of8zQ1VQUSi+Q+EZI
MnaIYKXB9UV94hgDqng+cKtU+3Ak56WKQO41UclaxtibZmhNVWvLJ4cNV/YhTAcI
L2CdsRP2/0Evt4JUWaD4ecY5ae9BTYtyq6edPDSGXXYd8rGBKlqT1+x87+c2Sxge
zGSqyiFQ9EW4UnE7knNAczyhGzEVivxdgBTHCNpH2ymAhNerbRBwPFP/KaQcI4Am
+VRKStQf1H29lyg6CGa4ZBXl0SVx1W/nZ2JhNipdlhMcLWOM+lRwWSKOw7s6TfoN
oj0qi0PeqWCwGKU54HwX8QuKj1oz+2rwI5Z4kY2dCt5SPpmkcFzJ0mnT02XUfcEE
eqIlLyNLIzxUV2HTH+pjkEI4EloCI7KNuuPvc3XCiDD8vOpi7sjCdCshvWUGJG0J
EtpHMYpJt4LCOwqCRbnl5vm6x3GNwNJoY0gU8vl8ZGHnmWzfss1L5DsZWG+bDE+k
54mUe0LDVFQJHOyMyloHBnpps4Hdn0h4gTxFeekzb0McOGVCidHyg/oH+gpcz/6b
u3+w73A0xtCIGmrTEv5Jy/87J6jBJltGDZiWk42cdyRjnaQrz5cMXfwZZxEcv7Lg
5ZFOX8UPY0IouX62srPoyzkTGKdRBlBKwahkrMdh1CNvgABTuBZ4dpDMH/CVkizN
kI3Qn4++sfK4apPNGABwyAciSZT/n0qtZnZlUW0U2+1x+elkCI0YE1XnFO/4kFsb
TDx3pBIYPv3b4pqTRDrQm+r6KAT4a5wDpty51JHrNMoGjOV1395q2zCdzRuonTpt
1NYY0ntK8MTEenK/ZcYx5qj/z0Dhb8fQfz4vBO7zU0wGe17/GD7Xgm4p1/BzZQLT
tDzsTs0xLVxXGuETyUpmTpE6QBpzhmgfTpbxUWfhTYXvEU/6iYnPSbJ25BJtZnoy
VzAa6rZdPnL9LM8Pv5eo2Y1JiNEkxRgBXQAEEZD8LdzAVEhn+lOUxZ8wspIJm9BU
8YcNO/Y7UzAz006p0/jIy7ZWH6Z1jfEo2r+BVsu/cTlvpQu1E/QXKra5OoUc1LM1
zahV0EBBvs0XMinPP3XOz3yMCprKSvYtLGzL6oIP92QqNMfVd9e2L3Q54LhHJmpl
bNpVlHZ2Qjkqa2/VEytWBmIiParWpWhLteaw6S2oKinTwA35Bmz93u+tDOzC+tBp
fF6XpRURGcugpmuUa/o952Wk/9kKyxYnqFk0WOH4QtmqdMDi8VxYh1nf8kYxxyuC
T/N2NPez4tVzwUFiZDlnOQBjMXBcY59fHG0tJiDyQ3wEDM/gWQSEpwIeFZ6Ht9jD
uTjHNQBmbc7heRxaTlJqfxGa2r9cCQ3YUmpXtc52N4J8APMDiX3QY23crpweC82/
XAYZFSZ8+dhwIlXEdjhpYBf8fC8HfgyZBVCc9mMefvntrWE2ddy6Dc+34rDewa2u
QRyOPWBwiSb27w6yshwWbAiIHIDuXxnu2jSNUO1S05JwbpdVxb8HMSf/ySDRLF5e
m+J5Q/tm5M1c3PBOeJpAaUsMRLJdkw7TBqv4exA0ELez/VaDSj20G4zsZqBye9wT
K7IOauX11z63cAsw2gcY5WQ3GvvR0oUzIRpnozXrCu4pfQuwNfeHWyEa6FFFaKNy
syXQp6dvo/FuqFttG/XWLkX2ABQ6C+1mh57b9ckCnxqYAtu3gWLbjRY9yVtsVWv+
kryYYhz17Qx3gG6KHyCdH+x/xXGngSgh2B2vwmXg4Uqspag3tUkSA2NOh73LJNy1
pynAk2VdYERA5w2/R7G+FopLIEI+dqqBkZ0WH4UuNhM/nDlF22rLeO42kitxAOLr
y4mbJM7GxodlMVWwNTCcruQ5vFERRcRGXj9gxjqXIu4tlS+bz5+i8BV2a9habZsq
Gtg+PcoufQiFWwhC75CeG8SX5Y17wGLsQ5zagCmTqT082Nkb+fXZiq1icHP40MBT
KMVSE4YlmYzDFrZ/a5b0qqwgaIDyNqwD0D66jxOUtGhLADaQE1t+Y999vpUe/YU+
oaaEurb9sIj/TJP2sy5rvrF2JtScupD8gPqpK1b9xLnYpztLO0K4YwVCtUNBPPHR
RZX7FrPgq8z2144fY7whpmlOi0eIecbmKQ3NtCd6qtrP8gQKyH14vB6/88YbdcqP
Kmi67bWLBQpG87y+LrKMn57VTK/aw0ZWTiFFnnpF5pOJ9nQmZiqCETb8PuosZLj0
oUviij3sIbQfYTMaREkddcRqt/APIsr8I5oIKG1HflSnxrAUy4BNr6E6G0gwsamR
3YHTYIsj1JrKlkj7YOS+zJc8YGRg7CMBN9+hKeco3t6KxfVsvefZJPfemkhgAGJ2
YAqtv+Akv7A358UIvKh27ptRnxTrCK8Nknh5zSZydc6oxBoZ+PTuRhvqj8d1DqC8
ktZ2prbjjBnmpPSvSKjU2Fqj86wTW9nuMsY77JkTSsmrAO+FYHE/2xAOv/a9JgKo
Xb54OQSL2SvIvCxmdkwTD3sNRCg2ZSYPSCOuNGXDkZATmHiOls/dlWX7IuLbtXiq
Sc8FJaQM5M3mUybhcze7p8t0i+HLYxrx+tFBamugiJlSOcYsgwiAGBSkK+gSEo2x
MmfxDjVMDLt75kzP3Qi9X7jiywD/TF6NY8gG7f+mcpeuMvQUHiPNCaLajvFjrT6u
IcpIyXWlzln3FTrECYqhPlG2H8/biNLvqiTMFAXR5b+Z5Dhe8WSPD0ZIHeC5wVyb
jcNV8+TJOvHubYwhbwvZ2ZojmnUW35iIj/qUfZp2OWSfM42Bx+R0xPtSawq2l4H0
SiA4sXyjMPc/smr9sxCDoI50uLqRDDigQJo3bqiZIBUXSkIGDtXLmD/7YUvM2MkD
wV0NLSSv4HyDmv8GovGgCCVQVDc/ksRxAkx+xiiorNWrC1p1l1QRPFDFn1RPVswr
5NYoDPM0+C3NOLE13C8IjnZ2nNdrzw3iB1SeroslmEp/y1ot/WsfJzFg9vn5zHkQ
X8vJSI6JnAybd4CCF+ECFpNz1s91hZ2XLfVPyMq9OQrwfhb7cJpD6pv99msb9hdM
/npchL2dg3X/eUirxBzNa0iS64xQODXZoCn5JEh3KH0nHv6mJShKib0iZz4VF9/A
DhGfym+OGqsWzYAhgYyFcrl70QaIF4tnPRFk2jnWln1kYOV5y4xVqNw0a9Sv9yvH
8Vzkrux9ite90pvRoCuxMOAGFw0evPvxWEZoAQnPUL8nWA4phnCLR/tybN+dXLAF
DXbT3rX5dDLnaqS221XZffk8KgLXdck8KCr5TUImvEWh1aClJVApkoj3vSTO92ax
a6tUs60xiKkmZFVZgaJTh7Vrmlkkz2FQZ7VdbAALBnOR8uFnAboTJPUIvhh5FHR5
MokCzwmAnY8lMBpp6hTXduyjjpEZ60EFs3buEhJLcgGVuXLXhI4WKlvyz7AaTtS6
gCDssXfXxbrg6OKzVwisR3oyGbCqOT8oaNOU1z6hRYD41UhoGzwsyxAhdinAwoJi
FYx4Ei7V/KUMFnYXBKLBiPNeDvd+AZBFkLQhQcITH8EA7dv7Faru9l4IB9a176Y5
DLrHdqgGPsow8rj88tNNNKmG0KXMV88TKqL1GA/kY/Fy6J4eRHZ4QfWtnw9Rcpxy
ZKLTrKGzVhXSfJKpOCPpLA4sF/Uex9kmNl43z/1L5vlxfH7oVVh2Lkg0EoQGHXzc
hBj57rEf0JT22hQ6brF0lFmPXvHxcq6easKjVWMFWQStqzwnT7wO60P4aKkNr+eM
iyzInIr0aI6NvyO24FLpZnC5ovJA/cfxZcdfgebfJ95G9R0VxXuH1kGu/Pk1eRRq
ZLuGI3UDUfKNrfhdhElQ2goQtVMvHxnlcgmmDZQwqBn0FOa1Ww+0ZbQ2Vnd/Mkfj
oEZ8sE3gSUJ9HxR5enl8QDkOm7ID408PyuX6GrohgZP1W8FHpejeT3y7c8ccKglM
0ymzvheOQtETp3NAlCgYBgBDPmyKEYdEEzNsk+riDl1z6UOPr3gKlpKwieLEoRVf
FSnE4hRqu8p9pm1cOAspqRvJcCl1Qcpy/xt9/26K+TywddmMx/0n5tJKmmpeIMqA
IvL/5E68pyovAhEkJ3WpLNSRqzd4Lh9qUuoU21uri1TrXMGnO5rWua1bzihxWcOG
QWKbtQYMBJJ0As/eaLhcGRortWhSaKQp5jB3gbWeSbUngtUrdzlqVByBbB56VzZS
tYiXD+TUCf1E1MZNshQd1uIgiDygv4QksgmbrsHH3eMQluFePpNdmF8WJsConufk
iIyjB4ixUEIN8llD+EsC7Mog3M3pziE7ffZHBdq7eJDK/6Z/P1wwobF3EDECn7W1
+ltBFcUvb79Bfk7zd8M34AUewe286yMf615vRJ7/dBB2gaKCF2buxMIgOxAeekAi
Wed+6+h5H6jV+nSRFy3QW3Ylvy0dv6LmZZjgMWqGzkTpF/Img7bZcQynWzhxn8j8
b9mrGkSs/SsCcihmJvsM5z+7hG14gPysY6vHGfE5rNDG9ysCfji5R3Vy3g2q4h8r
/6hHdqL+QczG/v0M+pBLjeNp6nSi31nnR/SLiyYz9kPSXjLukEmqlFzA+CvUxSPG
q3oKDUG06EK7u2A4cEVi17i1LWD7Ggzu313qYGyGF9RcnbvqlN9sGIS0Ij8WYegl
xf8R+iVle3aySnoIOIzkjGwo3s1jcuMXLzkk8Pza7USvsCovcnqMkP+ZeNsDwp6x
mwbUMZBBBHUkcpDQQoJ5eF+mDR3Mpeg8Mywh08FtoKsUkpJKSzhIgJmkKoXktgxd
cLzTvYntMlUNwuPGauzVj9p2L7+XbG78AoSgMC9+n6j6Sx3XHohDwuE74UuNVvQf
CVi4l+AWZKf9h1FCKsAdwkG3eYbUbttYASXf/Xk+ohZg420dJReh8CMIAvOuw/Cl
KlMxtHn6XyvKanJBtzh00tz7OAveaSG4Rv7Mg6WelOZfwRdsEvJsb6yyNRSqdZY1
06BRhx5pyjk6Ybxdk8+/dWNQaGWnq8YaHybRZOOq4ghmn1I8RUcTuAVRool1h4Rx
i914Wld99JX7LDx7zQUIcpICIuslwQEKWyKuf5ZTrPLC0FYu+l0UzcLPVnRzOvm3
1KXXi0+VnywmTAoZK8rqt0phbPEOfCz0YE4utjBJH+TSEqjVR2ICMMFFAAKDY2tV
W3Dng49R7MW/HMFEhoEcmJdgCkhBsvxhrlfc2fxa1za0bCkICl1pXygJ0YLeM7hq
pkmxzkryrsdSAGhPI/P3HS6hbnwGQQCYsGu0XnH630N6eZYzFwN7VMtIzgAa0vtb
FQdUVAsrtAXZmyMGyLGK3EJDjDpLZvnhW0xyfM4KxSYCprMNJ0HKHFrDtamHbvLx
kU1V/VpxRRTVAWQhawgFKyUbbBp4m5qwsc64FN/eoeWG5VLQLj/Xn9jrpRyCREeE
477TofQM5Wt1gn38UiFiUfFT/ZwOdwsH9sZtyBQD5F0zGsYlguR0ya58899sE4ig
R4r4alXqGErC6iOYd6A/8y4RWPygsts3X27d2fFq7X6YhFS/xNPNed84kJT5Wkos
FHgFlb98BZt1gKF+kXnj//xc6Ld+V3AMJ0EghxYL5NcMBq8DiJxIvqDMNIlwfoQ0
Mq9GmnCxNNnIRnb6e58b09tm1Ahhtkx6EW8ktqnQMHp7h5PvTBx+3i2bKcOM7v5I
i1Hl356zu4CNKNAhtOtjNp0FRv8yxnIGIK497Gq8MMPsARp2vK2u8KfcCSOOeAFq
Q1Zfu9+56sG4dTzKQlRwyyVsxWU5f9GPwdTvZ1ZdrPaqFf/Q0lEFS86Bb2P5wKIq
6linkXBWJYgmq6mC9/pCscmq8AdFBfnzkJtC0cjAZ9WjOsejD7dxxN3z6sBp69w8
WIwGY8wPFuFmTA4v5TpT9HUeDMV6LkfgOu/p2jvPkj/WLCHY2KudCWbr0qDsrqat
qoyPKQaWCWAvB5rvnjNLxZvRQzA5HItjYQ3sV9k0xKR9uGkGtjSFj3hshQ4nW2Jy
AmFI6HNNOO8CeBC9ovKKD54KfZw2hfBTqSsh7HHKMi0CDHVZ4odu1WB2aptt3kHd
NlcjRj61jHzdJjd8sDyFZtmIlp1CKHeSSSgq+Lgg9NtWq/x+c1qEqJgwGILiy6Vt
b/xot/KvRbzNFVMlatZASpL8ePZY9d5eWnblr1V1uvE28bsiuVEOHT1de0qdCihp
Hvjr97ucLVqWTBpxLSmJ5m+0XpBWkGHAp3vG7CDCLDSk+OYTI9Z9177PiuXg/MY8
LFgGJ3yFusu5oUZI9jolPJDMGHfFc8Ce5J3GYCeFrBcazBVvo4YvBMf2RTe/T+uZ
AqL4kXuPw9WaGwDIc0B192dj8YBEc3dvp5QW1P2lbV5sBzfYxEpejWn3YsL+NjGd
haQhhDEqz6hnGi8R6+oneQ7KaNzZp+45RcVRxM3Jxh2nzoT8GABbfUAdepUNPjd/
0NxSLEYiS2HrZeP6/3flR14z3k9AnzcA1uCnQ9bre+VlOVSk5Cc61acVEvWtKGIi
/qGmW6gZ8L4S+kn+qG2X5EHjv2t2ghlehRDKoLWylbd0kFXBVbSg14DcdKEhYoFk
3VRxy2GTJSF5nTqTI7STw2DPZ+vK6U0uNsGS5T79hxQBKn/R7A6v5NeecY8FLdX9
27c21lIGaZTQDtOIFNIu2Saez+fw+Vn9igC5JGYxoNYEkZiBWEfxxH+NTzujqos5
T8d9KR2UQqUs5MQtEtxD+85FajRd7ZyOOUnOTPjRbtlFmf2emr7AJK6hmmQqaHrp
2KTa2XOt7AaEMoAus65xNKx4ckA5oQnKw96Mn6J4JNN0fnNUXXulEnEand5QGaVM
N+9I1t43YefeGaW7fwi4GTNsCQXMAUvcvIs3qqFfspEyUcV7TEKL3JokacRCxTcV
SWX/RyM7PUaQJxzS1q66Etj5zDJ0wOIxZLFOFcdNaM6DUbMRnDrKZt18I/pVj6lj
vP3kRYgZ1v9FfeVoeU0QeFPY3yDr83lc0jYmRRRXYLTADnv9ANSV0LfGFbo9Qzvd
SAQpDCg7irxvrKOJMVAuO45+h4b1NMeSCzR1Uu7i6NLjal11EXYaxd//z5+CZFVc
pznDqY3LlKe+PJr40nSHTVSe8ipNKU8cXlFbr0YMbbuFxDppylJegChBRlyqz6wL
2RL57na987OGKVfWVOca63TtwSOf9MkTV+IKkBPh8WOIEoQvSCHhd75NGXLlEeb1
ixdX1VtM5i/Gci2ZnDVtJkUaFbHNX8iOzV8NT1f3M67fBm1I/sjxpSjnRrUWBAPX
IHyTkDaMHQkCMJGKAJFp6qKDwLMy5x0BC8zVeSrrT9AgmqM6xBSdUXSpfjjg0fvv
JUqH/Wv7zFZ7sVjMmdTez+AQ0x4+djlU2D+kRaUFzTIpd0oWP2e8cE/gaPSGwwU4
RjFdlikZdpqdHFVgJO2K91BAuhULdrwJukV7vzEeJ/L+YGRpxOFf2kNf1rvGKYOY
bM+FM7MeDTHN8XSecxZlUsGQjfIBFPbuiI0W+6cxE/HSOA4PY5TKJphstq+eUQNn
4ZCGXVWW/g3BBOHNHh/nN+XKeEJMVMMgiXB46DC5MJOT1t0stJXGvmoYYGCQmbez
saoZRUmSrfM3n5PlU3jVEP6Ph6MVsx8+hjqFkJ3JrqDZf7Xbsoey7tULhganyLP6
RyOCDjFVVycCyLEwVHyi/46DD0x8+/6DoY/yT4D64OmHjhAHo17YYvFCgvhOkI/A
d6jBwYdPbXC0NDDzwNWQLNIaq4lNBX4kGW/Ex/NQvdac0n+pNKcsizGDemUypChK
Nmey7Dm6lksPpCXqg9qxPirCd+UgKqWI6A4Rv6S5uH2PzO/dIjcU584uV+g/IkDV
lKIvJyb2yr4dzbfAbfIZE19MC2ROdC6n7e6bOAOBxDgRIiJ927HpfakV5hvqw6tf
JqGjPkimnseQv+l33tD0Ey05dJ642SpvYN5R5SBkN15mEpvLzinBh7GOOvbXDeZK
o+tO3HAqSZkD/K6napl9lCQoK+KawlSznGPTZNDp2czHsiltM84zhdSO/CyyMJ02
WVHflS6o/Tf/MC1iX7+AfKBPwGctwpRIQTei/9mudpbiJIFdHbI5JraaPlHbbsyw
Pcvg5ot6qp9lnDwrstTk1wd9RBkbph+wqinIqQZdzzaSX6IxjPs6H7LKJEmHyHxD
ZsBh6RnY3py2zFSk4MvOYtUBTirq9dMBUlh1SBigMQesnJnn60n4iauBlxd0xOB6
q+Q9eKr1eowoxOoJ5JZQW+orkDjc/eyVqcNU20mMIXlHI415EH9fKozExXnECPVO
lpjMn3Hk8WnlL31HvXjczeV//+vwLFhB7kNxJOZajY/FR5zr/NbXl0Q0jmu6rXHY
z8H521/d/vV3mbSegixUU0PmYcy4LZR4LYipkyYS6q1llk3Izn/QVB/h4tYy+mGi
p89UyoJ/GNrG2DuZ0jz8e1le+0f+LX1X1zGEbL+os4/L3Brc2mJYwrFMOCFGCpx6
x6ZpvqRsWyZ65tPNAlvoQwAcp6l9Pq+NmrpC4Ikp4GnXfDIDSmTeCw+Sxd508jog
tYQYhWWU9OKCf3I5gWtAwaOe92wFnxuJsVldwIGkqDXBcv9KOFACnqXgoM9BsFIU
5ifP9l/LgqZa6y7F9ATSF9/rxJrHAMmDfOMzswgewG9XoPyfkW6WiyBCwiqwmMEB
VPJtQARjZiRC1uyARALTF0M8JduJ+qtUYwfy93Bxd7+Y0BWYEqiM7AYp4pWabuTg
tebwm195e2lekA8RQzGOqzQpkH+11eMPbJ5+lm93Driw9kUD2sj0Msrq1DWOfeEh
nzcW2HpiTBrdCbQM9+3FHeMkhkcUmsWD5syy+L0pOtukHSgexmWTktWOa4Gyu2Uq
oz6myNALGzxQegrjguvo+0O1i/wdNiYrtrQmoZAEQR2WcVZA1+2xP+8PlOHAjqQq
NBlAPncp9J7gx607vxXJB6mmISgsG4ilSF9zKkASSEr/NJwGzk45B2w+wOYJ19vv
F1DgINX9zEvJXEiG0CpgNMO5q2TXhUBHFw8V8/v8CuX39KwLS4rlzT2+Hh7BYltV
QQiDXECFt1c8riicNf1hXGHkRfLgAiNVWZEu3yrjy+5vncGe1VYC4VKuk0nyKVnk
hlohvRaCPkZnpiv6rwPVE4Yn60tFjJ06rmPgUbYbaM57xoPfGov2sfTTLHhS7CdN
3SWr0VwulI9LzN3lNVn6JZuw3ggcU3vbYYG8LVDeLxTx12Gkt139a0aDQWBhMFWP
4furJj7U3KT1qtK3DipYYEpWJ6Vbme+Pt9FtYZ8pZbztUJ0UwzsjvpDJiQv14Rdy
58h9OTrUDgu3CjLPPPMWkbCcQHJEfCJVxoNCtqRzuGva74R3M/Dc1MRut4/BoXuv
bFdNZq388D37NYSdIB1RxTtch7JMKmO7azHw6BTiJVxD6KFlEOP3nv6xP35Y7UrY
tc8RQ7m+1nkRNve+8hXhaLc8HrlSkMXkZO/H/guzKDRcho+UN0WbhFb4f0s2g4aQ
AgLJGLj2R6hLT3I/dLux4AekfiVNkZbBwi96CyA0gbV4bTNjklPotS4INeG4yLPZ
I0SRH8PwrYWkOxgIb74iNF2V3JtdxOMdImQWlwk5LZaBUex06TQjUTeRuZt6NO8J
KpBMeFwo+Tw/0ZN8X/lCzez1FhqKHvLVXaDVVceRVgfQSOxHV7ZLekgTcwPmH9pR
+YEPHEiLDTlseK/uQwfSzW6wKtZ/xL4CYyDI3XxPPVl+C0TyLh51cK4k1NPYk0CM
Bbdr6hWwFh6vKcNQe/XuQxFnLi5EFNmMa2vH2yqT6F1RhUDAk9A8KpSQFhVM6Ojz
Pl5uUsQFkUj77pYcOA6AQkBknwYt5SvBe/97EWw3XF2opvPi7WiTyPUvxJqz5zSn
HtWdPEtCMRvFIDquW9xdZqiZft40n0NKtHM5LNnPArab5vY5mQV8fmv7pFB2HMqF
NpylhrSI2Z5YbbHQb/7A5h4+6OTObZuK+lVNrY6sM2ZbD1QBorYHlvFo6VgAAOm5
By4BdH/txo6SuZEAVtr/ssRwsQnsH3cwINY2Kyl82BVxOznQyjBcI0Cq1rwuYrlt
GcBZawzPkjr+UHl9ixfWKFGB3ThEcI74+AHyZzeRw6IGjlFk71pmXlIc12Y5h4K+
BhgiinC9cpQDs+F2UcPymF7YwfHWeSIonCedDvw/63VQs0F5PbFzKb6OE8n7psaw
6/q7fbY7gNfv/qCFBj1sxVcwuRLRU7WRwp8+vUmn/9BibrmV2tHVhU6SeKoVP32T
XB9rkRDRzCnBiEG3Y8pnNHYuwxTNX97fJAUDJgUVEf9cKNHxLg1SlwU4FzAoKwUH
HaKWqCxzV3KW7z4u1QpV1BM6tDmv4Mmy/Lv6qXjgEXkUtFHfKS6k2Ilo9Hn7EC62
1dyYyJ4zKkty9mCeUN+2Ia/U8x5OWKpLmwtO81U+Bem4lalUDRVa12iJMKYyCAoK
ojgmY0p6/jYV43J7ZMVQkKOjBu0j+vv801wErRx/AvYTvLeXXiBA1+T13xiDhENF
79QuqZoUeTE4rlmrFjo/GpnxpM/pMXI2/CEW/+1orf9H0gNLSTPQTt1zBCPb3+zf
gjQccScvorB8BDfc7hsY2VZ6Q7eru0Xo9zNj24+pyyzcWNsOSmRZ7aGsz6qVD1/s
Vz/uVDgODBrYuKJw2oFgiwedJ+JKYIkbEI+tu0JtC9iAW2kvZfw4lo3KU3404aCO
Wa63r6HLwX4T65v9Xo0o5jySx1ngRc8d1G0NvELaEZyIGo54vIl3gCpoZrRF8JwD
BhDTI7Iv5qxRG6CpWDtklql2BUJozE7YbjZm4qekLRazJg1NNm0Ac+tJjSCpaRea
zsZ6PZc3Fh8AaZnhd8SfjU8aVHKTaKMRJd6YtczDYY5MjcFJjrYj/PsxRtDfXTqH
wBCcuzt5GxNYAVnPVh0tbpdsOcvlqRKb6I2AQpmvMN7oKbb3csDUQLbkGuDotSpP
GAzdAX06EW7/kobt/LV8jKxsBi1gNZ1DOPOxDuYzFQjjfwflm1tdSClWeFdjsLNr
ZlAf6R+5ZZn171bUZxfmNqBOOSeQqNgFS90I7uazU7dgWW3BnXlICV4dsY9H4kaf
edk2CAkwaj4yUaic6h7pi16PNiLFSmxHyqnoUiNqA6LbMc9WmCOL527IUXdIznn0
z0oNDqR87vavxpPfUiF+ynldFUCu8OYVhRqMgPOsUh/2iKCKQvRAnVldY7F/F7Xu
gawhS4sV+koimwi1jtmgtHOUMFm3ccG8R9DQBmbJwFY4avzgnebQ/7ueSsL2N/Ne
0peUuTkxqVBiyK+QRSJXPKxthJ6VtGOl276quvN03RtYoJV7vqinqNwS5SUcsFmx
Eko9b51UT4L9pndVwfIaxhcGUz1vXTTxklMA8gP22GU6IkO6p1qZA4bMQFloTAM4
w3HxQgNKsWL7hvN7kh/QO6I121JsZVZv9SNNCrrI3854MdgNzZWOCZkE2DfNPrDN
I8TYJv6eBTy9n7mKUoClBNCeRsp0ixWSU3AySR18DtNvd4Pa0jXMJjBdHbfvOZZG
nCKaStDiw9PZ0i/HoW565DqwLpThNH4OihSCGZgsFnTBvwshyBS3SaWVrYrjsYN9
PthIgtTO1giDfZuD6z2q7WgfLJv/8G1MdC1W0B8HcKwYFpJvE1kFEer5DbNt7OUn
wbgmNEZ6QYxWhxanfh5ayklk65aoYfK8ZMHxgwAKQAYVQdGe7gF2ccQYGsUy4B0X
1BQBLJhV9TEVFvJjFfwLpzqVCkmxO3sIh+J++Qd1ngZ9ipRNPDV4zHDGFngZeKkk
bA2T7jeyYDn4F1JJb+qiXpWcB+vWSni8qgEm6ILRW+WgwunsR2jIJinAVrJllKhq
zUXl6BSrPTGbln7WAur5wu4Vto2wtB4jtglK+HIKXtVOtAe9w77MyEgB4LMaG7Uk
+CNU7u1bEFj10VA7QsrRNvdFyUn3rMnJ7IrX1KFEZlOqW5sxZ9wuM3hll2u9KHnv
ehfGfQk+YZY7oQcMRBIOGP7vCoFGMOxxHLsP5yLu/sYYkT0vkuBJ5H7fWAaXcdrM
pv32HkJvJgKmxMQfpKg4fzQPFoEU8SQSxOVPVaQZhvQsz6wi5B2pPCbztv6OjPkE
V8F+PKGVVKFcTmZRdNM/BIRGS1GFxe9y9TROXGO0wKDY9EqWiDj+dyHoWL3QEATJ
shsLlaKCR1HHSFnXihLws/Wlgb+crPtjhUG+CtLKABolkPv2/CyyvSIvIPzpfaxY
WCSsabmf5J22ojBtaHAQw/oqlJq4J8uo1u1Mfn6fdcS2Ygib28NHB/9GvMcPsKFg
mTrQtL9YjU1FVgDaNoZalbs5Es+ddF5HOfuU/zPh9MpoPx614qpAWPuaVq/YyPtg
ACIuT8TTUC7gvXgfjUhhbv6sTGA01Od755YJUP9b8ktSc54i1ARVpHo2tAk592PB
/TPfgu6+uIHfRQ4aExUHPuu9NuFzHl4fuvDK9XsUTnkIjY82dhhp5NK54fW5Dlg8
NqAwEweTKHfWd+ocwviUEw==
`protect end_protected