`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
dYVY1GBMsK1ODCn3ZUp8SoAWP8Fvt20jOclKciHf7Ysn2OlvHpNHbXI7BFbSBeZ8
c0HSNxtSIQSCmTTcVbiOe5bNYdnShY74EmVDlUagwaODhK9Urx30VHPfg7K0Q8Dj
u4EuL8LzGtWyNpPuuYUPfH/EWWJz8j2B3GlAugKl7fR1RciktYEXyNArDzj2i2Lo
icoQhkynNgC7v9DkMLR1BxAwtrFrckccZalCrbzlnjwD/DOLPtfjLaczesJPkKoa
xZJUnnMJHmZHdGCWDxS1eicDF7kXXzsE1BA2jAX7HQtg/mw+vmEQXKqvkKy9tRtW
yhUEHOXSIVFkC6gJ+buK9Q==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="SgR4h9hEc61j3UcDg7JP89NUc7gPf41F4aolx7zbZ/Y="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
PcTZf+e633x3tw5Pd+98Hvg8K8pEx1TP/UFyHup9OvIvZyp7VdJ/eQ7Czw0TCb/d
NGL0fQmqipTyP1VBR/CwCDPv8pUq9mWdoIhPzGBVMq1ZfAiLygNMWUwFu0/xPfyw
rAKvJfKF1tLDCsja4oREz1+w00FDmJ2gsQcbY/9d4Lw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="fB5pBzxyhRsqq3gFtq6qZ5Drx26WwP+GzJuJsgJq2oo="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 37808 )
`protect data_block
Pw0LuTSwA3gmWF21w7rVYBcj97hqvAcf4dxm1w8M8xOO9V5Zp53fD6281Uk66by2
V+2le3pjRQ4JkfVvu0vvltrqFdWvBln4SM9xPIyOvOgxR9dZ/mACNvSM4sNQA0B/
jQTg7+iVGf71qmS2kysHxasIsPzVEG2qU32O3CQ94XUprc1zkAQo2eWcwRz1MVHt
xeBxNT9+avTKbyRKMNvW2VWDPuZPnEvw0AOsUVsGFbzNAy72Ig9Ix0sF9opOiCYi
aTSBDVRCoIZmSmm6Q+zDE7Kgqu6bt8+ZrJqaZ4HpRQJvr2VC5emCYyAa4e3gXgbb
1yzmB5t8RCzvN8gAI52Te0BDO4IdqcOx5JlzRfF3G1p3PCNURVXKyNZ5VGsbxqTt
3ciQ4O2JYkCkqvNeT+LqJXwlEBhdI0nDMhdS0gMNZUAn8VP5wdxdz4ya8zaFMzWD
YARnjnT527tXgrg01G6sDP9YLP00Eyk5dd6OwyOmD5Oi3yw1EC6vJbddgbnV0/nh
4lqsFM3GUt5sizP4L556Kis5cZzaLdyr3PV634LTvzukCU6qKoF1wneEbn4Gzh7M
HefcfW3roeozForNQOYChOc4rvGx0hnf3axnUP0ro5yKNZBNspO3AGQr7i401nin
WMCHZF4E3x5bgEtLLITYm3KVZp3/g4N1AL396JHRY8liVKmmvokxHqlJgllrE2YR
FLBGt0nMzd5TusBglaZ0JynVHk2axv2ZSiQoC94486ID4unks4V5OYu9VgNSFu2v
5Put95H+eybAPqgQ7R0UmjQ5I5ViIYKjRRr7YJHRroQyvjP8a35G0ZeWiabEm4up
52Iw92qCzbRbPTUpVlcKUwLJEd7VUZtivjk2qzQmc4hhriirHcI7anW3zzYOIuq3
TAu/P05D7znj4TB5yo6zfvpf8++89iWnXCb8H+JmuZaQLTqWRMazqj9oCFqnUhAj
JedYKqn7zMHjJKRgOa31jJVIzs8a5TRXLCXfmvJq3XwHSFNBVNHsVbITm/ATcK65
0mCspBdG217R6VY2Y1Yn6quhesrfjIJN++Pru5pdrIHj+ponmSsZxxTiXAJVnlss
jaxcderpcjK6AM1AnsoJVx6B/gK6FC5IVwvarXO76zg7wX2AaQOIl8E3cl/uNCvh
hOjZxy5+zjpT+3qvHoTWyX3n0i5jjChUdLRX6wsiW7QjlcVgG9lKh/dA44iBBolN
FpApykrK2luLSF4OHiHgY+3mTxYuw345fTFli87rdvOiws5EQ7KzyV3mouYSGlP6
AC7vkWQoTguV3PRPy745+EYEOawUTWyGFWImqjj2C2+QIVEKqVkydN0luzt+tPhi
hMAfaAcB5snp6nhPUyBJS5sDdKT+TiFSp3bU+xSz3qDAKhC+FxCg5vfRc/Y6QGJS
4hP9ikHXPfqLvfBzh5nuRMHbXUzFr5mIVTLmm0nD5BrBmxcOp+u5LxT8blmWRlgW
bhS9oKoVW3s3AwF2WsQYfD+khJ1sDalOgF4MBygxJeykbI99coJMLMntQ90eA7NU
kcD72yegAHVusjDBT6UZDA2HiX3JbHH2E/hplgICFbAqiNHxIJoUborJmff80TDR
KAzpH7wUjK36nK6BY/v/C8eubwLUcG/89Sq0aSFz3PdZCjYrobeDZabz0qJLkOaz
DqE67yAkcjMX/xuVaxqULDLoWse2c3DR1D/5bxeb9pZL8OSdx3mM49X/pN23xALW
PVpK80tgVpxJ7SfV2WQ2v/RLRe7xqAekde2MwEh+cnqtJobIUN+l64IHMhylsy+t
1yVy1h8tqNR1Hh+6x6bK7eIBve8x8yNrVcltHqZXXi9sdB+HtrlYEAMJ4m9meT+i
tTldha36XvTnZD97OzILWdUDV2T316/s3AKV7PpIHtbtK/Xt8YSz1Xte6tsMc1+3
55PJ0rWmyOlnUUXERVaYAlEOcViaZ2rsPMLs9/DgKFgsuEzLO2nOXCRequw489eI
XNW20X/0fave2t2jRt9qQzerIc/rLwq1omNIa754JchYOZzjyXPbmcNbu6FM0LQT
ioz+t4rQWFHYvQjn3mUYuNOzeLZhJjhApK9beehHSdLlPfysXJ5qjNVsvGQjP8KS
nbRhDM5u9Hq+LXAevHh0Pkb5GkLFOtDtMs0aUvsA8s5Mt0NyDtZYkDn4SB3ENTfh
bnJx0nZU9XBXA5lIkaFDQ/gzF219hOfAUDRKcraxg31Lwk7yb1Nm/jHOC0MErwLR
2lkr2KxSKwcRn9YMmkQfENa17A/uXRIUYip19M7HXT2vh58yppTTnkdQLbhrAP/t
UIrPStBFQ3PdAeqm7UJOVTL9Yg8bh6TQsNS7JHooYkr81g+vTk5cVkLFQ4jUtpYG
a7kHqqoGBIWp1B8XTgBESrpz/edoAKt59Vw1AQf093F/CrH+SNZF65nLY4m6Kq9c
5n+3DfgMVqEGLXcQnWRp7jq0/ixWqFUwx/J+2RBmS4PcyMQEKo5WDY2AAMmzEy1u
VkD6gdDmPYsvFff8vaDSIcQC2RJIYw2KIewzpUTvGSXrydXqEfU2BSlaSElBCN4d
aK+JTtfwaUyeL447myxm+eVE/2Uzz/ki9QaxrCEOOxASW4laDhTNn2/leaRlqwCl
BOYOXsavegJwUgQREgnPxadjmF+uFb6hEDU0M0u6uHLTz2PXdXiWOTY/WB0q5NGd
gA/te4iDs5XygRAszttVIffndxWGpWseTKxYMWo6r9AGTFubJNdwgyNLQtfn5Wpz
kNuqswEXjQCqmLrY+Ry+l8YTwRCJ+7zpYSYiZ0l2VKAOx3iFF2aAMKKo33wAjiTT
Rlj9B87NfjFAIviddt2rCPfge7InBkotfviFgm3r18pKrg+wWWVd+ZbImqos71HV
HfkXmfKLwUUrlPoS4N3iL6uziWcnev3Q5xQ69RS7jf/owTzgFMJBPWXlGTPjgT+M
J6aH1KXFYcuIFa0IiUfxLwuGuRWURVtyY0ZAYDD3JXZU6r3+98h21r6KZ15hq0Op
a28jPPqOCXId8LqDdY1I/o5HYXu9MnendsGhaaJti8DtjLOyT5LoyEz5rvxfJeO8
eni0f/228NXbnbPQhdemDQ5XPc7L3qygfG7T+S0mDErhPyQHp2JiJm+ML0gqFjlp
Ne+N8b7WHyocZVYylqZOV/yu2SkFbqEIoyjwBK3TbnKSMJRz2eu7cUVPmO1/QM6Q
yYpQjhep8sWbLQBI6RYlmuxrrLedppcJv/Ss9rdzxxDAeKKcrmcvw6DujkZeudqG
fMJ5qyUK2shcjE2GH6T+0ss0w/M89CtIwTses9aLY4tFl/F/BnqnfHje4eXsllaw
OK5DcOhXCfEe9X5LrYQQJDXKgk38MhnI/+wkx4JDcd10nlAbScpYPHREhHfKdhsf
MtEJ5bpC49MNY1+yWCO7LFHE3NauS461CtT0C0DKoQ/IHGjzKVXQy5fpMUhpJj+H
Lfi7Qav4KBxfwvhTfKgwf543cFostBYE/h4TngiigvcCD80mL32M1pxNrdCiAGJn
369qc+xtUtzVKpLWFhEBVoiKCEC6E4qKoBuKzCq8FgwMavrAIZbhYqSfSrCSyo/w
d+dRsygo++MG5Dnyxfy0ILL1bRTtCddXMq6b8xPA6SywWZ6YghmGkL7cTQFzKXi/
EY/m1wiMq2VJYnLG+NpXZPCtMIvcQUxJsS4tts/zlCdyx0WjScU5NPHvFwqkUS2m
cPuLmpSj3N/Wy9f6xnoCLbXizzuTvJPU6vijoTA/PPDcojHJAUmso1OnDwGHX9Ea
73KVMfKxm+1NOmTI0yu7h+0ShV+dAEwEmE6mBOTG8HGXOg7/FZP6Ltf4ruGAAQEB
upeFYsm5ex0G1hNgOL8hDUB6AwE22IgOf5FqdSD3d7LkhsWtpaFiOqx2b7E4NFvV
JDH2W2h8VjMcb19vXKYKy7guwWE/A/1I/jirXGf2gPQ4xEby0Y68JQSC4lP1cobw
swiqYDEU/5pDDl8aqEIomd9N4BnLzZJqGu7ghhNJljq9K9ZwTAg/wdfVq3yPZLmf
t+Up03tmHlgf8YRId3/bUPh2KqOWdU/Qg1R8cCCq5pBlK1NYs+5ajko/gdWFzMeN
qrQPJ8rlu8KBqEdOteIzfP+CZV9WJv2mJXpTnfIMU0LQHUKmNH8lC7RCuzvWi5QU
52FLGAMJwaOGanNwqS/bYML8WAhSiRskb5d24K/vTQIzH5EWYupx0PxUWi6udcBR
2pplzqFfTTaIHr/CdCIKmNa/NB+ksWiKKPPGCWyzCxL/x4Zd9IwU0XA7M71hekhN
7zGDDPmhQPfAXiDHeUYVGBvYZPZSxBuY3e9lHYtxPcjXW8eVS0vajw+BOlrUbt+t
uY5czTQqOHveTLiLTB3DTgqzUf4pfhE6vDn0kn4ZwABxPP7ASbCGYMTGDAxQFSXD
K5AFYhAvyrS0TTPs9Ql9F5rGx5zklBD1j25PJdIk88udikFnClRaKIWBiwdT7Ps5
5FGbOBwoH3VACn2bco6e7+QfjUUCA45sNxyBeqe9KMkD3JiepGUOivs6QV8VqkFy
0+DQmwAnWZLd1vo8HcRbflV4qKxtuDiw5jGIGTArV2kBFYSjL5ztPmLlnQLUs/zI
ysK1hzZ3McV/XsB4Gd2wGDKa7Ypb1iGpBE1/lJj4xUywd8+25P40ReLGul4xBcQs
Jk8kNIz4XK0oKppgO749dxVfv1qRHqXMRY5bBk78OAaDh2WzrzzuPAm/+/T0nLor
XTGrG+C4HR1U51Ltopv4w36f/sfHipkvBEQ6F+zAukUIOgnCsscdN+2974Zmmf97
QB3bIfoLw+jWt7SB2XMlgLm/WkuRgDl2xv8frP5mRnKTOHzWsu70TH7Lw7aKxmRB
KygjMYkSbsTuaqaxJ/8Y/inSXjX4EtSBid0ImwcPPiSWpUitDRTsxgnFpDodjDwF
L+udq68eWxJwZIoOiVu720wScZ8uv0BBLNurfqu7fnSkr4OheSuEztEJt7ouLpUR
YAM+s2XVmLvfwuVPMNtNQBtAdJfhOcUa23kIyJGIoVta75Q82Al8oOyE8N3uayjA
VAmjQrznXr/hPY7nBOk/E60gN6/smXH8AdXXqG7THmRuMJl+TceT43LbJgM647Z2
L7VLfvmxyTO8rYSgdk4tolimUPC9t8zp5DoqksDGqkuI+CDxutgt6p3iex5JaFf7
zh55FCZqREhdb+4DDtAak0mQ7R9kEnL9wH0Oh2Cg52YOS+eIYBGZFMf5kh2m8X3b
+dB6XpMBknLlZhwl/SQiVm6dWITo7mOlI6WO//6+rkPlRsZhChL1gp2DMcQcK7Yq
gndOCh6lJXWkpoj9gwtLxhqHYgTq6rwpOVu0IbqyzIy3VdpxrT0f8swl7QnFAOxl
HDgSTi9A+0v94vtPwlB0c9DP+PrMG+WqV0xO8H3s9+Jv+VXFRhabZ36Nren3YriS
1ZmPE/+W9JI++CVrqAYAWv3hSGAgY7UcCHiDhapUYXQpjz1Zyh36ypEA2OLhgIiN
x+GjbNFb4FO6NkGg5TfHi6VKdj+zZ5TlWJO2HFTwJp5oXA8NYwaIvPu8ElnghrCt
FmJVhyXK0ROOqmucwjlFgbblloca6Dstl/auEEnm0jn8SpeZJ+sOIIWTsTWTypmO
jmtIcSF7nn1ftBeE/HIT6ZxSz6MaoN+sSEfzNsA8pzK2LTa/rRohjUNiVEVodifL
DWOdf7bOXQ/6Hl17GsetXBl5dDJ0qljm4N1yXdw/oBnjOZ1YsHPkCtXOGjLBZBd9
SrPWQ2//b4B3MZxyaIP8COxowFif7Afp0bXQZm5F7N1Yahe7g0LQRVEg0W7eImxn
FHFb2VFSHBOdgTeipNkyfLnKZ28HE87ivbglEi9lYVhVKds8kXp1mkxFz+ufmKPe
Q8yssOVt4r4uyFnGEo69Ji3cyHtFe1v8nGNSIfNVcUtuH//0cd7il/w/0HUlUXtD
/8595CEPpLvEbqgb7KG86PJYMGpC5xczv511e4Y0dAIEbpuBOSWP67LY88e6UUr8
/6cuqOU+mpUStfvj92/D77wn5CUKzdOOFepJ9vzmRu668VLjlek/7pZ1x4dJqGKj
0I12Zl+8UB6UB/V6//D0VxOKowniuWgaVBE3mcnl7Fn5mtxICn9FlxbjAHT+nCHz
R2UkDfmrd9csT725YyToYZvp4GLodaXgnMh5hq0b6Gp7T0aSP4835eieD6w1EKH1
yItqASzZYS9wFdDoUg1bwJaEk9SA+5ZMrfJiQgVRBelEW6fEau4g+RK6s+DRskDl
Kl53k+KTkkxwGIp8OZL4H7+8wpAvffMw9VmbTCZC0dmme/A7TnVQV+aBaO7tWxm2
KBC8mElrT7AIWiFymMY79e/kDr92QbYwTqe1L7CbX5+fHi07pNy2kPNQI+wqzZqx
+DnNZVinJwWyIR9tyLacN1Ap9xw79T9NFVE6ThKRNWiVT6iLtX7japXdpqUv6+aA
DyNz9QXLEi4k/TpNkzQCQJoj90Mkd8CHXPQx1Z5zq2ivPWDfyZ09Zho3CHudizwK
y8IL9/iGXu4DU9GdlI+T36eZ6XpqDTns/hca1VqVlffGpM10ig4F55PDoTP/wVub
vYAtCUjFwnXEpt+VbrYF/k2n7jE56scFYKucsaY+BW+8+FFUVcjjmzvbFcWHIBsy
AcjrEIV+LOzRhsuzqw0shHVXUJwEqRYeRzwGv63xRwoiIlEWdr7MB3vzyGEbyCAX
+wghV3oC5N3NYr/HG84/Wl9DdfIRkXHz7a/WWPCLHL2osvEpUlBcuaqepSCDp8YF
yy/7PWVWJjLXL/2qFPqVKPhEkOq8G87hKFFs1qSRIgPNKheJwF2fsIJatdbfJIr7
dA1wReDXWnK4gZIsihJYFaA1/hA+AXPio7YmZuVpLPaIBdX4hXuXAXaQmqUJKj17
KOU30yhQGX651bVZsLVtmn0NaAXyO5pooVFthMVtsS3WqwjqNNS6A+WBJ3w9zVbl
DoQtkuUY84S0/CR9VM5Iu0V/ppoh2CcOadnKYfqys9tLn0XkozvSUyXctFxQekBH
I6+V7wlad8zMyK0gouhhOpxw8MLIGxm0uQWCUS1Oh3tjqQuXpwfacNOH25krtjY5
f1mpAFLdgijoMjOHQ8pNZFSOIHMv1e5zsOuUWZJJyzLjF9rkQ8d5oDhrIjngjdwT
s/1TfujQOJcIqvR0EBTIXVgveRkt2gkney6orJ7d46oyoi7HmlLUgyGQLGgut+6P
MA+q17HO2V/hACxNmg7oaL9KgSWk7SG3Z/349ZPvhA6BfzWFUD+3zl/bpoGRQpiE
LTAa1E26+GqHvy3K1I7wPnzyqN4S+cCzzf+axrXbmNBfPd76B54O4b+FvOa2uSgK
/z624mQzlp5pwJInIddoCGVD4S5zfYC21JErajJWoLAAbGDfm4KrcamSJLiwDe5W
/9geNtx4gwHNnFxpJlTedo/vOUWlmZ5spruMoHwEbSgJSQo1enRlu57of//XzAXE
TDYzrS4n3LkC5PM09xIcGTE3+kVQ+nd895mujQEkTFcVVroLh9gTOEZzB2munLFf
XcTZ68GaIWAm7u1VpsBepwVGpwkht3hAJWI0KI92mmqyboUJujs33PdDdiEy/6rP
qwVuwXBum7h+F3NS/ZGGBRTOYikrpAp41UjNFHmMO1xyGie3tDf/Oovhh7XIHENl
8n+zW+Tbd5DcWnU+cBMl+1kdJcIBgIhuDWqB4FBmGtcR/iMiOopQg6oFE0oisrOl
11l2GgsW4UExZwL/KVLVrXQg93LSzVeil3oHHdPahAU0bpSwRznguKKJfwq4j3rb
FmISgRZnMY7HOnJZql7drxDYe4tBZpHUqutayq0jEt36EtrLV3A/BVf/MF+SiBIK
V4wHtdfc8Hbk0FO1flqIbmrHWYhrzrm9rE+Fj5NInHgwfnx+baeoKBmK8RW68w47
e+3n3t1ICSj/r57gaNi27odYp5WtyTfgREs+iFPMInUtpbwcV50JL4ikeSPL4BWt
2cTAHu2ZfraV7F7/6gmNVtPSxOxzXNQ9fQM+lvCNG6GPjwW3BLvibqB8lCJSWRrr
i4SClPYnrzQUTpGL1RxiEhieii0UuY/ZlR8A/DwvgYA9Rk7oo8Vl/c27VaX5VWOw
T5qRm1HKN7gWdhZ0LSQU4EkkundgDNSW63UUq8UzyQyH6lRhSFYhmcj0VH/G89fj
Rv4xlMkAZCSlCeUtMHb3W18PA0Fvg1GubYbKOoigD/YdxF1oFu1cHTxkme8ucgoV
DBS06tcuSW8KgqSHXIHbyD2VG0MdnpKjV1Skj1uXwc1MbHhLkz6/uKU2EKNPy2FQ
Z55t922Y7pwpan65/HlaD9k+EzQVvTcwGH0uD802YdjR5H2h1DxvUKE1ou8yh4xB
/T49oWnG6zSgeVDqAwU9sMBE2mBvT4l+0RW4FdES9Qhkt6glpm4yiOwM9LwWtMfZ
ZbWOmSdA0jA0MfQVSizwh7mBWBrvlCvHn/8PAZQphsAoOvaG8i2IKceGpejAvzvJ
n7N+YmQcgpKF5Bi1L4iBv1KQ+RlS7gVODwk/+kgm8GXLcGAGVkeC/iXakBZp7M6O
eecQiljV+qEIHa/KxdyN9EPuZ8eRdbabqAfOo7CVeQoC8XVI1S+MGucE9gwvjqdr
fxBLI/wdKxYNhQnNgVyCbvP0mznWzuRQqS1+mW6E8gFASc9MIk+QTSwHdfAUjYFA
RtkhKAQXFrN5BUpwMa2+K7gwz98v/LgUczWTdur6ZwDcUQ29CHn1jGcWzQ7/GNDS
g1y049Nr5jDzB5eo8pBqJDPskeEToirNYvaktNTmXMzkfWd1fuo1yGsxn4+8FE8i
T5HrvcrGyOXWFBP3AitRUmVdx5UgIDKV5L4oJKGnhsprMu54bcJLXTAhnizKZS9p
6D3RoMwCotTO2SmAIPwCjZ0+Om40a/L4kShCUKGlGY3nrtXNn9JSXuN2YBV3/E2a
JbnBhJ4nTDZVvU1mowy+xGBzjZQYM5pyfHS7tCPtmQHIDS5NOlSNA577HDe7hJpO
mAu4Tjdq0KEgHA5UNsMf+NkcDMCMo5/yROGKnZ0VJordSlQdj00VRONFnxD9HZhs
MqZ2SrsLaTdw6oyDmDdijmE9H4M0endUV03umYPKJXinmvBUzPrGKoxSS3wIyAnx
amtcs3fSVfKUgdjfsYvogQYlacjcj7vvg8a/YdZwn6usN0GD3xQnblT69xhay1CP
v94RHlsNRQNheoeWKts0VPt6SP1REYQ4wFrAR5XCgBlE+s0Kibj2lGMnfDhUSCWs
8vwPlgMkk+debvsEjeMn47ngvNUt0JYLqy+vS1I6/ALTAQCMfxxiV1g9jKnpXNqG
pJiql8xiOTZVGtUk6e11PJ/OKTkUMHyOaTSMeHVEmHAV3dSuBBDRqfbxP0wjIQHj
fW0XQOLvJb5LKz6nEOvjGfK2V+eU3dYkYEXv4AXPlMJqmtmR1dLcPsb6PNm2zJf+
EUbDr7C0OA07Fw9oaSjPI1x2S3npS7JGbZBmrmvAqsrIDy7KxTX2JMnjjRJy1fkt
D36ewqy04Xgg/63vIkeLIlBpicSB9tgoKeTut1L30Z17nxFeqgiZ4N5LBV87mHvK
t/R+0kaQLvauGObVKuechpRGCQTiF7PsVkUoZoSWR2rmm3+kASKO26Dt+8zNrXqJ
5+Tb7ZdWIxQkDrcuxD8I6VeEGYq+pMxwtkxydwH1Ms7X3ZijPmMJfT/f7b9bNC0P
xd5A/y+pBy+X/Rexpj3AOLK+KgEuCDjwW0bT9tdAJIMik2LsT2/CdIu64RK6Mcas
FStvzx5oSbq1bs551YvlmmUOP/cEib1fvVvvjjmjJzKLQs0mYos1adlWEW5tsbWD
u38nFNQxx4qQgnPbeAAKq3I1weslUPklpVBBfhS+zWrakJW5EzwdGAyLtw0NqE/y
TqBb1b/vZpPrMC4zJZM68Bm6d9uh38JbYDlSiKkovqkO2ymbhkVr4yzbf2W0Ckoe
XpzDeY2OMLPABn9C9K6EtIW2ozox7w1eeObDQFe22eEQfkkfPjfJ3NcAOv0dT/sA
aRPqeuS8SmYU24V4F/L8csG67lQFWgak42QLke5fQB0qR9sas1TrkfIry2Z0nox4
YtzPwyw04BHQd3teVRS7pnNJeppV04MdRs8n06djXSnMSFSxbULJF3uv0keyaJjj
f8b1kb1TaKHgD2dV1KdYLm/wQtyQIEKZdFydTk3QDOaYynpO7h0s69eNZa/E0lVp
Qouk9Qf3a7HdUsBfj3Ho5Sdf81qR+J6FFNbcCbp3SB74IMAWN6PjgMs0xay1aaPO
u+dYRQl6F9UUeZfPljUqFvYLwVIdgty41E1uL82VTGxauR2cRCKTuFLnBGl4+ZRo
+TzP/207OzF+qsTBnn1ymMEvnzlpd7qRWzsYVWc/Ax3a7SdMUYc70nRhM8kSADF6
1JDB4KQd9csjN/xLs90E+FA3pRGss8tOJED1acKBHj2IDCiwM8yGeWoy3uUVQQCw
ZmiPw9IfEpLETbDHG2qBQzlgKckjjqVLKnTj3mK1mdxpCc/XnO1UKbcrJX2F0EuI
ldGVb1xr+JqplzH//g2VSfYQRkFY6NpRkp7dfJjDTyHDPg/mHg77ZUSgaLA8A5Pf
V7GuIyDpUVLYhQN/UdW9HL0iqleoQDoWnTAqw+7tq/g3tjAxk9EbWGWvwLprTJAW
nH39Uk2Ok+QFgXTKkdH+gesnHd7W1o/Fk87WfjNsRvCiGqxyYDQxRWQAgrdrNoV9
dhKzljJPKimQUJiwtUxCePykzojYcdgQpEPtYD0ZLgk7pHUf4YLPKWWY/S+kZGpD
VbAwtNADIIxROsw+Gg4bhdo+/poeB5uht3v/4mB/C0tyOk9LXP39p1QBqbVfroFx
H5kbyqgGsJOUwkZc4qJtBW+N0KvO1HJOgyRfX/ox04VSItin+2YMQgc0XSWc4PAW
AUXGgYHVm8hX2iSj6ljcw0a7gLaVgORp5Bb583o5SV366BcS0x6wt5pqNkhXLpoC
ru3f5AnULQRS2l7wqpXsStY20Zh3O2ILOIrQYGUBmps7/Qo8F4wkbKj92XDd4+jc
J5z5oiL+aJQbKdymvcMpjS0mqVK8800MwKJPnXRX82kjhzP40EZOmcRdwqZF+7d2
BHVuy4fdaaR1Xz/KryDFPXhTsiRkRyzBmAHFskB2fh10IltWCfePz2DEopmP0xS+
E4iyAUW3ecrQ2p/bGci888rM8nJOzFTa4dj3ZSwFGOBKwYKz9HMD1PwT8IbbOwdl
L17B1ssXxah6wKOq9OuXG5E51TVeQzH0G0fOtHAV5OnKiplCtS4Ac/hJFSt9ckDH
/ocp3nAmCTCjitfNJXxGOYh5NbM5lgwstoyNS0zVzU66ce4ZgXQDANm738BS+nYk
KlU5wUjqEQUrgzyHtMU+3JvT2rUMhzOph7uebKUNVCvNJNWI+cCAj7UbDvYJSM3t
AGn8uoz8wQYM8u43kAniWiQ9cZ6AbMKgOz+FIV1iFQbXI8Ozq3+iq3g3aQyLnDg2
eQCElNba8wC1plHeT+FM+EyFmyShFD/pCmOjnL4dtsWVlmaDfRRYHVfbcsS7eefH
/iKdlsGGhIkdx/I1hjRtOjDxN/n5nzDsY1+VWg3JQDg3NtgKEBIrfJd2LiVskgR1
vFLEpyMB2dzO5hQSZviqVfSnSB9KecrKycRuV9sxI9IBvTNi9UqW9nrkPExqD/JZ
Zwm6qB5zipQjHYg2h/ny0Uff0L1zlaXDWh5AxA8zodruBua07vJ4dmgOUwSceHn3
Z9FyJjRdQEhrs+CQnxHtnPj6H7Jd7Q3czqIMwO198mteKSQuPWl6LpfsSkUQS2CJ
3jISkfM10zzxjRFfoorgDyy9pDzE5wEGMTy0kYXrcIB714pPAu4q4ZOxOlFgmTRN
bpbUws897dTxyzHpG9/s+ioygnClCI6tA7gyQu5mO4SEbedt3swUfvP8OFWNoICU
6Y6jJ6ZyRlQvd0csIAZXb9ezR9kgbzTcKlQl8EiZNlYfxu+EMzsH2lEItDu9SOzk
YTHW5ddsEbiU+7JeUyH/W5eORBXhVYYbE4gnGJ2UgQtzwKFdV//5m8550LL92Vi/
pItYtocIRDPNxCFRG5d5UYmAkPOwJ8HIfKDOTgqHjTPLpyrP8E6ruJUx0K7MVljj
AfCVuiTp+jquUiBetYUYnlYnwm5e69zm50x9J/FKdYX1i1ktAE8l97gTQtgJxs97
ef7Fg2jIDiv7uBjLi6ej6x/amNC1yTofd0nIngo/V1OlIHsFuGP25j3KAevryMyp
xv2e9vxYFGiN+XKKR3ijae8v+d5ig2hPTsGMr8KvWjy6NM+M87mCZg/c/Nq7GBrc
89KhPXn8rVyuGeLWfIut31rBSYxamX9qd31LnjcKboyNN/BYa4FmWgqMCFxU30be
hgc20+HRrjZzEUKHAJE6YCmdQfzzgmnetQ7FEHnWGcgrVZsAcwch1DhSei0wSAgN
TX5bgjVU/BcLODYpBHYgMybwYcitkygCyDXvrKFsRcNlkLljwS3r/lIGMvhKolFw
aNMwhXB7/uhnwnICNyLnZsklnnnbHe4GJ89c/GnelaD4FE0tTMjWB7MYpfkDxdS2
YiT3xEuAkvoDBZ40Nv/XuJeUNeMMSQgLTxRFBFf5E+7Arb5Cp8KEGjYKgwuayH7a
LZP6yA9s1G+yrw8ne2jz8QeN5KOYJnlNM3B1nHM3JvIFmJEeIF+m1H8famqPu/oa
nD0Ydwe3GCXyRWCLp1ftf7RAmce0EAocDnzgMcPr5WqRffpiWh8AqsUeum2hXQhx
7FsCK20MR/zdawd33f/83Lc3XUImJYO6iSlZhocnXh1gHODgd6ZIZg7XQzuAzHMI
a4kBtPg1se4Jl0sIOHgYHM7pddWwFhdpxxHw7mZXrG6cZPOnY2XioxEZRfTBfhEk
1odwHroiiYUTqYzLPPVZQZ5cs7BB1WCddd9mtj533Lt8ZRZ6FmVCEiG+KFzQszhj
NhkPQH8JLTyWD3UKT48wxF02XN+kaQqd0WYbQVZA9Z8+lS5kA9NGWd+8MZ2MrRr5
eBKb0PR1XoJCQnPe5RI0H2aB9hmttT147qD4bv6yxfMar0rvCx3UjVa8GBJoOQXI
Bkf0X88N50GUeofk4gvcqQbg9NwZoDfNUby6rmm1qHuOnzvIMI8V9Q/P6tlWlqfe
cCmGdAgxq2W2ycV37wQg/fQfkH7rVmlfBJruJEVivl7OjgLXnYjN4EVrBUJNFbnd
LkE1tqQZZWKXb/rYg7RPm/mfTw+5xPk2T3ACVH5jS5cFtXjIt59bq0FpTV/FrtJQ
x4p8u3Kp9BXEcxE8qB43pFhmsCyqPFGChVFpsc/DPO2ftZJUtKAEaSG+5A+dV42x
WppgduaEQiwa8GsQ6LdMHCHuSi2YYdF2q076prw+l04urSQY/ev90QGrdQIKa/Hc
lDcGllTwNCrhNj67Wem3lrQikGj5lALR8IakIx04D3MM1sIh65pFBkvvZhVdyuqb
rgHQQpdcCcXsboCYXb7d5/P7OlQOQvbuRNFVbR2vgwH5s9E3pRXpl8ov062DQI9e
RLBe/JbqIfTb9ji+uSmy2+wgbqHCNeC/J2GdJC6UHUi2u01V0Kwhvpx18t4Quxr0
Iw3anbF/VppxGquY5/K0VqRlnSV/CNwe7Fkf2QUJmIGvT9bEAb9tqhPaB/8CJhRt
jaIBapmlhs+DUKLNY4EecVsriB/7GhbUqZpXyUVhT3fX8QJnAsXJdq4JqZBiFydL
1tuKMVHaoBnY5QS4oHKrU4CTsEpO1GYGp+h0Uamb39VsdR73QtQgpejUfyM0SFLg
ts64N+an0jzlYXu2x5o8PXvNtDGrVDgicrhlH3s4elRXPLnawm5YgIsJzwTlcAF7
ra1/FfMte3g+byLTEWby+6sPYOaP/LQLCRJae31kwu37BT3DpE/V5nJeBYPUa7BF
F5Kr/Y0NiBgWSvpWvWxPNcqwk5N8oUSNLd+ttvQDL6phvBZ81N1twZEPtTG8OqTN
6rB9CBtC0UFAoV4WHlJ1R2tmFl4Zb7tvuSNijp3b4Y6JkaGP58qh9jxiq4UJyopx
SBx4/XEd/OP9jk9jFQhUxJOepraYY6bMOS51tdde1C9uwKvVBY3HHvuMzkHLTW6O
JWkF983p0vJzoPOVFAjOkQijegD02whpdKha0ErZGhZwQsV0nnkafxrs/YrpBFmP
qltU1okwMBEROmF+nKuBJRds4BTJEOMeVuH3srS14y1tLtox+rwSStaIBxWwsEr9
fmpUudAUO+hptOzR5nwZOTkpeKByyp4QXgefEtbpJk3JlECgf9FnOzFxvgSDf4qh
ycXjUZb3lGgKRUrxX1upl47oDkqpGbUqAJNVfNGT4u2c8/hPQdAu9BY3Gppdhdj3
BJYtUiVYeuAhXiMKcTcDDDK601wujnt+K5xJ9I+PnVpaIR8o5bsbMt3BA0Z2hdOt
z4EXFRhv7SNAj1D602DRvXEz/4bdU4K+zPHe0WZ5Io42w+BdwjEyPJNKcRNjrgNn
d9Oj8rrjRPH6ZstIyBvvuRCuBa58mkZlE0lZbDG0sLAYUWcWXsU99rfMAC8gtIDO
O+4PdxHQAjSCXkcgfF94Z92nknuSx2Ti/bWsDUVRXOz7BMMYMeEJ3e1K9mHvTCRu
hubbgR/U+M4tNN256tvNUEL6HQTceyhI4BuEMCDQDytBxgVCEiv66CUJUNNowH6H
MrWfdfWXxrQzTqX97Fwn9CB66gNHm5NSjFFYMbjXdgms0s9FFZjC7KmSY5dfOdiO
EX2F54ouWUbOOs8xwYvdpd5QuhqH1pZaLKz0ZzXq8Ar/K+n9v9AZ2xSH96MmxzXE
L0mBXXIiKCI8r+9p244kCGFcXzSlSZfB1VqjP5wYHHjbe0dS4Ze5DlJX8p4tya6b
F9MXcpH1qdRCMsEspu3lWG96GrwMyCzT/p1P2+T8Ov+QI+YO2Zhwrs8UUvgJXqCU
CvpJ7o0AXdBfi5Xkc3LRGZnYkhB8Vc/7BnrvZoL6jUudndO3gHRwxXr0Ryq9CUfB
AVTC/1THQfgwS3zT/2VqLhLprtTiNvZRzBPoB0Zkzu/f2cgrSipPxZJP+XUU6Xk4
ucCKgILEPB+eWjFJxq1aZleBMCJNBSx49jfqbDF1fUDfxazZAZN0hw1oOJHHfLq8
3iBD1RL/CodEufTHY2a2rfXfSVg2Xt7gRblys67kC486E3ORm2AlyOi7uj4Yp3k6
VlJLqapLxfI2Fal/9z5Fl5CaZQ+OPZddTLsIfZ014OXvY9OuApWJdvwhdAfHD1B+
NJHrU7H8wsXGiiU6pxhbHhknxgMSYmzpko91gnqoCgdKMcsHRWSeTPpvTbiQarZa
oPgmVgWDUzb5E/7nHkvFswvl+lW/D13KnLg+UMY/82fxQluLSzbyAQ3OwXmZhrPR
jNsJWwcS6PwtfbxWTrLGeBVF63KFLXJBjmlAIsvTz3YYF8yfF3/9xscRXq41Zn2c
Mf5X+6fteoKbT+4PxR2GEQODuM6ATMYkTJqOvDZQNVeplf+n5Z7S5ZIKNt4sFKCV
2y8OphJ8QKp5M82j3zuNujPgu/X8LWoPmOnzyk2QWgitg3zfiWBeZ79nzm3Va+U1
cjNtFzFwKFEbTVViCnbR2aovgsA8AW3Vn5Tt7nkJfq6JHn0oxY4DGiSSzDwL1IcZ
atJno3PayIcfPZ+sF/qsPHpGKtSHZzntmD1xEhXGqroTFr4guLunxzr4Xux+n8uI
YkY3GZLRMBswxs1sihE03C6ZZx2f1j7YFkVWVkF4EnOdSPEkazqMi4PzNk0QguWy
gXWp//zahJwEaQXFQ9W0JYFl0hnaxRlxcD2pu1cFb6X8O08Qw1CgilclYFEtvmME
5wcUA54ZXFGUxFhZDP4FKbrfl2+3Ywhy9GLpX5ZVto+xpYyWwBmhcjS1TD44oqvv
1B3XaG2QY4HLM0m9nCfE55i2EewecFzesGvm7bAkLzRJJm5ouTcGNdhSxi2z3HBm
AxktmaeQYIay/FqtcwbRAfA9O342mNgWMb4p/Duizps8g/BToMz4B9nydbQt9gvP
PVJXuOltMv3770IUxGTDZwp0O1Eh2GjvOesR8rVQT2BmuPpxTEVphJ08HLjS2WRn
r1oV4jApXs60DRjABHkhltIIIH2Uw5PFdEAUbZzH8BnlId5Oufy2+CNcOcWnqNA0
0Z4Z1iZwb6x0CR4A74K1k8YV7MRqNPBSK5A9sPfd/GHRubG55k9mN/UYMNdvUWum
HKJl3+jp6pqt2JtIfVS58wYjC0GUrxxSecb9wJkpEDboUZMfzXvPGJkqExFKo9Ed
5kme9GXkmz8PHqIWK97ZUkOPMRdDSM06hPFSLlAfXiYOfMAjuR6Qp5JbdEH/EZxt
KYpeG9cbTChZuh8dj7YVv4bvr13uytLQ5DddKGk7n6GXut5RtBuM52Nx4Ol27nl0
HvKGb0KYpbtcoBtE8Qmw6TXFlYvWpl+ibSfWdh6ZViA9VlirLEcCR9HvBalYwhyV
DQn09EsWVlVyDBmm1JJgvP7AJ/a2/8bzWesnKbgaqt7UBjct+3X3BKyXyi+RyUoB
wYvhNh/NUxO2EcnBkyRwq4graeTTMW1HOG6kG3U9/9avIUcETfezQdhcpJSyyRjf
LEzgBhqE3QPc9dCjQ2Y0/A4h7iKv4jp5sXgwQKda1xLqVPaQZNf5cXUzZxVHM01L
vLpPruBfvqHlQjYH9ecNZCMv6frcwHVDT1HaSdTmPT0mMMBreZKod86WZQXXOgCm
BRrbt/oe/q6sdIlITCG27ZhbtJS6SzgEjMhBzk6ULP3O0jOPxrF2THuFtD3/GpSI
hNJagRr/mgiInvhwUk/Axtxwe5uzDLtqnts5OlxARtg3i+3uOLWLdmZn+Qm6EMBk
R35cTzbvCW8B19U5nmfsJK8FFF5aAYrjr3FYLPW66SRns31dZH3+b6DLEwY+YwTr
zWc/wEMZOIt6sy5EgtEr0D2bFtLyQTf1PZ1+dzY4+azNuyebsufpWX8rcaQl7l0i
dS23AxWdZ388tX6xLLlb1so0xwbM//ferxc8IpYcGggNn7PnPQ3WBM/YEG8uNqDA
OgxYtXF2S88fhu7qBKwHxm7Ozeyi4KafbRbAFE0XGkDXDD/fWmzQ8dEVV6g3GtMr
FCV1IJKZU9MbNuXhf5VBCJ36Z+2WyG7oh1jgVPtPEuD/EOm9KSqO1aZ3DomLnOVI
/A6DSxYQoN9uPQxsejmXMilksbx+jdT3Lz0XN5TYsY4tfvXS3PnUwN5gvh/6x7qv
xjUy8NcOdHm2+yj/CPiXXiUhiQthphhi3KDMVMocZxejVN7tEyRbi5FivbsZUPxd
MNySfk6BMKTSc9dta2C7xcsP6scUGX3vl6NW5lSbs2/JlYlcjD9vkJxfcuPCnxq2
in+TFn/fRAsc3M0+x8b8acEgD7YhLMLr4kmaz6GZxy6yKrytoItyYpboUdN0NpYR
T4QXMPtMsoJeMO4mX+DX2tIfRdeK9yGbsbFXqSyobdAg1wOCaPTPuFu+SM2nutok
1Zv+gSJwIY0nSI6zuw17PBbwS1KSk+E5a++jtk/lcTmz7FeoFNulsbfSNN7rm05C
EHPklgAee9UbEHurSYXMEVX6Npf+SQAWSCZd3GAmycO7qpDIj8EW1G6lODolXXx+
t6I2i/Pfw5M41N8YaQFv6m7LfZW8jma6cnxqcNluRVdMU/Kwcz+oVs7UugdonFjR
ElEtLX0oXrAapXQF041zs/4kxohux7YwC6pMEY9fI3svjCTTDQIuDp54tepYo8k/
a/5nuip0V0beS3Rl5kfIlL8LFmJ3ZS91uJeLa99GbnapbO3imMCHNlboa5hfvQ9z
11IbSw4oXfBXQ5IrOmGQZWlrPc46/dCxVmlksp0Ip9r1SF59uK9zFDZevI34y+Pv
zCCQy6NebNqhJ6/wy9vG22RUW4lkM/naJJUiQD6ar1NHqLGMEO1eMbBYNxUG/LER
EeUTP8FMEaHT/irMzsO2fWcqpLaro7JbeHJubg2e1puNd4qUFgghXSI2Z/dZ1ATj
qGEY0CVyZWTITmInPvFWe0TvhSKr4+5MANXRKrXWnwTITirk4eNLYAbnfI5r4SLe
Tl5zTvodvPoflbsHewWdda97DMbBmKznW6lYM8SHg1T5tgDyIrOws7ZT9uPwmr2R
E5a5gNbEGg5ma4sVWjKFKFfCy2rP/2b4eB0zq2MwfnT/pMCjNpnhF+RVk2R9ar41
9omWXvKDAKYMx08DMoma7inbdNS5S1+tkkRKfI8Nj5R6Y+VEzYVqDRiyzng5zlHf
Qf9Ue7IbCYZw8NQ2vMPP2eYRbCLhqsoJckojU7aVM1FS0H59AgpkgY7nvtUb4BEA
quHy0KVwiFknA1sDTRpspyx8XVHEMNiSHIhUc0+XuI+Mmu/DffDZR3qLhKRCO2gC
zKEcQtTzpzCOUh1imQgYInNkI4HLGKWIeZ2AyL+b71q5SydiQLMWC4T2NscCEDA9
4PHveSaez/xshJbR+D9KdWyhDSLE4pRCGvMLvZyJXYr9Xyl2/ZdsmqZ0w4CFD8ct
FEL0iF/7MeKJ/EQQjyR1zqQWgxoCMf+kTUUfjOsPWskFKvm3wRx1cEizTZd4fHvB
Y7ex1KKU9qrS3FKNcrydHkyWa85ko9lSzk0BTWnjgptGpjAo/XzK1GwSlSjaxpn5
M9J6ytKuseAWusoMhw5c9MWgloe//kNVCmIaUVVtCV2Gw00fDfRTqYc8WXxIYIWY
KYeS8RidF8DYSDwBF3julGtiS3cJMvp/7maauADng8B7PYBwfkqDOhX+mYX7cjO6
yaqtf7Abh0j5/SqTd2h5hfn8hYVMplGuY79XCYU9el++pOeFfdG1WNYaMtYPOK7w
VDqd/Iz7vd0AuNnniSK5hhxEyJZKivyg27MPv06fRVTzi9JVbkS1lIrwaQH80X0G
kuFujBWSl6cXANBi1BLJH2efahb6/G+YClYfSK8b/tdPBBw5Po3XjQ1PqRVhVro8
gW0NZrwBLjCzTXRiHkiY1orVvV2m7tMXg1x0r6CE5y8p89nXPzOWr1MBmtPZ2xnn
eiSd+wcKySSwRXiEPSvEz8eIJmnmZBuSt1hSOIuH9T6cBDDi+wM5SWgu8nnl1mIX
g5fBqZFXLjTrDMrYMXyi5dEIrLjIrma6/Q1QeKHOjPkXpc/rPilx3T0cDsE0z6Zo
vqF+Ees21f1NAurc9zMqBeRM1JECJ0S+Em/F5I5qRsVrsraS4gdC82DfSCcbcAuv
N4rVjZDCM+UinH9iCpxBmkwfmd1jkoGQKiw064iUNtEVhS3n2pWuer4QSGLsi2WE
dlJwovBsYlXI8Bwf7xpVq6iSQGqsDyPI6DRou2diAARLDejLzQ8m2kTEOJCmGhro
CeKPa1mOwJnQdk0qQ6xLYdxD3r0fB/uCO9N7LCMuwxlr2xlBy0k19kajw686OqmT
Wxl1jTK3n10sFF79dAYb6rEWDKIkl73aRLZAnY4CbSD61qaAFQoY8rPhyd2bwmTx
BJ3Ke5B92NNqMpUlDE5mXGaYxB4/TKzTHMWa6Xrh1CKNGjk49dChDw4BTxkIla33
ChKbgz+zAVQWRgL7tZXupwsILN/C7bl9ghTBkYCm1AfpBlhpec7ik2N3JmnKoOle
tat27MAClRXbaycTaJyVdnOgZC/FW4QwqCM5TZCxR/CQ++zA2s9Rq1mm+FOSxAr7
Koo9/YF6DqO+FKbYA8c6jr6wn09O1aNEeJXr3MWdadFbXNyPPMRwFOzIiE4DAWJD
vM4MYhk436OtEJdM+XsNfw4Z8xYLs+FzzXBQ54oIDkuC73ri44wTaOi55IerjL7I
XQK4RbcFT6dG041syY7f2NcJeefgGsW53ZCWIlpgBEP7cwkW2zLYIW/B9CtVPLbc
Y8wRQnaBTG+ezqb9u9DqfcaXCnmvHC9kCElN1aQZ+KyLkjbXj3S5FtxFQi1yMHoF
W18qaFSJXmfzr8MhtJglaa1leKfcX7f4kiRsbpVzoMagkkieETkagQJTRgG40/jw
Tt2xw06S+jlmbSxGjVvFbmDebaMkIbbLzk1suZW2RZxhFoGA99IVxjVRZV2+t/Y5
1lqqgv/+5btbBk5hLx0katlwfVkdWI8++8t1xJJqHNBpfsgfEOAaz0yataVWNBrf
ssyfyyMLa9HIZeM4sJphFY8z95aBJANCu1fYPBxlfzfMULItILjhwc9u0qcIZ5Rp
rpmy+uBOrUh3jWFC9A5NwUZe9D16qlx/WdAMr9tXvJ5RAcre9tNALY0ImUdPRgBI
XeuT5AInUmBjJmQAM06RgsiboefvTAbbEvGkqgJ8FCqMY5/Zp5pKVNagh6Skccx6
LhVmp+hmdP3uI2dveXlrusobomDoRXuR+FJH8lygoaHNFfz1wwbsJpvBiOZ9/n6f
Z1NWkhfvR5a1mpG7k6zeOC58S+vdxwkVddazUuB2dA+tEdKhryqu3JDtl9QGtWJb
orzXLgdU6FVwGvDzHSLRA29m3XfDObo5vk5/Uc6YgrTYJXEw3Ym75OPA5asKhx3X
dXhKdq/24L/RVOKPk1B4ME6nSSWtsXQ615eMRmkNYFoFiHmL/tUwv2HzC6QDS9rN
kaICrSfejfN7whzoEkd2vrSNbPnmX6x4un3X+BBEPq0swhWRRe5DpXbPwlpjMk25
hc9UUgqACjsKLutPAfDARglGNC1bgpROIogdA+zb4Et0XjJyH6HmxdnPNiK+oPlU
TweEOPpYL3QnBIDv0qxMCupRWH+pqR9I9EeoXtJvqnocNcBQ58ygEl2LGVIai5fT
Kf3CgI/bDsM5CwgXalb+ZaO5MY4nCA7XrxOuM/yVBN5Zpidday/uUaHFa4mKa3zL
OfiAVT601ojpTxMGt0MxWkcr18v1N4DqdDAeQc9U5F8zY3QoNKjTj9EgO4vDYb/m
BiwGU8NiAGHft/q5dnXFaoYjtm08xDK+QByOHAVBlqkBgDhnWoKFmp7e5Ub6knvX
lzvcpqyyOCn3DLd9I729b+H0g7/kqS1oEQs65dpty9Km187XKfPN/MVzihs3U+4J
Y5Hm0qwKzENd4srpWFtS5UH/Bfu54Jm1Dhn6bmqsZRuQyVYtDI7PFnVEa1rnhR5m
OMiocLjrmielDd0+I8lYKKfsKpRHlsf3MnCBHjsxq0iGs+wYt2hgRflWxgqxrAv8
lCQ9iipJbXEDd5MbEFDjFc5xPMPzuQ8gJJl1tQw+QILVrv7ZovwWYCphO48OM3jk
TT1/XqO3YQlH7lNJlYFSyMla4nLBOqgQXCSLiZDpOK33hYUx4ouFYGmBSP5rThce
q///A2OIJmDQdkSa3EHCpBsSTa1FU2wAdz3ZRwvBL5hIwdhs9kCj8Tcqpw55qNk7
q6koLrET54l4VwBN4PEnLzeG9FJLL0pKDNv3L2/rjItx3D4RIEwvXKYgL4gPQGro
KtD03oAkMyOTAyjI/9WNT8icUHfWlqWAiid8Vj/TphYPpQFDYJzYCv2EeUSDRE7i
0Lgwd9J/EHwPD/RflKSOcV6s8w6Lw6X7uY1zGbMpO+Lex4IsdzneTIoBLN3ITyq9
iH84zqMsic8kX56kZ+910To2xFCanHoxrqf8SRP8W0qr1YSe5Cx2mwg4DMF6R1sR
9OALwfgkZxMbCWekUvLZvuLt9+QHJfQmMbYNpKfZGLOnboGGoDiwLU0foGdMc5e8
QkJW27LATZtarxKjDf86zCB4K4s4bDEt819eUAOSVheR63iD7hmHfqO9vSEv33wf
56QKngC+0qDp0YSSIZ/2x03pn359ujSgVzUvnGufdP9ureCFKCBlQzcSoILNjOPr
6lWGoFsCybKnB1juSP3uh5YJ5cUV3H6Vq9EtDtxdV49MBuCqOa2FdB6ViNDTICHM
CXHbsPgbWJJzz1FYhThFMV86U1CLRLipXpqZHc894heOSURtVnK6Q3oVrl9ALJNx
LtLKJXbT5giVoAjPTG+dCAj/kIHWNYez9cdUdZ2lfr00NHH731raS9apBunf2Eh0
E6Nfr0ct6yYnd7opi7Jlc50aw3yfALTyLIr+Siv5igDxZiG84bEDWLb5CNqEoK2c
Em4R52pQoZDU6YxYLxGY0MJwG/sqSOearIp+0hCg8AlKjIW80MyfJEIm7BnybGMC
h1CL3RSE6DoeHzwegArlpZa3lxc0fUZlgVQ8I1TogoqLuz67PwV51vGjFNe429t5
BTSYAAKPggECyHBZ0TfU7F9VcziCIdTd0JpKh2dloKHko13QA1rKJFf+y3VViqIF
fdtYJjyomiRtPD1+kzCy9KOQ4rdQqCjZqS/UuyjFKR2LQXVUURjTRP3imoZGuWaC
nRLeF0MtnefN4qoNjHpLRw7IE7EdN+cZs2jlhArpRHCE+D2kmaVXw6SzaCF2f71r
M3/hU8k5YUm4mzscISrAQTa8EoMyShWwsHTjR4JeN/dzGcijFuyDK1hluG5ol/sU
kR6HALH74OgMesQieR7B2R/f3gXG/oukHxuSwx5pWS2jdtc2Q4gR6LZtmD+j+v6P
G13ErGGaXmRtSjsPl+D+UL63BgMPSCoWy3gvHHxz9U8ZsWTxgiL6ShdLTO82Ub7F
tArgJG+v0A2AJPaFwjWgoif2TaldwEQCMG2RCH17bHr3p9NZ5thnnLQ+WmAH6kQ8
HtAupp0QfzELu9Uf7JDYTCbmTKdaVFDYxpSU+AAiNn+SIxbWnwBQE6ZVPsZvUnR3
4QhD0zbCwMGnDW4u/fWDwU1pR1by5tu32MFJyo+oAuYmLxm1epPy1t/2+I5fL6c+
p2Fq+c4PXlEvLluGsOyTaD+tjBOMJgo3NlkdR7wTzR3aeQ0Mp1AyHFBzE3mPmmjN
sUzKG+AZ1msks1nUPtgpLwORpT5txBZ5frC7xAf+X+o7OBzA/9PdzVY7mvrvMUq0
fngIFHIjfB9mFYQIpiLjODVYXGG3pSD4u27ekp9kRX4hRqwYGjp/Kj57TOocGJNy
hsTh5n+iaNHk1Cae3cZglg/gy3LHhIa4IDli4fiZUSDvR727x3C5GghutwU11v9W
Tqf044L++KOzygnunrqpT/RbBrVa4p93aveT5p9t79Z1ovV38sK0doLiIWlAtj/O
00dFTXfPcnJktrODuwijrUECBZ/iXj3UPuWizFjIo3s0cziY1w4zlmCpUaZH2KJ+
ogqEUJVc07ST1bxc/wKb4R3M2vXCVZZ7zxKGrC9SAhFjrmQwG5gcVniP1+5OYQ5h
f5hkDPenYt5Y1HW3z9mkuTldTmt3lgNmSVTldWPsO3d/wvNl8W5Mgw0LyX7ANnlY
D+GuAm8N+odyz1pizwfq/L/HgIeF8rJ9jEeP84scSS/VDZ6cIpkbY2pr8SFx1IDv
5bUIl+AEPhfFyQbhfGCAI7HaukTFZO6pTcQCgweJOepKWHVsn9JbWa4rRhfjda6C
H4j+Hy4KJMuu3kUj+XPClT03tLP9ExgZCFXJ8vo6PTcn4SxrRZ3lBcAWaMFEBNVZ
jeGBfcsQgQP3yQ6qqml4FbGMjDQ78No/X99RMw2uzV3VXjfqcyPy1rb+TAd6WD+o
gNd1mpG4zdqVMFSsjH1aRmEKZHHORsT8s8gO6VPKtEwpZRt6e5CkxuPuaaUT+HKI
EkmdEJqp3VVZ7oiVVO1xY56KaMG+zLg44RBgekVitrMUk/OW8doKkuFu5z8lnM5v
0Dl7wsmUnU77aB4j7FYmmcfPNXP9VhwD+qGCRyemHuDVnNf4NYClpM8LnNwCDwQ6
XaONnxdWm6bj7HKgw+tKt3SWNRZPYM5JiHS7xBM/JTPCxVf7MFSRJzOPI14RcZdj
8PDGn/4FPc0Q6lAOaIhcyBSh5SSyozHQZ1xLd6GEMVjzK4yVgtqUnA8En7kIzPbu
lApYH8cBHc7G4xMWd748nKrupUNuHWnE7p10tBDKdUKVGiGbfJ3n5BMYQpJulKkm
tANuKP30IbYpdqQQwo23ppeEb19EdAAq/w1ewEhc9ZjPLmbpWuk+PqkxL8QKZ1O8
uDnLJtkCnbLUMmbd+k/pV9/usEr16gNloDF860Qp94O7bGhOUnXGVHKsQIjjSTzB
68dD/RFauw4JJ+SEaUBMseQc08gFBqTa7vf9OFPRPCVUax1DF5zS/ygLCpnFFNcm
2EceSrjqf9pFfuCHvFA9Ttvl6xeyfy6EriAvSPRHETl1hTuy6lRTvMvuw5R60hCg
CFr6fof9LoLYj+IQ1yGCXa5QYXl8DtlxfCtsmlwS1Z9PU7l58WwJrLYeUH0TgMOp
rKDylPA0e6z3QPUAb4digScg6mWGuneiKJ+9XFQ+KH0Kr0mvN41rjW/TaHpmpEK2
EDXv7iAsccwJ7vg84Kqta/Vh/inDB4TO9TDmKbz3sC912TOlpHYgcmO+bkA7L6yK
+eH5xWOGpqChe5KhUJ/rYO0vUEYqXWbY1xEPiRUjSPvs4i87Av6FO02S25auOhlI
kQYlYFidNV/zGS8xZngusSW6ZF/1LizTVCd/6wgOE1pAlMSeMIH90g6pYWeeQ2aY
t60+seVY50GzXQwNx4t/RzYHilO9AphBS+2e66iezC/nl/s3snT9PTfsTJJ07swi
7whoOmTVDTZQTMasCW+qOlOpl7vBKzxogRW0tl/uVDtfk3tXgrpy30En3HHySoxq
nLZVhXbUAzKY9HirjZyEs7KT7keB5uWhGVHvfyaVy7agKHrpeRuA3uCOZFQVJEyF
FUpgjKnej6crz6GBDwW7usdzY/MtGxYInoWaf4kdgqmpyeDWUvQX1LTVbuaDcNoz
QW+6L6aRFnCLr2hNZQ1DHcU8jN7eBF1IC8wKZEHEWguUNVhR7o0Ie3S0CuSkH5QQ
Oj8ir0op+a2SwGwAhC3p0OFn74tvPcwv3WUfQkWKDAb/ydHU0F+c8itbVYQcAPvO
3r5E+gt8eUVQjviQm7Wz5/v2HhgN6tsEPhPP1JFpxy2N/cl+HTsJP1HhTfMe11KN
kClIWcYDsrNwE08IWGTczV+LYIYwAJWMyEwy+BxQ6AuUNMa7Y0X6+vuguynsNEvu
mugdmNhE8Y8XohToE4a7JNYzbiHjvBx9eJeEYHfBvCVRjB2o2zRe5KlzC6oD/Iq5
6OJipb0T4IF8ijuhdidbKKQ/inbByPsLT6Zn5Cr/r6fOWFVCMnYYNBB/WTtWsAcr
NYMzWLpONpDUr9/Y3G08MFJFK7Mv5/MzJJ6oJX94IIV5cJpLmYyt7X9J+dYfWY9z
r6P8lr8S1bPtjyhq9Eo9/naOe2o35Lr6t1gCk5yItM+v8VAzoxksGd6QgQbc3XJb
EmakgnfQm84U4b6CLUOWjRexvCPCioWCiLd5knO7k0Yb+q8dPUqCYx9ECpvAYEJ1
mg/Nexk/qdmT1hgAaDCeq/A4WyUr21wIbZRmoKJsdnC0ZIWuVkp5HKg3ruPmeEot
F6MB53+gpD2Imksh2Gi7Cmxk4uk1NA+qgDr8hOP6JmjRSeZHaTNrl/qy0vSysxIs
H8zi7lnOIOVu8N4niugCgTWDrhzucGIMDDaDUivH9IdF6w25Zfreo6lvLXfnpFek
3EHNWGbjXZJj9Q98HNiuo8d955sUIrH8o0f/HiEj64MoBhi600TAT43SomCKCPUm
innoSAtq72Z+9gAjIhX9WzeF/cSfwF36BOPdQZa2hqphJHZ9Di6V12bj5gnzj29z
JX+N4jlbDAFB+XrO8wI3mLvwTGqllr92/3cdyaxWgoHM0/diTBVPUcwkMZNtAkjl
EcW6RzVX/pYwLPzsHPEECjAxfU3wxgqMCwcRUPsdKNraD6x3jz2kUO76+whaSSVm
7oM6tMIsYr/K6gp7WHjUC8HACnGH79fHI6r+FAzi3U0Q84rUvM7br4pL8LY98WMW
A8G4ajvlunBKqrRlkv6/z8c8U1m9mvjQocg2G5B0q90/BhoXxlCbw6ahePJ/QMAh
Rm8kWaNjWdGwNE5uxoAQepAs+zRIAI9NKPZIS6waN233JQEYxZG5ZwN+QXE0pUrb
29EORfgPThij/5UsFG5HCklR4HtWL0dEyRZGX0ojqlFZ/jSquoHS/lo/N7s4aATG
AazWyC9C0TYOTNBYtpWIAmvGnF28Ps8YVjhmSBRxdAvKk/PqEhjJ3OqXLORPleJM
PP1WVYf+PDEVCVVDIsgWbGwl2211hJyE2pO7eiGhty0hj6aZLv/USEb4OTOCOhXY
0wFTsVjR8nFgs7tF/hBZ09m6gdVBSu7ZWx7hIfsJRRy+BbBP/Wcljf2bUQX7a8qb
Wkl+nN6iyttxixIpPzzKDffTEwc057nzoT2fIoaJHEZGlTfuE8kKJHpZFFdrUmrU
G5Yrlz5ZsNlXILivfvxwknHguIe2erelxj9bJz7s7bpkzUsLeTsonIGUCNy54duP
bito0Lt1sW0YsFXMXAO24RtgicPN4SQQ1I0wdcQCtNRYY7hHyeThbGRRKa3gcxUB
d4X3zTwgUOkq0EOzAI5yQ8SA9YQoNTOaeu1114ZubH2KXjf7MaM77j9Ib+Q5d0Di
BmXxcak6ikLmORwGi+JB0jbTIAl2rNaFwC6NIjYoo4kvMizh24V2wApdn4jS3CO5
A1sAOsrYCWpmcWbbepIFjjwkwR9LGyPRA9+CEvx9R8HaeukDy0RhvPjHQ6rUIpVN
UG5RK2vrrzYnr2qeDlqSbO9VAVmylt+k6/G8xxIkyjSl25LzaAwZk41IWEdAFF+i
+CH+bf/QElf6ystHv9eKRKuLZ+Tecp1FlfVBiWtCju29x2/nZD3GohmHBQl3ivcB
lw4zmg+FdZFlk/OnKfknJ7OuPf6FDCXSi4kOa1AsTrTGNglllkiaSpt593X6S3U/
PEnv7NNpE88IvcjnZ+/fYtqt9gRni3Brs/ddca0JLNt/5MhBcXCZhR9IhjJRHwoq
8A1O65kKb6kfdHeT8/YhNYPtpUMilXcdwfDf71cGIsMMv88Zs9E7r02Oiaql4Qd8
ABBahmxh/Q/AUj+znb7j3ulMm4IOkMPxGUugRqCPrM9RBEytRWQ6MYWpy1Vc8oW+
C2/lkzer2RjXqZMLHST3ftLwo7uZ7cfE3WlrUYA6a4jqE5iUNzvuzyuEpd97CyFD
Illo59Bq4BpSAVeTO/Sm9ghtfeCttmvS2hmn8ga+3eCAfDZJ1PNM0+7AwGHoT/Cn
cEYEc4UZRWX2lSYQW8PP28mrh5rI8I6WLFRLvUsUcjqAF45de910Soad+VoeRGg7
xbbM6LU8MYYe4nukpHaryeEcyzTX97C9WFg8EoBDCAIgmq3zEzn4tIILW6hkG/ic
0gEXSVfF72+K/b3ER6nY+46SXtf5HMSf0eBYfX3GPz6fLrNHMQnIyE8xQCyZVVHU
FwxA3/hDXkEn6NBge94caEx/a6mbaDzRmQ2Uwzm00nDy6nTxwuYUut+PM8+WiuNV
2S/kPbLcp3r0VNXMqLrOaWpv0pyuTF3lgb3AazpaMCXCFL02nnhssVQ4y/TyyVtA
Rh34RBLffWuxcjUFkXdTp4QTHkFBNMxpkfbT4xutr2SOyl2NZeu8V85d6txtxfDe
uSbQ6s0/zT4KdVxImqcIaU4cjy15ojcAVtII/u49ccuuiRaj0N3oFtHPzdytW67Q
SMQ7hH01Siwd7BF6pCQdBkI1rTPvDpUgmFdb4nV58PP7Dxx/2so6C2iPIvlK7NYi
d2y6KSk9qoJAxgsUtpvqg1FEEmNmaQKtBZss+9t6WipaUSbeMDlnJE4obGQDrich
NE5HhO22fyRsg73I/74g7YOfpvF6PsXFCiZNaf63ushU4tw7X0cSMkx7PAOfDMKB
7L/+mh9fvCUJ0OUNF4ErR/u0YQyof+YvCJ/5x3t6b299d4YVRC3SlpkxBSHoGg88
L0opfQPQTZsJQdsXnpfHJgdkLCGj/a0jLLpHCCxVWrZa7r1jisFoOM06ptiKW18V
mR4/4jv9fFfbTflZUYvOZI+AYiIRWZuYYXpFaW9RZM6kOdbQnuN5UuonbYDh1lEv
iFiA0KXQZaD52ynXoTIB7uMc1qDu5r9eqSudwsdfbCcpZpAOuDdVl5W5XEuQoBPS
emI6DwbRZnjj4yOepTNJyZEOU0xM5IWkoOHSm5LWFzMxa9TdFyE2uZzqer0cj4Vz
1lLclqPhi29jqYnaoHTRNjWEqRMxttAWZmL0l3YPJ/HH5uKtXxrfuHHXWOLwCKCD
JvIpn98D3Hgmr79+zEVMXreIY53J6+8sKMYFpr8L7Jg7cMpmV4OZYsTpzkJ8lt+s
5vjakmmZMqw1S6t+N+4ORvRcfG3ysRwa6wnHrAL4XUcWmrPtaRfdeJxSJi8PoTJU
pEOPGDB6GNqe8OoPKpCFsuBLcAfIrn7IGtd/moIVHBEcuK9XOJLvAbiE7vMhUXOh
iZQbYqOEY+BtDmokWG2YBjW1y6cXouA/Q+AL3KIQ6370v+jJM7x2ELHSzJva53ZS
GjqbEMGFrgDJJxPhIBCtNzmQMM52DSTihDoX2soaFtacMhAym6piFhypN15ywj6R
brC1aujKTqTkN94K7Il+6fZEH3//njKv7smOXrQJBHkUBkS5518AtK5h0279FAam
jnG2oY8n0KGm5azY8FjIghUGM67oqV+eAEHYZ2tuBa1KQmToSJPKDMhY2v3hEzDz
tWN8LxsQtOxqZYgCcleXlOLHHKLhooUWhxi+zTKJaIjolvJqRgR4OoJIpMU86jLH
Qu2DPeN2BYDRVM2USO79H33xYA1Mo/yOVDVacBQ+AyUNLCmuWAe2JbFbeuUzqgox
wDJf7PxIYztXE2uc4+WhFu5Aiy+qcXiqBOuMQSHpQxErCUJpMaFfkepgE7/wP14J
xmWRGaTiI7lQJqa8VUptONK3un4Z0ddQ8JJeW1rHo+uneW0dFkaOUJWaWrp3a39M
Pb/OvrYvY6sPJ3UyY2lXdVxwqjqFJgG8hjrpZXQAdve1Ik5K3gXYU8gcTsR5SFfS
uTedDtWB/sDqz60/4rRmsaxO58bAYb/aRFPII/pRUOBOrw3izlKjIK0Vz1cWYJS8
cxK/t8WoUZ9wiqfPJDnzYYMvuUevr09HC+Djg70a/fMPOC1rTCUjF5hqQWgMN4ci
aEJohEP9UnzIKEHaqaDx8RFZ/UocFnsVP4OzppzJug/7/zgTsAdtNpkvQYE+x8ck
MY3sMeguTx+n4jvgzkD0slJzxbRJr/AKOGJfACyzpFtnBzBr64g764+Htr/VEbuf
B3q1twwuqgno0S0EzSdrxckWwvAvu/aGpnIjM+69aF8fx+vrEtIdAQEsIq+mJwcg
ZWu4bjKpGr5ZTGt+MNuWH6hqFTMj+6mn3e5VBRPqEkJCPJFLyA293e+HV/ZksIGt
C+hv0t96brw/+SfnpcT2e2qF+AUQlu2xdpg66MgviV4VE6XLV2+ahclP5iTQC1Gw
6TQhELJP+QsASQMnqKOuVF4H8Oi0yMsCA0+zO/1ZnJAGXMoo1WV2G2iylm6aX7O5
ubeLPWGQQ3l4oJ5Jl1TJm1jba9Wa+4k7UUUg/hIGk70oQ3i41uGWsGgD16rrAkc0
a9OB6hpmPOCI9MiahRbj6UZnwmORYgc5qDLr4Mk9RVOlvrL+SRW9wXrV/McQcgAW
h3vLL0itaIiRO0rU1QU0NrQonQ3BvOplEdK+PilGLJjMzjTRIhtEISY/nZfJCV4x
9S99XTr8EnOZwE3B8SCkNudoojFAgkYAvEvDWDMuq5DcFXU7opBCcIR6YAZHo68R
ZuX0qpms32Fc9pcsIN1mYXqW+mExVHm2X7tuYDvtNmKps5CPPNax42tDQHUx6cq7
A5n0+EKfVLn0dvn7NJeHTeUXhUwEzJHU1gjc8s08ziiiCdbYdqLRg4Hh5ql6AriO
itS3P/EXcPAs5qDLEDLPV8SfRb/oyTx7WNDt+d0WRLVXZmKdxooD9SgyxHKfGMZC
PwiWSob6IoZiE3b8p2IcYZzeDoYk4HzcbilaDfiSpNZH+HEw8S1wb2jYHS2r5n1l
Q+9mReynI6EIyrb+pa7awUgvLfUIM+ht8Zt3uS1Skf/HbtjfJu9Kvrz6xUS9GLYe
0iRtcFb5fAvrSBAyU4iHs9jUMSZ9bPQMl4dtyZTuNkY8vrZbUg5C2tJIyn9i46eu
8M/WJguidXLNPSKnlO3nRQNMkWM1lfdB52KyqBoKt/lSXA+ddtCJwUpXoIgO1QIO
QjdZXuUm+NnSwRO+Pyy6Om2HKBD7Gzt69jwnOJSCpof7Y+Ol2DCSW/xPJ/a8JO9x
5ihQUsM3fR3dUEOhKjEGeIxRBk0GJHCvwyf9da99CObRV5CsBEH/3YOZjo7I96UQ
ygj7oOtOKRhLtWM6Z5YL/uZKB/pHK1nY/teNHpwG94zRMWsbatl0stm3f3peeEge
oQnTdIBtSUJpFjd1AblNu8wlt6w+MozlysYXD3UBvGsnYf/9atU9F0izlymlfnIG
XbTAuJK3HmxCYx6SxFg+w0U/Cu0rjvkIelqlR0SUPf7s+kSILVHzYzjn1bZ7k7Gi
1S7+OME7OQ4M0KZJFTOauHjLaz54UxzcVMErxHiVs03fKxRlijgf5WdV/qbJ5SGQ
YDiDn5/GT5LdNCExAU5Wlf9TPv28Ga6GVj9MQ2LcH+V8ezxmPR079Lkk6MIvA5B6
SRfBYy6UFvI1z8bbp16qaN6qc9dAid1DEP2Cfz5oV2tckX/VOzmfw0QhRRHidXKM
+nL8CGc3RcMnflgvR2VI0kKqchgLLLK0wTPwLuKUuy/c6Z12btwhpgLD8St6984f
9Ypx1SHE6zcMowzW/5p4GPFp+PuyyOfFl0ncTR2oPKRARQFc8yRvQvYtWmz1kK7U
KtWRWEo+L9VGoDB8AwqKTe5v5taxLl03Jpt0zgfq2Ge5g4x1pE7s5m3IGYqqve5N
ZSCRykzM93eBxqv1+oFd45ebeQSYV5UxWBvmWVkFUjSmiVWTXoMLE1so7jcrV6kB
tf6Syc2LHzpa18U+FS+AL35D66b8D2u4IrSu+Fr9ppz2KL2o7uZNfVj0q/2qTB3Y
7WLuLj3VPU1Z6pq+1DIEocOGCVIjIc/VkAgbLpWZZBlBV2emxUbnLO3x6GphYLgc
hFZAY0akfP8Uorx2+a4hxeo9EzVF+IlgpFOw9e0WS9+GKydUBm98zhpKn2+J1Z91
aQr5uZ1l2pNx9RKnwoeardPFNIQyB4xTTxIox73p/KRI6oYOqEppfK7XRI1D73f3
yaFS38ui8siJa6IuD5OhxgcEuxKXpwEhoIIemHHePvbKlXmn4C00np4s/YSLnedC
R3fHgGHWjygiaOuB6n2tS/YVLNzqSCApJVLlSh3ircXEJXlYwnYhmOeczo0X+k2b
oqu0uFgf/CwbK+D9DRVCB/lvverr7lOh9+r+DZ+QBkSdm9ztwuFL2qwKNiMtZPNE
DZIsncd4Ep1aQUUn+tZcrixvjFZC5e9NOo30BnVs4eD+7SOfqcQcTLL4TQKubyaa
OiPbX9kWyhUPtyP+xSe6djDtaVJnm1PBjPkDkhYRPlDLd/SOR+himDhIm6iD8xaM
Xlo8ncygemMHw0N+p1J4qpqeGx0nRsCwTTnVBBWapu4B0BWT5/jn3LUzj9bnYbMz
3V7ls0T72/WU0ucIh9WvIQK+GNpTBMCQCNKbMM9qrxoAXG3lSqDHFZGJG6+RiB8n
kSckgVwCItePwA/yWlCHLJx1vcyuEAV5n2l0K908xH2iIdohrDnJJVmuMsxNI9+H
s+TrjfeZlQH7qbahBDWuS4q+0FAP+XRyYUlnG/aFs8714QwRUruX9d3DXAaeVxwu
H+AoSG8PdHn8SHh1UKGcaCVuDmRajqGQz7eSFRLNkt+AeWEmkx1J5DaGggfJwq6d
unOk0/IxndRCGwW/0uCjO3kk2K3/E9pIHy+U7p5m8escHVTF6/nUjymqiNC0ZY4W
wfRj+cziEukOTEMcRr5EvPO4cCl0kN9veX2rh39xjRD5svANYcHIHsgbNJjhQgSC
fXnzfL7pOoaOv7RUiZgY2DO/PnkmkTY9q5VxxfCmpgBvbRxCCQvv9FcXDeP26RKL
TZaxojRx+mgPJajIkXLUe1TKGu0y0Syku564AZASX2710DCp+NilXPUGO9gn7b+A
pyPWpbzwH4MNePXqBB0dVILXmcetDgiEUcz47oX7r8uAKLmE/289Cej8mgSsO2H9
zEJwBqNQXmNZbYd79rb7fiZ2QPl6t40iDwzJ7SOWQmu07KhHzrHYHd0yM2+J9UF+
awYzm1c+a11w4yQWQrF/FY/D24ACcTONYxUivkJMFBPKEgugFVzeziEh4ISdDLmp
HV12okXHDfq0AQw48MgcFs6Ww9ZRTgXqBOEQXAEf+3b8qbguXTt/JICl1Vo4TOUs
B8wYwszItsRVMNW8sMrUETdmHI666x/r9Djg0dlp322wTVg6ddmfKSZf1PBf+Ofe
0Xfc+jJ50z89Je45GGjf36f7aRovpoarmI/7XsgS+xnTilJ+C0Lch4AWl2uQRuaA
WzrKgd+k2Qz2MKU7FZtSLvHxKxtJ12NkmKSbmUYRT9zJXxzm8rYob7BFE6yObe5v
BTiY8gqNcTW7NS7QLuMUxnEsYP8/EhD7M5aZHAqewdKHbJWxnj9M46TzDZvlqZc2
HOjAdiuD5uzl5Pe3pmn8mc0s8ZOyrQaDSnIIc8Cnh96nJowEl9RHCJeT3+J8J2GS
1LD/ht1wmdXvG+VulAhe5L29X4EvgSvyNO95sBdxRxickhw3KU/8CMxkExB4vEkh
SSPl6MWDcQdqD0ifF+L1gW10o1EMdyANyrW2pKdiQxJWp7mHUiDJU+JReUVaRuHY
LRafoDo5G9e6pNJWsYfljehppBx8hMUd2DJlIbX86ETjSsucqMh7H+mm5s6h+E5L
DQsbl8NT90XJlrjluDs6JJGN8Zlqtc3w3pGEGn7Q8+rtRCZ3UZl0rItNlPfIakKO
305BymCnHRAQiIOrALySyjSmVPELBkYjWEb+xVk36LawISqXLGDtz1JZunMeRC2O
Rkrpo6NloOuIqiM9IPRztC8eltZEM8Cgwxwhy6NcXiDnjHbWmgKppZu7UhUMH2Zj
Hv679ypbVgHCFM36//xqIspo/1OPMZZZydkwgnYd9bhjkKdbL69mwDluD2fYguUA
tCGOsrqnbLo6LqWxDq/9oAbG9mlVALBcm4FSB9vwjQKc5JjNt80gI/Vm1n/LNu/Z
VGy8QP3SWmj0ztFLxeWst6n+eZhuna9knezT+vGxo6vXDAttLcr//H+Zx4Mu6b9d
SBHae73D2b0awiV0QzBqNBOni+yav9+HKkEUMovZy6zUZw4/FxVTlDY7O+lmWQs0
OzIJrbIZ6A+aEQmhvGfp65aR+MPMxkPK+44zGnGJF9r1jA+eXbrI+teu6MpGgaPr
JhDmfloedWIReOdokDvTW+9BAZcG9JBNoMNh21h8NAudUqu4W9DOfdSix/WFqkzG
EBvKD2KOERb6G0+Ptg2jRP9pFZVnYukG11FhVd3oeoghinP71QptaEvNX2nX5XB0
sxHYkO45YOwSvLrhUGokph6eCGZJsSTiDCr5bhVs5KgC1H8qZls8mJnc2DLnNleg
Q8kMTekbKvFldgVkGYpdayksmfo7DBd59VNwMNb26uazs/fO50+P5L5HKAi7UCzT
Dhbe3t7Xh27d0BLzWVHtIcykuFRP/SpjM638Z3TOkGbaiQwsUUjB/YRSMENv43Me
7DkUbN/KAWT+O0IJF7EN4oDLpOo7cPNcPhppe+9DiruR1an/nWAWNEBDZuMrOsWz
ufsvbflju+CMmh3E0LDEjDGU9nVI4rDmOBNnehHFuwkxqE5XkTV4phSqg+W9wSO+
rstP/W3VlTtvG1vp7qC5uxR7kq3T8ZSm2B6Xp/555FUrrQd5dEqdBlg6gqczE7og
qI2g6mIGdannv9QhA7Sa3RgLcWsabuGRqJp1Wijb4pVs9Qnyu23/00Jeh2jbYIFF
xeRUcE7w/3d+W1ezBgFbScVkPuVATEmoDnSJow6AmUJC8Fx0L5cowrvTbR82RUHN
YSQ2Vwyafn1Pk8kGgq767GqYm+MTWRIx7MKRsAIvqP8i/NaaB/kbIOyhEx9CeTeG
ftAk2+SeXbg35ZuV3D2iyt2d5bg1343IbQRKeMLjlfwjGB9Wo0J3b0ivR2OKJZiY
7OywLxIziCRg0+lZmeAX34Yjo27mbs0UK0G8PrYZ58u1NhMGBl87qHBo0ZM/wVFx
tgAItzmRw3dWvqFjkEuWnU2mjetq0YxmrVIqdnpyb7JlhD1Kf4gVj8TUVP+gy2ph
XFSF9JvaARzRbdyYOB6U0QxYbcto7CJQI6c93Hj7dj1GMoZVOE3+cAn8cHUiDao+
XPWrubJGQEutJZMMi/H4GREot+hNhystdx0E14uL48NUAqiUoCCgRiPcC/lS+op7
+GGLJ8m7oOhnWRCOGvXvLx1uHDMOakkiOlTtgsOOUJzK72FzF4H1Lq0pvPkZDqiM
by3tg1UFJIuTuc04eTD69k9DYiA/wcMMVdJTkKxXdtTV138aXxc1QGd2WRdtbVyE
YCM9UvOrppYDcsdn2emWrZ2KW4tFgnq0sT+4y7+3mYHLUVdLKKP2pF+fi07o2kHE
UF96Xbe7HDuTD/gvLFKYNfZiZL5TfA+pe15Sq6kHUdGK2j8ukUAs0QJGHQ5VIej/
H5Abv4PLotp26aQiUZ7Xt5L7lUwK929zOPqFTPxCNnCg/I3fhM8usZUvz9ch6oZb
GR9k3lTECTerX9GyRVibKyYIJdTWpFp+7kqFNFdQfalAnoP2FNnBMJY49FDFSb7X
IlTR++6Vj2LtMFbzslYE0pX1R91tau0Khn7JYEUlMqjS8uOX/0uGLY97ou+2orIo
+sBvrhUk7dMhWF37TufP+QncxuYH4lSe0NIV8S2MltdH6CQEG3rX1zNfmtJmlWPt
RV8Je612fPpsl+yBL1+RIB4KHqUQbM0uCrHQoS2tggzlHolV3of+v2saJMcGKV84
XPnaoXJuRPAhc2ivHiCs2PUJz0FhbdDmaWJwHwgTQNQTlHB418NV7fzP0H+hvIk2
H/10rVhYfiuSDAiz9hLMYRLKeTyWpQQDHNS2nhqHSiWcPdrKnBo6nbhx2UDO+qhQ
KhAMWj9QF0rqSBcI6ecNZLEjk8yH4ZbtnPJtI4nvihExrbQYJuT5vrnfwC/LBzm3
rnnhtE40+znFh+8b82HCfWql1NZeA76WkZtbLvo/C4aApkUmjWp+Y7MqkUgHszkl
DGSv1jqtkwBVEYFKxw4PR+6URRUrqlc2YsPurrpekkZA7S0mMHUUxkz1jvir5CmZ
JeDCWkv4bGmnDpjDpQWIiZhd6lCaQoB24Iz5i2p56+hr3HyRovkMiMGFMJ5q+3pj
CtiK2px1rNZvispumUjIlHD6FBn4tXtENS3E41w95I86K0fyozmwlSbqeW0PhuMy
ZOJJkwGoE0J31P35B6/nwGWMcZdJRNYuAE7uNqu5VXK36MsuXGbxTcrRmkT/IQpm
g1etKv8Jx5xCSCgATaKPx9WL9nvdjVnTnSYRDfEXZwfIvA7CG7TMwd+D9Ih1jjkC
RR3JuKb//W5QG80eCWV4UEWyddZhhRGwN17hjLIPwZF1c6KlWQLFY1qTDTZbsbC7
mhCFU6478jqYcJA7e2CrBQ5s4bKle3rB3d6/Gfpe93+JZ5BO89eHRyXUcetLeiB+
buScqvwPfS2+PEuYVlyXpD5XSHv6URS7dsAxJLJL/bgfsTTTaMxPWQZ1JTc7kzC0
lQqF37Cs5c+EmQl65wA537jQw4YItOuswRaVqBUVtOL1CTQGT9RL6a62h91U9rjF
T9kTO0j0b69DXpLZ8ag9wYGuN4yKI64I8agmSUGoLXoLrsO5oEoIrUFhaf5nP/Ao
/w2jNSzhyRaOpcP7bl53BOI2zpcNz3wFRuSWh8doZy+fDCymR+bef9jOVUksLzXB
mF6VTIdz6lZWTlkMppBFC9s6fP4m0ylxY0ivyfAX+nG88tDXc4qSGf/7ECdVQGrU
mCH7Pr6gDKgv/Q6C+qEqkk3zCuKPTjWJr2BVHQAu2MBcYBJN6daEeUzXZepXZ88e
+0iGf29EC2QjRxTgWNzu+JZh/EtbPIJq7zc1rOYYKLftMxGbX6vVxVWSA07ROxEI
xt/mYdtDdXznMdxRv6vWFif7yifid8rneRDVRChQClWfzLRZwiyyfxdoIF/0XehP
De7NWZ6QRxaOxZMXALziPlKYLjH+HG9SvCrNUSDcvbo8UWJ4+3ereGprSB/XVZIQ
dL1Oi02ThHR9sdthhH3wOJGbHpFEikxuLvoGPFZnmFKjITC9mxafa5G7c5r5SFJP
AeHzgK/bzPxLcD/ExUSyjv+jmfOKIXqabWc68CLZ/ygrhWfzzrrrmx8uawe5z1Cz
LE9dV1CFacPw3TROVbT99h7M0+3SwKlKEEk2fLprJUjJX2dcWvR2Pw9ZC8jP6u8J
6Y4YKOrsXpnV8lKhuxVyBPJbBa3I8FWUe8xtIfNkc3s/shLVhnN7XN+4z53KPbih
7K98urJ04IDer1Ne1tik6uRwxiYXpTOQx2UQtSuzP1GgvxmMBnbVYbI6+JdJpiaM
x8s85AgRyKAPAjHnUZv63dCcmjegFtdt+mVH7klI3Bv51u+2UOydgE/fbsQvwsNM
oqL7f4sJiv6p/SpxWXcqczKRcYjgUs59s23Xl0LEJ8gfycwYEGQ071yKaw+cP1E/
KXSyNTyFwfEaJN5S1zldMIS0PHunMBgCxEJfaPXBx6v6ZW9d+QRDspMKMMXlRZse
z1CASAnJDj+UO90vHxoXA9R2oC5THh0zzrYURemK+wWn76tjlX0iv94DyMiDltMi
IQ9bhEGrDMikzJpXAicfg5BvGlvFzQduGXG7hUQueAHKDzXVeodrmYrGzJJhbDNn
4de1XFx6InxouITR29JUzPPKFI/XDx46aB5WChft4EgZCnDPSwy6BI044+upitdu
nu9X6a+APQhy882umpTt4DtXDjBZ2FNfuodJOTVj6X4w6LpuIh6PUWICHMLWHbID
rrUw2xCtmnId/lx9ZQ6ShVHV1h/20lMIlXjPiZo1Wtby843+l9iNYzTy/y5BigqX
wSaUx3Hp6MiCOo0Z7KFGc7hZ+kdvAiyaz6BOm2xCzC301o3S4J5q1XSuR+bLhfro
ZwmxAEMYin5m9bxTW8wpIUTjdMr/jZPvc3Aa2id2pir19d6fc0eiexgydpJq/uJm
xx7LGmRkSy+p0G4R5fNX8JY+uFK2GVihoTAKl1zPFR1lJ1Ud6HAt5c8olMGnmRNI
Vh3jprX+Km4Do85WkjzsZZDN7I+8sc3Cj+Ary9HZRzyQoYv492e7zD0me/R2fX97
gMA3///Jejq1kWSA2b2eps0unT5G8PHUOvVae/l8YgN5o3mFfjrdyeXSoA7T6ePL
6tAYtAREtTwJUdHz+tKafiR4b2r3hXwMkZz9fWEWyBftuPCUeyToGsMOMRGXpgmS
ux2EBVBP3yeSGudHjnBXgHd/TKdptL2rdO2VzKE6Tpg+zDz2+c38WLyPSMjxzqpw
R7tNM2Z0TapABNXOFsX8traHtGzkFcz0V40ns5J4sG33Wfu1I4mlXKwQ/gn625NI
THXcOC2CWnOq6aJp9uXcsetdt/erCgFY2W0qELjAwcZtD05qLjwbxHMe7TFqfX64
bFMwRupjbNFNgBrlDUoXDVI9V66gOoF0DxCYkBpq623FNkaRX9iTY4NVctlXOb9F
XSrf2iHdR2dyyr+Le1ZLPa613UqJgdIKobNx0NvALalFEoWnM9bejEA+5pBGHOpA
OxIIqKisqw8u0+rnD4tYzJliV3YZ62fckIIEukgJmzdQfdtxblsvJeZkKlXFjREz
ZVWQePMrN/Ww1jnchinNtKgbadcy7uY31Eu4uO9fDI9SUNBWyfS/VqYuxAXFcEHU
hUubWBtyENloDS7DnVahegMQaA/A/tq67kjk0lZM1SCX3syImDdfWG2nspMPK8db
2guB2LCbv9U2lbCZRaHmzOCV7ZTKfnNMohJp3nxhAhs1bqq1u91qvepNIn/gozR2
1KUL2gmgnn6yKsbVrX1EW4TxicFg3EVNsPON7jjK9ROxp2bo48aSTbOQehmUMYNo
064OprYiH0483AewB0I7FYGomSWUuUDFEdT24PQU3aoZRFge8ipRhv7mmTSawG2m
liNoDGMvBeWelMymXV5Nk4GwPDj8mljjD4ioc8I8yPBgV4iJhOX7ESmLFIwgACOQ
OuLSJIPt5FvgkqzcB0/u9KIS1+9emn/fsZ8QEx8LNShn8w1qgg51twgkpMcLeG3I
bs9TYWUxqBDK4V7BZC+V0ipqYlW+ZRsIbZG914k6R4VpRPHsAtPFhCKsLFUMPNpF
YalV5Y7v2nJRUFkWad8TiAjLot/HOHR68LPKsKLes4uJwbSQSWCCNQXfJUumA/Ts
kPj4bYqAOXka62Mad5hyLNsoxYWFsVUvI3Isul5M7bTJOOH7L6TmUVo59p+NRe1D
Efvm8GSgkBKR2ZFD4rMVW0kBbJD1Ojf/g0Zag1cIPqCdbO1Os26/Qe3tYH0ksMdi
wpXQmwH5ZxiwM/S+NnN8s+etFSTKTwZCO1MXvyQooH5GSxacjGe8ZsLFkXsADeSn
l4CIIy9BTL+vAYNNmFUGK9f3UZfky6oPWDrvqB+FYFnA/JQMckM9mV3MUs4qkguO
8yIpn//UQIN7wz08l3vPnafUmY+SYDzsLI6uXd/hTwsZUZhH7UASybd1ji3I2/cJ
bmmgBLgB+yErP/vumnMJPeKdRH/HYejEnROXtESB8y/7ANsGlSlLqprtQPliuuIH
g3IyMVxrCnN37xNBXjHaOiVw5DdRKNDp6LX7pCLaHFWATue4DQcrehao6i9UiJGc
GkDMMxLhr4/pSt+DLg+yNOt0GFXV5crMWLslNFJrsAJRlcXZpPYzpjRZXTN+QL/L
6WtE/BA4lkUKTPSlPSj0rFNrkPsHNLI2h+Ptj77YrRHD60MZbGLfyimWMDgGN+gg
HPxoqxGcBxX20VLrOQgAu2X9WnctFdKoMPFfyJ1S+BKh+0+xW2W1AE8Hh9ntBWY0
Rkhdn0HT7DFcxULcvnpks87t0fr/sWJKWNdlWRHVnkA2q9tvzd4d2qSWWh7hd++Z
atLrBy43i0lO05Xo3SXGHSHOQO6iEQQTIIE2kKRSg/uRMgh+QJZPEPJrZk/KlqFw
6QtEQjV2/baxYSRJpSZwmpGJzHB/fpgVKZDU32Y5hp5vd5Fr05rv3pRv9/weqoq8
7ox+YuaVN2F9Tv4yE1Cag1m0OVwWhgVrmU/0WZP5EquahsBQQSju1AsreeH9vITX
11E0M4834JZ5vvC0fNsDqvHInt4chORseKF6a/DI4KS/laFULhhlfWHPdD+tZYGI
MsUm0jNiB9rq6JfEjhGXTzzFNPC7J+8IPCfZfJo8deDup2Mk/Oxm0CLsqCSBA+Ad
phGipspKDZ8MX/hFFvQ3AtogR2w22HKBhve6BgrHW4m5tL5lfhLDPFQbhpZtaC2z
D9WQXvrpUUtdeuVWMLxOkQNJXuv+VzGPIZPxdzF1Zhn9apLK2m0468Ck/lsEH9Qi
z8kVyMAJdopR+Y5PPqAYZhwEH+6QOtvLeAuyCjNC5La5xb9J29OjE+B3UcEZPHLK
R7Uvmhf/imrcL6sUgcRJwZ6Fi3CSPJAxrnNzr1cWpPqKxYUaa4BVL+BaeO0tPeUI
Z/umJqiCsTG8Mt/BovIt2F07QrwACfJ9vhRy4ttGaDJYJK0GFkM3wYDTGc7Hiuqb
EI2Gx9RMZNsw95Dqs0iF3dod+UUvOmDjgePsizUYkJgi0Md2chliOIp47vMm0Ru2
djkq4T6IkLQU+tlhMsbAJx6y1eFsfVdtpJNx+4rUFVW7G4LxKxxjmSXxkpsKsO8h
NeEGwWkQQIsVxhxj9sYukA/630od8Olh97GkSJryYHngYamr0Z0okx7PiMbDHsYO
dKGzOV0XfhLLatFEw/4XnJqoCb2nnGku74cwCO4NQmgRW0ZtSxTMkXi3fn1+L8Lu
+YsXX68rOc2lKHiVRzes/rLubc2y8KU3dlIky14b315GmuUjyzwhKhYAsDaiMR5m
Te3YHw7xq68DFio9NcxQH6BBDZWzMK098ZyekENxmlMqoAvrborTRpK9RWog2Vue
5ifWYTVc0H/4HvmjEqwwP0f7dGpw6uMnpojK8vLDthjs9t/Mv/LdWQH77YjqKAE6
S93p75GiLwaLLatz7VITvq9YSe3SoCuRY22UzEPV+ccOKjI2Q6opXdMZ9qXqic6e
wmmY+m9iFk+WQ4GobKgFiw3K1TJfR4j7lO0hhNnrnRixwR7x2riFxGyaYbhYZ+3r
mwmZZiHbVvPbmiCjthRzw3Aom/ZwL80E387XDaj76FmdkpqiC+qOn76UCaYbNE7L
RKvfnn7fKZ/aTnEUDKdR/N6lMQGef8dhLmaNAqVvOJ+dEuFA38x7DaGcRPfaKWXh
ZYhFyCy5Pn0JFeGu5qodnm/UVrY6wDU86hGmfXxn53X/ShfkrhI3eFoo/BU0yoEq
n5Ikm3yJXtxF0YXKOwmBqtf4uEh/aoW78N8Q+ryE04XvbNFDPh3+tkK6NX2gUsci
96oqOG8L4TBI2NX9jdSrlvtVlev8lLgRoOvozKS8zFGXkU22BLEAoc1PdEoD2EWL
yQUw20/94Rv8ga7027Ou3C/0chRwu8llT4U/TZ4j3tm13O4+xhODvLecNaFarUPR
CMOEXKi3vKv+iUAjErnzw/EDHn5rcHGlLDgXetk/iEJWYmBRc5bhD1b6+nrC477o
OyPQTubuvLnNwPXBaec2xOBvVytZg9UDhj8mHb1iyr7bjPK8j/DLjDNvUwTFWENp
aaTIn84/RT9Wb1pOsP80P13I5dA8sVVOWLO53IFqJheeLfR2LChBMpsAcrTHW7Ox
dSvLsqlsF8IfHFPFUFrGiaKxB1cAqyy7Up1jJm1cMiUGXLhcy0TerDOShPPs8O3S
wpSxHvRctvSzZ2l90cAJpNsbmWr1WdXBYjyzQR+zp3456gkulIvMZSfGH0EVX68g
B8RCcWQZmVRtpdQuHUFmlXZ/HEqrtTl60Yjlxai3amX6H/gv06JfPXEFOZWCnlgS
Dp/VjLpV8oCkowzGdWJaqz1wTuoAQTZ1mzrl7DDsWtjA87ZMKcYe0bdcHPdIyTVp
U0zmQpG0M2h8YLT1wwmj5cHcOY4bbjBqbArlkBNgIkO5tgVbKIANWRgZu6P0+Sw9
NT1EF1nl9DxfB0C3Gr/YTf9BHy58f572BqubMzbpAZDAzX+3vuyUl+yQ3rTIsiUw
4CP1HjODOqLWH6EQ6s/MaxpJN4I39D4jbQdQiYIJc6XUqHGUsmAVFYDuBdaEWFb7
+lY2L2TDo5lTdZhajYyiKmi0xjvoVxSRInF5DZk6gHLziNSHHJ0fWj0GF7ic/s/D
O1KuXeLS9brj71k1Sbk0B2qOYfDHXJyhynmgiO/i3EopHh9As60bvV7mEzNZH60i
h7zaUorxpgdWhEzBAElW1r6WGFnwtraGRDW0M/F8Tl8dQxFsSjuHNQ6eNqml5CgW
fd6qAJug+39E62bV3ZmZ1GUiNAWOl/mXnTy4QeJ03sDEtATV2An4I9CyHBje8gaA
Fg0jw0J8CLoI+Lii4iOxjxJBDo53vhXhbYcgRbEjNc1toolR6mOsCgvOWANjoWW8
I12tAZvKKE7s18xtG0pDRTBgi7XSGdRmHGYX2FmoXp9SfMuQ1ItlvUS5FjAjgG1R
GbC/15ooeQ5pJE+H0dj6xz7cIdXvHghZ8ZcTqvl22tWEQYL7x/oq4RFmyzf07UF5
37Ka/fQnOpdKJO9Uhd6H0ICzdDGnD6g8wKGuUTAl9GaLTSfvz9wDZVb0kFxUwauK
duy7Meu4dP8jy+PSmQtSY0K1TyR+yTvBgiusnP4ouOaBsiU+TVcfWVCEvLKDBKko
G8i9AKu/iBZSq0Cd4+ISoDOCXYWzCBhqCQF5+ARDdS9Pmg9b+xi3J9Qf63NG4x4y
9bcyqk7tS1vx8MIYvCxCxT1wWWRXUMXRMGjV9w+d00SViFLYtVpdenZzKe1lxOSB
jY0ZpBs41mlsupth1QBbRAN32OPV7ZDVjNNTqVz9K4W5TjN22mKrYS3AyoBVKq1Y
bBT6hTZQWvDkbvBgteIK8JD06hKI/TI5CxW/a4MG8u0VP0lIjQIWqj97sqsKmcxP
753za6W1PEX+abcebhdWXiD8Zc5mbPUBpy2mk1immjwtAFdGxD8pSwAQ9SKGW1jc
QrSpwbw/W/y+QyQROWT9U0pGqZNtlKJnmk+XhEHCtbUubO2p3P4tN95n4XUnFbF3
dpd5jvdwZnml1c/1FEYr2PbeeGHZs6OIwXcTBFLKvtUDbtH93p2QjGKh4M7umoix
XziS8gYqCeMrQ6llV+ECYDqaT4lEVKmKYPuGLg+PvFm9PzCXYUhyOmahZNCQjy2M
7YM0oW4wdOz4MBdAHac42xqGI4Mlz5nkj6MD+XY7CeD7Ms+Gw2haW5H6qiqVfrOB
RRliw/SAi9g1ipx082zVEvqqFkDUpfcgdVn99WLvahB+FduETUTyr3+SX35EpHYL
tA59Gu+fi1SnavMmmvGyEdj4kiMAy6RGPxxvrqR6l7eWlkBQp5zLIGTdEesCWq5h
24o7KpQwVuZJ/SfD6vy2M+r0PmpjX6kf2JlyC2xfFxmbp03gP5ZWBdPn1hEp4GH/
kHjlLLLXviYwhQT6//rRYlTz7TB9ry+voe0TVo079TdLzskH19fkwfrGoZpkWbdt
nw1SMD++2ukrQ0i/Jd6F0SWZbYvoKEAfFZMKtcfTO/IxPb+iFT0G08c/Rjb8cxiy
sK13AGs88BDTJG5zBKrPryd+96eTsiSLNNQTbPqSF1dlQ0xrpSUl5TL+qQ6UQJwO
EjCQqi3Tp/PW6Xk1j+qoJRKjwW+kQT+MmKEEmkxZ2F20xr62ytnRE5YVS9+3A5P1
d4Ryl6FBCBlt+wtbNVoCFNtYQikb71AR+4PTnxp1baqNN3iNwKWPVM+RmYraDfaX
SxpX3hwuHZ6AcOiQUl6kPuYogoJEKfO12+Cj6Cv4LFLoE2DowI+zWVWcroN/taeq
aGeFIQfXD8KTV35fmIhDRd3/vX5lCQMddB92KzCDdpVURUjA04VzqUn99pjeZp4l
vUaSLLgJ4e4jXDpxMU5r1xccHf3jo3eI0kg6XNDCEcf1IR0CyzjblnN8pPWcRn5r
OTpV8kRJmnNb0yoifUwUz1l8TuXDoXQztQ3NVVLrux+FB+FcBBjEf1RhjbJJ8SrN
LqzOVrU7WSiIFgfYyPvqdUg3D+HccJrrVwem4o0mVqDyhxjalkSrdA1+tK9lhIoo
2yWxDXtvHw/TAY/B4TCrkHNBVBhCmGV3Yp+wzVfEpt6OIyNZTQxBasgoFgzBHANa
qGSostaAB7lVH2sG1pJ/CMcnaKp83VgSzwGjvJJaJUtnfrMDNFO3kMJtR14cK3v/
hfJ/TI80ageCtUkRtbDR3Fv0ZSOmnmbX5G5oW3A6KYvAQ7fXXopALuq7f0NnXXi7
78xXaUgKaR692G9zJ4a7gCoy1qM9paGhy63TX2yXglL1BpH2xLKw93ZJfCUmL2Ci
y+Lt79UHiY6y5HNQXdKwHb7r64JY8V6EAN8cu0z+RahbR+xxaMSVbE+CHJr2kIQK
Q3GR8M2DDYay/GhRkzBuH2DlDOv2uAe5umyZ7OpJMehYoupINWR9MGl/+VpEJHmA
MgXxFxJagoU0XXVR51Me4Ug3OfHveSvR0hW2dqnfz9FppRoNb8FRxIueSM7BYKtv
KWqZJMP6G4RP6mH4jrnIublyWb3/u6GV127E4QSdb3Ou9kX5XG7lpbHvcztnxlGv
QsxRpH4VQuZPw+FLOjLLg7u8fICxY9WNg1nil7WtFf35jEgKehjX9rH6MXuqA1AQ
spXRjnwrg94AgtuKJjd2zhlQ19V83+aLIzoy/TY/ZAbE7nrl7UT7nkuMpDdPYHDm
a0YQQEalF6r4u+2gMtLfMuodlgDK3Rrd5bRSXmkVDH7yZYoe35UcgMonCJQEBlnK
bYecTmHB0bClfElH2/JRwdFReDNFVUCA9NspW6QZD/vmI1foyM+8AybdONktQQve
jVvhSANcHAudtPJSplXlnYjy4NLRRcVk9S6M3M5wgRJ8WzkpuNSKdtxbtUOzPDh4
pRmw+T9kRG/aojyWV4P01gkZA8qZYk8qY+hLvctcooxe4JU2wDuy7yXqc7Ncqe9G
ZygLDwrIdv1IogcVX/lduD6BHSsQLvP6zHF7jVTuG+RBGbFL9Bqud5CN/OZoxwSk
6qTTV23IHa+8/Q2xracJN4bPFht3lKLMeYh1xNm62j1gROz6uPKcrMv9Dn77MOqg
bYtMtuUzbUyXsBiggCdzeGLjjn2uTZ1KM7Slt685Q1DFLPPvcjkr4fTdRpuMgTvH
ci+kFd9VZdIVKg1IAhEV1bX8D16T1WOMfsxNpNo+8+QBRqHiUNYpakHKoENmFQqP
IViW4knt+gIj4uTCedsOxYotr35xHscWrYtdsTOOkgUoDDEo0k8wcMMUpZ+dy3h7
0a7r79+SEIRDyae5UFOt1PQGy6nwIPhKMdJluCGlRh+ZuJf6z2JMuNQAxRUCQ3po
b8+qBUOfZnXWZjo+vZ5dMa3dy8UVyEMiRyyAZJFPxuq5yI6/uNiVsDrJFarPAwsW
hJO9qQkOkHVvNklhab1WHtB5pe81KSU8Sm8A2RB0TJ7Suihhgh/d6PmcOBJycIY7
R/V40Cy52Dl1ingIYpepsQzNW8hZDsDLPdsmRneFhLKmxAeQhpGx/qw5Kzhksgew
II9ScxmY5mkbgGjDbrRfn+qhH+s/UQF7I+KvTH6N7vTPuN3kxI4pQlZi0fVPoakv
F7lNJbdhe6IZTzHDy8ue2KGlSJsYN1TqMPmHD43vW6f/sL62hNWBXILKs0CmRtXI
jnu+3v9lGv1z1Po7j+NQ5Y4NVV0fOmjwHpEYX5Pvf4ORO98/EtUJZqlBJhqxtXCU
VspD9E0HSMYQcI9RMnCvIUtrleAGqFQ7cPv5icJsM3E2VYaxROjlfFpYVfLCbz1w
60IZ+tBfjeqjEzLNBIJLohP1NLThkQ60U6HbA72nz1NTjalxElPKVrGfTnKWp1ai
JQu3NbiGBX6E2DM2sKkYxw1Eu12YnnLZnB+Ne87H8EgshNDFturVD/ASQPw0OGS0
mJljjitA4KjtwHUvIjQ0w0kNqCMEf0EJtU/aH161FjGBpqOGIYjb6b8j4VN4QII/
XFFze4YGjCAyVGarpl/gQdl37c4YF7tX3cRBhnSdaLBwARHkUbttBPaAaLHT+WS/
t5aEKsFVyFNzjH1Ow0fheus7mzZ8fkDjX/FWBE/lGtRlOcRQSwMfK99XwNN33Fei
Pq+ZfalOgT1SyfBrjrV261tAXI0sTFPFu4V1cLBLmwlRYmtgt/3WPDpjZgltOlQ0
d1kgcsAEZ1h4Vj5CBjG5DIbOUt9vpZPKtLtnxzqHSO6cDXu0+Kyf4a3SwpbkvKbl
Bf9BWx94WmV/03VVmhfQ8Brn6AGxdraQPTAaCRldPGnaks8DgMNOOJgdx3puyO22
gjWEsNYb2bW9QkhMP46iPQiFsD6kbkUf8Tz9lIcYPw/TTXabL912m+u9xnKzJ4jp
8lhyJOb1syOW5UMkrbxQVLjsmDum82sdtXASEub4zU2hNRNnYP7mC+99NOTqOOvG
KLcHqOsvcz6Z/LJn/Yl1/GkeRtekiBThxaeM0cGti6zIgdkF+3a97zU4D2yKs72g
wzAXX66dvz4vw024Jaf8u+GJ8Y2z3uoQpScD0EP+QKeWwmxYnZ+dVd4xPjCa40Lm
RObCO/pHf7LaOCklF3blreLNKkfWYIb/YIhdCL/xkyJ5Rg3ExpCqA3KQNxpHv1lu
AObd3wJ1D78WAb+4/QyfIWocT4J9RiFVKh88j0+I8Ul/ukKzyjCLVIOegcHop6Pn
yavZZBevz5UGgt4JOnBtmXQT4ronJWgYgXTqm2BtJWsCE97caI9XvrJc4Q9+j3wb
BCqNCkBfGwZvRcIqTgvvK3ZYLDS46swgpiJbCg1xEgm9ZPmdG7t74whTVAOwzqib
MVnDdJAFkNlsWJUF0YDyPl9gvHrQArOc/kzJuY3Tpk4aOpAZ7wpzKe2gLyNCLtjs
UdRexWyEFXUj7JWKLiqxTk/ETyR3EpZnWGmh6An0HNw6jIIecPk+WM5uu3dX7lpP
PL9AMt/S7wfTxq+iPlHRITgUMKZE3fpmzN6iCeAv2HiHjr/3928R9Gq4gP4PLIRc
WC2HFj1dOhVg13otYTaGZX8i8XQjOVesDwIZJBJmUpd4fhm6kTI/aTHzw2O3I0y9
Px4ORGTHm4nPBos/2n/yU/Fn68nDV/Vh/L6qHZtgA7Sj3ndfiZUi8DYApb2RXfYX
HzY5gigm4fMBHEBT6D8mCwDdOtpHwhmF4Ehz8B3QD8PqGlAhXdgAS7QESKTBDAc9
qW7UB12t8nRBEnSMDz/oCKsPi/AmDwxU1GM5L5SQYNlCpPLWWDk9QN0pSE0NzmXi
MkUFIAZZS9sn2FBb9saU1ijgQlfKsBZ3x+uE1ICjers8BBYabqHnAhS9dPHiblL2
q/y8UhP1LVaMFss2nCBujWdoJdwuBlfVhZX6HjtIE3XIDb4BKGASCOD2a6MkrmW+
cOgU/4WQsVtmb3ZvXWP9qL643zGGloxb3ECvb7OrE3chfqvqvD5zyXmw+jiO2HoD
b4lqn3mn2KbidxZtZmhRSDpnAFQbpq9kTa1NLJBIDs4MX15vVyV40bWo2LAyI6+k
tNz7aChZ3pTO2avEvMgGhlpVPxJDlsZ+Bq8Gdlg77l7wT4ZZdxs4sFYk+0EWbXOc
5bQ+Hs5c6YuC3nxEgeLM/CazSFShq4LwjPAwxVd2pXLWaJ5u5/1pE1gw3Eu+vm6t
UG8fjJDVbaLFxCBlTC/bjEAnySIaWy4iEB83rGqpOuJbQUwP+7CBqy/O1pDh5R0L
75hPdwPH932svoFX4uHi9Sa1JrS0hfWDa0D7f7+VD1gzWry82IHNNWrIQ+Bfulvt
urZnk5spbcOkbTNPnaqjZcwCvIV0yX3MjpUcADHSvvKFCM0+t17CVtbLEdeE3jR2
rJ5+rHEY3iGrrY3cPgqXZfBCpBfl6Wno+ifvxUck8AzzZpVv98ScgQYL9vNU6GIb
zzT93SNuE9nRXAf1zI8sIsjiDoM7IgrnXFchs/of80Shzp4EbmGLCl28p23auI8l
BxJNTsZd48u20s7XONGtrzB/tC12+w1hmO20UbeKl667XtIPEkW+PnaWyuc8ZCxV
fVROgXV5wIRrsfOih5J3cD1kTD0oeqjApXA83pdwGQQVGJ0iuyJWTm4C2NNk07mb
0hP+IdVdKktYAkEta32elG7ocskrJwHOaRbC+Pg7I8zi8K1RT7HrewOZBPEw5XkU
g+HPFcaOeWnky8tHnh7L/NQ7/dV+WDoiojcvkVl7ZR6gbNTIDa7vKOiECOI+uc7t
UV4oE6L+YewiBnAqD7v1ifYTnIaVXuqHmgZVw4UwuUh9gLPspWpeaVLXm+6P2iCH
cks8b5SeMZUGh2Neaev4DvRu8WjoC/3BDrvTDyP03V5AMFFKmG0IavjkI1fDHiaV
mW6WoBvxKJRcaxJNP8zSt1Cmk2fte2qAU9tnZM29dlTB7PLVLq6sLwEs3cGdFp1W
rqrqUJmyh0NVlY68AzLdHsAyolmeRjWZar8NQtuQPjCYmWvHkfJbr6aVu0QzdFpN
aYHRykv0mt9G3St6ufBn3lUouLMl/8nPZyPFQuAAo3d6zXxRDThvolRaH2Hh7Iim
m8oKNA04wByU4LJE6d3qWRXf8mVF+8zzbUNqpBnYFWvwKzcQmNM656aFZWdT3YHo
qgPHy7eY5aI9G3zLmLWW4YWHZaGTh9eJ3c6XHB9afIQQGbsBgq8ySqGdnm4E1VZ3
wsl5mXPDrvqwkfDKMkWLZVIBlaB0rZ1pEVFh2xp4vx/jaK7bmlUTu24lNlOxlw4c
NqnNB2hlxva46ZE6s3qqBHMPsD8Efk6K3GNeGiaXMQzwFrl6GISQ7VO8XwT1fExx
Rea457SG3bGoz62HvGka3Uy5yPNYzs0XoEXFKkMNShdFHLeoS6Tc333eKK0YtILF
2Cl0kuhzCWjXDPSCE/Pg736ND/oXnsii35sCxtqf/jJvE0S/MEn0uP9vNHPo81gZ
ERlwTEnN2WycpHQg2DwGAuQ/7xL3EizdBX9TjP2D1HFxOxiB/AV+YdrOnfTT2dDB
A45odgx2xGYcU1KBvAgp0FoaCWj9Q4VYPEYXbSPlrQex7bLvKancOeGbVRjIcte5
rDIc0X0UPOJnWDs0ioZIAYtkenuSStmP2k+zztAr+R+RcxJKXNziirpmwkluvAJa
+BGdTuaPzvASvfRqezTgVGlqgYWMU/mIb8G5d7Ps08tKC4FMIs7L2p6zaiY5XZ8E
ps/qyi2wIWP723wOUMP3CmXuZOupr6tmrsZMjp8LypcCloPgdQX2RAhzXVy7KwU6
Hb9l3qHcN327JaFLGaduSeCS3H96YdqjjNZ07VGmyt4A5OMgXumEDLstTO17HEu+
kFvUr+EWaqI7uD4Co5QHJea1yOug6EsVo5SV6qoKTNk0g+wE+x6+zIvY9J8ypIba
yCEpxhHvLb7u8373Iy34ltRq3HWZmuQFWQdd6s+zcGx9jDjeabEQAz7RXph5es6R
aDwzt9C8OauS4NtwIKyEZx9ir2ah6Dpn/kUOA3FjZc7x3Ep4g7Qzg2Z3jNHTVRJi
NBmuIYsHn1ZnWKO+XCsV0FFEDZmyRdTceavdd57hYtftWL2V3f413aLZeqNmDIVY
4zjvdibV952+Io8VPYXnYpVDxOCp4zPx2C2M1C+ABiokqZRYYHg9ke1WKie9bzqK
22Uj9uI/8yH7eN2fCD7YwxmgYgTjTpXN83wB8IPyuoFj/g4kDFtYPIJTwHg8eSHw
jTx/oTAFRmwhP/fCDePDJoLRiBM+BdQD3zMapJr8u80BtmyFJxzGMx3BL3v1r0Jj
hVV0lgeyPOUafcHaXhy2Gmkw4Ot2x3Rs2HNHoP7zuTA3xeM56mhl5XpSRrk3LJ0g
xOiUWczPWCBSuRRQPVA+W4Nk4jXswYHHDyE86WiKfqCA+gL1gwb20B6DcbLGyEwG
TSJNB3mnd+gc/CjbmWNaI/SYB7i4G3l/9aGAtZZYTnu53WdClvkAJhrdgjE/LQzE
3Z6o/TL+G1Iw2/hqZ0kgT3eMtebooU15jLMnD3qYNlWJvMb5tmXh6yGezZvO2v11
ZTOTkbh34deDqz+Oh2NLG1hlQd0cOAmwmoaViTD78fmPJ/FXPm8ihvLUaA4l7gj1
TPszqgovdayQBMLx47VKu1QOetBzugyis8e1IT6W2/0VllaMkuYkwGM3CV4itbKD
YhkKoS2lWx3DTh43MpqportJqE36k2OQXxc6YlD4e/nF12Lx46cM5gw+lO/zETFw
Yyzv3lmnguQ+qcozEysMlUfl6PVXczjlCWbzSKZwCiNN7pQPswAhngDxnz7bLoBU
d1vClztbjOn4V7p6M8Vj+b3TP74S6BnBYvnZ6HQD3EZcI5YEjAYYJ98YsTrKmGyD
1ENHFipKcRXaO8H72r54F2yqAQAwgqRWLk1QvdRMDV2c3ViH76MLE3+FV+NF7poX
56S11KRM+gUqjfx1cM0uDQpqkE4icY/5vKKQPBEtiODrvtISybI+wM2TQbysZ+Lt
PSOt7nAsZN6oXHlfZ09IxuwFbLSy31jCAMUWPPkgj5SAK2NO8OQN5nx0ru/TRKYh
GyGRMjYG2PyvDCv1QQNIJSVJzwPsfK3lNF13JGbuxKh/DIQQxj/gm1JphSW9cpFt
rtEScWCcNG281T4ffIrUWAhrej+rTyB65Npoxe1bzsbVv0PLIPtSyzJC0ZazR91P
uYHjv/KK1B+bFWeRNM3mlf5LtznnzTCA8lkBMz/Qy6Z9UzWm1wmv1O0slqnxgrCs
Su/P794IBXu/RZVE3K4Ym8Wx+vLkbQP6+nWNfJ1F/4xSCOWoLL0oCYn0iPCAPUo4
g6wbb87O2CiN9EoW0H0mC5cgzw5Xy48wK8zuTa4X/w96ofCScTHpVww0I7ZI3MIc
ZYHc80BcvHBhUrweCUd1t/RpyfbPESm6DzSkjOqbhFCxQ1ENmorosVif0QAeM34T
x6Gk0UDs8sTbBdK0K7I7Usu+gwIPy+4EDHBX935ozpL4C9j/6ZIFd5Y4MKcPuikb
0R4lfamPlYdYONKk2rigGLdUPZfeU0pnrBNZhSEaJ7gxLIvRnpkz5WWqk0k+zPrS
qChaQnObY5Mj2sC0mmQ+3FAkMReJemKmfW8QuNzzq1TfsBPMeo/j8cSkjfoYk47u
+C6aUXvmrH66gYaQ5TkcAUMPDudXkIBUXe0D29tHQEo=
`protect end_protected
