`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
bo49trehcslJg4im271Q377QWe6zgGpw1iSHXV61aCd0DPUB9+U5vqExosmwglnR
6EIdorVY7zsfjqPqoS50ljy83z3GpEMeWK7/xAiZf9jImF+o/Ezj/1WPKRAKtVz5
yx8elM90r3yDxSLwGdthmYnPTuO++Yd1iL9oFQMV68GruGNnFuVq1XrB8Tt6EVye
vPGU7Q4gMNrvmlvEgevKN9Bs8+lgi/PKkdBpc9AW0dPirKg1RzZ8T2Wf1Mwp0XIH
YX7d5mHjUO75tWGxTIkjCUfGHCJlMvKz/K/WATUryLKzdtriJ9WuggQOHykb7lRU
fuVQKf4SrtBTco2G05uey1cwVdO3qWv7Cr/+5YwcBHLx/T/QcRdAFM7O7r+P2oem
dweiX6K7Tq1AhTzaP7yDeNV3wIgvYhgZTlnQYroXGbzaJ9WSRzfprvgCFU38neYA
K5R2qfBrq2RUVcq/WncAWXIWBqDFgLJeKVKVjLZlhZGNWHDg5D9h7D/Euplwp8/z
kUnvrBzWleQnWHzuNeBXrEzgBTmAJz78Kc2xjwe7/hKhLmp4mzPZ1YTVDbyczaFr
TPkN24wgu5lGRxKX+1Nl+SlYioT37Mi2c6OB1EYgLRd+lg+v+YhHZO/akJ+BvFND
968Wz5CHRzcLWA8lS87rx3GUgAaxG6aJYXZwMiNeKAayYcL6ohQPO0xAy4sgAZCA
AObNur5HL9JfBH+ejzGuSHxsws9Hx5XlXPqCIj7+PYdQz/pfaw5j86KteutBwG6U
twjm+lEA4GzCAs7lN7LsPTnyQjMJNGYxUSD7fikzyM1sdCHolxkryqg9XpmD3sHc
8uMsyh6scSDSZIl+Jr/YOjDQAkrjJZZw6A5t/Z8P7MqMysj8gLUHm1GBHhNRH5Rj
hVLEowhaVmFYnMSKj4Ff15RmnKXbBoKgvSvCJ7J/GbEiHvqc4VznsV6Xg2jpjhze
66tQc7tiij8ilKbgk/laLmj280OElwVfDdHJitu0AopcYRbvFjG9nPjLnmszelrG
chkWfvA73HEtSp+Jy3su3fI0YXKStEEi6carBT0IcuyLZeJkn7Vd7aL8R+rC9FaP
cTkjjWUPhNNh0+FbsXKvI6IZaMG2xBoORBzz5b9HmRBK1yrNHX9/+1cw5OL7MJKG
Vn6vcLE2yGaXl45asY6tgmREaRvMIWBo0ip/rHx7mfW0S0erQIL5ZA4ACITiRwpy
Ca087iFzH4MyuWFbcZkgYhNlbBEWLb1WJX/fhXnfdGgkiNY1D/OvVXG4XfizOKCe
cvdrQF9vY/LtNDv13MaqPbgHUYRG1CljDIqKAq6RBXbtOk9krY4oAdwnd7UPFmXW
OaGpxr6Xm6I5voTX4oVKGh+JW5p5Yvf1axaapOvF5mbGHxxmTaZp5F2mpmKasaO4
QhEoPxV30H0BS0SNC0wY8oYnQnZgwvHhr+iOaFPwwfCB0NbT1WLi8z76nrGq1XvA
pDQWR9xmKGccaMbKDzpNq/uSoqc7lmqYR48KzYg9D2ylNilrtKst5ASTyoo3LTUX
9lnvjD8QYN8lehwDyiFm2EVALpNWBcjr8kc7Uy7f9UJ229swFlXMo2cIOyKSB5qX
Rhlb1EcGzNvdLHrkDefFV3xb+t5fqTT39adb8IcQdUwXytMgfK0xWElnPvvttJL+
or01O5Z20GYcvyF1YX/tiEUrR1j7S8WcBa8TxxVJdh3tiHsVkI6z2yHNlTjrdfSZ
8ZZqjOntvLbTl/+p7J3DUlECgdDTpBdgraRXNN63e4DYWlL4+dTAWcJUfzPdQMgc
TWntgjCVaHNq8W3d7xGKbOnPgV7wvwY0YupzjPTDapiPHlnDVbbuWxtwwWooeqqp
WAdsMKflurz675MXwFQhe96W45c9ZpJHE4WyI/IcKhgV7e4PTzWWD+nFfxCaopa/
Wo1QzR/jVOh8m80Y/UYj7TO8aURwEdxx71kNKiCYS9kG/eCK4I/vhELP8N2bHuBP
+FGcxYySeDfeDEmaB6/Col0SNT0GusQqPjGib6/H7AUesWS+sTfD2h6gAz2sPSCr
Qn2lD1u4/r0LXmpJJAj0uB/ma+6RDmW2IU7ThLPge/UrzKER6D0pSnHpLXAzZFLe
/Ml6Mk7QjTYVzLxkSIpI9pxJF10hCcrIJa4e2fp0FqLe9JFBH2zM1bY8D0AVNkn5
dwv+E9efzle9/O0kZzsUjyk/WgbT2VAgSChUgculw8lugiMzAUFvM4wlx6ZZbt3W
W33xDVAbTylpx6h+Yh+fIwChBXvjm2H7vCyknglPFgf7OSHvmgjAyz6xo9i9f+Jn
PTGe3HqUSMLj/j60fiTQ3a8Bdaaswj38p62bMOj+H3ugCuvZrKZrp0kMU6GeCa55
oyB5wqFdzVxHCKlWpNKP44cZ+QglGFEocqZYzhvgUFwVV/gQwuElE5s+CZmr2XbI
YuMNaWyfcVFRKsk/IHnk2eytklL0ELhghnGuS4k39PhMIg59TQyAKGiEXHMA9DyN
0tTwUAI0mCg7GRbh//9Lc60/SEVaQJVdCstIZlhDeBsyTGscpaZxI39/90XGPdQq
mMTlIvaLJFQUo0TleKZWGN31YuvYyfnils6JG4Ppsy4GZilFW1oDdmSw8QPEtqjJ
ixE+hhpwh2gbNRa61Jph3dm2Il1J5jcx/cwB+NRKLOpxURHAG89EwoNx5cW/KTRr
bkTj8YOxS34zIRVRTLhL/X4cJ/BYSdqbAsSKJuGQ0GA+0ilroJqLKXuCQdfvZthN
fu2qFisiBHVlOFdjunWIjXAEuD05AePV/vmPANBg0mg4YfHUzS/WSHDh6xP22cA4
bWUVsGvzYFJBxwaebZ3qFxgV2FjDp7wxTzo6DcamVh7uJEaB6o52Bfb9K4mhqU16
uNWtHRWstTpLKZY25WlQ8tTejqAM7pP9NU+MUl9zIN48iJ6wOsiOMdht9Wj2eJTr
B3l8N67XpUT9CPkQu/85EI2W4BrxgBwQymGm+FQmh+DQ9FxVBE1gFtkExxWKhovF
NSjs9gARPJDVniLQW/2+Koyn9mWPrHmw29Okldxsgd3YyNwXak/trviLW9wxfAK1
L4FFoNxTGV4XFLKXvyIstDDE3TMLYNJoBh/Z6YXp7b/+0dBTt7XQXWsuadQckbGd
pL+uAYifScWh/yFKI1T+IiAo7LZegaZ4fVqt9UOsoYo7VkJElh5SN+ForeISbvIo
zoRodIuoTcrGt7sdtToL0hFtTvr8q9s+p6O6lAY7owkjL0CzwVzZYFOgPfOG21xY
Ah+lyFFRyGAxClRCO5SQVGgeOvm9hEFqSAsfaY3nKLhqYFmZUWudHCTGGCe8nohb
G3V7fWqY0Bxjx5dsXXdcWepHPzpuXhDoHgj31oElamR0TJAJS8ysv5W9Xat6pCSs
QUCThnP6OwJnZ8Ofi1O3JqIrQ940jdeVzUA/m2aWr0/mGchFDnRCglAdFIuguZVl
XdJSs82dgCb3nTGeLjeioos2nZJhomoNSDwplnBlCasGUVjZluuoZ7BtvsejhryN
jK4YcjSJa9cpmRZGsdRwrG5CYnbkYXrKqTrmeiLUxr5CD46dQn9MMw37w1BZ9IqW
2OfErXkJ5tVMqWgVKbVP2WhAlokZwRu7aiGsZvCDUI1hPJBjIwFYm8JBsci67NZx
BvKjvCvZF4XIeGHbRnbeEDa8MMowlh5Zmq6q4RoULIiuECv9a9iAMLfsStmApVE5
JE0ZmYIgIMPh9DhT1/k4bNd5vTNBpcsYvcPzapbmPyV5c5TGXqBl2JT/mZOBtBCf
z9Qet5OGK10rhtAKyJjesR7FF0bf1Po96A9kbUZ57LrSzvw+zaohVNYRQnnDBClS
qRB/IysNmyoGrPmZuyvE1lNI6afoNln/hv+GMO4cbU/nD3M8uQQnuCTdaiOiDE5t
SzwB10+kyI+K/neDwZ+od+Q2iVPeTTl1nlmBOXNPx4/T5DT3sEL6LBqMKbaRhRi2
0XweIjp8YDrdZxFkBuYv+xTm9VTCeOyIt/5HsqNO8lwM93hSrlzz6uSk6jux+jvG
L4/wmirYxZKe824yeVmtEVeJ4EUZMTo3dpwA83Wx+3cxNLIsQnJw6nSkGjKtbJs8
X9URK3duzDvGldu/Anvq9ytzgsa5T90aTMvoPOkKQecdeuh7FaIFxglGfgmkBEwI
IBc/SMAJT2/pQSvnHs7tthUHpFxdbzGJ4ayY30BhceZwxo5thpiQRUFXrKL23OhT
IZ6ThpmywHvO9ZDQBsQXvbCy/H0a2c+9BrTAGxmQ/zaKGHcLLSMysSjaQ0JCboHc
pVPZDL8YM1BhsIGaZDXqdYeIsIFccPgt9aQZWU+SPhvz15BdmhqW7Gxy4E5eezj+
JlzbVeqdWVRgccnM0g1jPiLmxZeRksPAqCLD5JDDMyw+W9iQiw3MdsR/utoc3lb9
31oKI885atJPb3/ntIL8HDGtl/zxRRZDW+29zVI89A+jkAfUMUyQowgzWj9FjGQv
MduoArtSDm2BhcOiCKqG0cA7KqEhjKGEwnwEf5COx711M3QpqroWwg6Nj6Sv68N/
rGk7OUxVQddJ+qLXmAAwRsU60Uhrcn+Ir1x6ttEZmv9H0/skv5TMZSg35wAvlnSe
AVIEwcBr9gboNlEiUk4ciG1OI0OEjhKPPy5YAdvGsSFZc4l0RZXp2xmmMIqeqaxd
AeCUPHswEB2FBD61ODM2J5CnXJtt4iltHUFRNGbEMzs+ABz7/8KJl+34irBxAFQc
wCJc+/fHjAEHiIJjdk8TNDzMqtfp1HShCDq2rHAFMTavdSEjxsgFnlfiQc9mZb3v
/a2yXHPdX8ZrBqg9eWXpWm5ht10j1TaF5M5/v9cmUu+rnFmplnVB4de0Zt8MG4W0
OQWsj1+6834UCsM5LCoSEjHaaGvk+A2Z6FK9wnxw0oT2vovYGnvKOD+VxdSdEPul
u/x3R9eqpkzJebVVPEir045SaznSLobDC/hwcemi9ZHR/3gV4n4sCovziLeTi5DS
/RnrSAem0NlF1FKdwjCZXUuk7reYedFPqSW3qomLvWt9+HcpGTc6e7Fg9yfj1x0d
pF0n3Ly77ENOWgKtrGZMW7GyDJ9INJ73p21umLrLhQNkJmphZFkqe9sWZJ83m/GL
25/ZLMVAOr9CsraZ1pZRrVgw0Z2qeRggTJnrvoMpJsE4ajUkGE9Zp0pJ/mc7Cr81
v4XpyPXMt1fVrd848gn1pf4xenBv9pQzvFVrBeeYImeTw6mGyHZSQyevZ3xgdpai
0vGNJW9Xg9PU3MhVvLxKkthYJ1W+HJEnExutQEkvtSz2FIquUKGWijW8JoUvq8fO
RdLKCrQo7TUj3E+qwI+TSNDxDeE4S6y2gbQIGCvY2/jo+VE/VoUR49c0qHkGWVN7
Hj65nZHeZPoSKLtNF2mSsTPGW8LLn/FI3K3jjUNmKyCV7R0jKKSkWkGqLpnpkAiI
Qy4qyqW+oUtclUket3nV6Wr7iow0Hbye86GRskkZdyIccyRNSI3Nj4jrWKmBH5m/
VGBNtfzPzuAIRNpByMcSf2pP0rcgvgmJu/PNa18dVlpRMhoyIvKHpBv06J3xIx4n
ob2pcjUhqoqUdyU+Ucho/sIDRXtSfZH50yVpciJDMGEyXvFU3BYTxM8sDBhC5Tlf
k1rCSugWJAitv+Hbfa7uNwl2kg1uLODuOjjeQWz9Cd8iRHO4LMW2zVAs5wqTASch
jCPQrajYTLZG5cbS5BVVfplx1aQPeSzMoqdBZcHtG97qEuYgmWScVLCr4/RYQYJw
9AUPtoZguJez3In3joDdPAPbEWiGVEABDNOL/oIeNGrMfcYGv0NOAB0CUMR6ZBdh
cqWusCAECv71TkPwZvbQ6AqwlJpEUvRaPPF05aegWaR9V1f50mkx4tVdWNWJS/B4
R4r8ClNVuSwBombvTKyBZMqmY7CRFmmkNEDdLQW/OC4kewjkQNJjejwZ98tyqHVy
IZIxCUVmidBZwwNFIZ/ep4E8KswGVYz0DC3ezmSoRRACNHdODCFL/XT1OmnfzfW1
VLWyRvgRUFowzKCI3B0Fs8tWLHQqCS9/W0swEEwr+xywuL8JUcfvtR9jRTbnEDan
jy15AqkNaA/cH5yxx9x2fuisgRygdNu+Q940R63CxbX/ZlxA9FmmGS0dVFQxtxzo
NX03uN/xSHyYMav/7VtX++DOguPqcABsspIpYRRnVOlqUyVJ3jP+bs1y1iLYbvI4
erMmcrJPLFm+zXtZZ/lLsJv6HBN44kBFYtISRFLn7Q1u1e5fwYD2sAsVpEW4EUOm
8NZmE+izh6oBkt2jbBKT7FkLcIlGmGHfVr5cTVeF1jgM1K4yQys/rvfxjCZ5rawg
EsVXIQVi9KnStCcAf2Bfhs6HXiwb/xDxz+wLCQn7B63UNRQ9tIaRENdfX3O1VO5M
TgtQAtXRA7AfR16Lim/hDvxenuiGU1x7rd6LK2BK6kuEUyJF6TJQBJYdluMDVF12
kerQlUHzVjHJLE797O94d9lcD4zfrQxzO+e0RdSdp9lT13TzL1qZWvh8Gk0/ZyjC
T7amU4ZnrxIqzkz7RUf9RH7w3Uce4sinsqZ3deVpc27qjDRnQX3+wB4qijeLmPKU
YepUS+LK8da/SCeHd5WWAnTS8eWxri0h+2eD6JD+gWj1OeMHf+NDtfmXGNN4Ipts
qkcXvy+A3yGLD1jtCvtu2Tbtxti8KtbBD1z6nNhfGSJaFiNERrbCDaKf69wBvO9E
YkOnvO2rrsQZKwORnla6LdjDEb6twDuKIxokGmKVae+xmnF3AMcYMYnE6v4/mmYf
RmT55PhStm/rtma/zJ2VKPUjXlk+TWLcIMrfdJPYYdHLJu3w1Etcb20TCnj9Ygut
+AmAV/rHTCBbyuPMy175ty85V3f45en++SN7bZxkAVxzNc7814pcd71tG9r8YPdj
1RAxdBLmjSK0t/wz6PlCMI0FKgZXOq7E49MYfGzuJWD9cB+4N40UWcb9Ep0eNolR
VwTRpi58OqAiVsZnR8r9TRAOJFinemSwDDNg3jPKbM0Elv1ojz/V66bvX6/QANZo
L1ukT2ZB/I/NHxVnQXS3/LIonE88p48XUx8PRON2QaVpdafqCGHA3BTkJIaCkfV9
CQ8CmBradUJvYxBss6jaX0HGyrPO/qMx5zPGBZ17tzF7TA8Y12BplRW0d5jUqc4j
meZPlOrM6EFMA4mXajmbQeq9cIbCATPMlLbx4LNhHccW2owdMOJPSS3M8GZ4zYsw
GGpLPe0JPgjfQIUlqUkjDHnOYNVvNmZ9fzobTv8X2fBXhEpOd67+JejYbNvSzATi
ld4uFQMxuvk5LqjAvYXO54JP2cNFvjs/P6Sk7gcQm6YgHmnhvbl0Q78/rRBhXROM
ZazXlaQT5VmqfoMH2lYfWvoUSNv9lcpxfjgJzX8jSxNc1uVCpWJe51g1HjEv0Tsq
sQtBu9l6K4SRGyfdIiIfCQhe63rEAjuQObT3Uvry9nR2VjfzAfG17I5Jp22JMDZG
2EPp7qcHwphIdag6ahTWTOaQFT2C0fBh59Dln68ytVBDcOAnCe73tC1IdTeVoWc+
k6On7bDT9nS77heGfll1I1tWb7Xw/TSxblERUj48YB6JpppWIjf5iUsi0zHRTYAc
4g8iU7fL2fFdQVxxbMdS5JAEOFkOhrin/kez5vz63E/ehxE+NiJikrGbrIzYB3bj
m3Ap2cjYeGgADHnYPHWa4IWwizlqZIRmYKBFyYzjorD30pi8ajVByjgGD4advCTZ
LQnUqzKW9vh/Jq+yeugkhC4XMXbLu4pGanobQe2caq0txrUBIVjTmDuNpO3eAQ7T
94hJ0SxxfDZaasTjMDZckTwTzwrQiYcTGey6DSEeX9ymf9Ve19SUixt4hGpvqTHC
IPQKiDdILLqDJtIkS+sWJqEEdKJTaHdwZb1cM+DNRtUUj+NvlpyYgMXeszA4iCfp
j7wV8JhPglsk8vsQq+Vy1taFohfkfsSwRCccaXHs3bWkFewuIXL8PjP/3xEPFTLX
Cf9CMWHz/VXK9vDDdftjUHovh+p579/SGStn9/UfhaEccZ2U6ZI7f7K8nr5GAvs6
e9gih9MXfYitkVtRc9RG9+n1XgllMSc50pl6M6In49FPaNsSDiFsiv88vxeN1MNY
hXHVjnHnBZM2SuZkkQ9jMRfWv5VLMkX28t2yQZuZWZBZ3Ir3+NvQ3Z++xF4ZKAGR
Z1nUUrdyPrOBsDyiJ6wVXTsgcIDrtIUTJALbt4df3Z+6otPy/jkX9uLahrrCmdVO
hRE3zDt8O4gI/3FVOKkEUTmmUyuFiLfxeJmVMmwvJTUzU63lvhsW5qpvqzxfy9hV
VWltfl+wjBvKJnVBumlpFtrV977632m5KrD6xz2fQM2mM6MxA9xeGhYe3J+PZBwv
JbYT7jNlRjjtnqp04kU1jA9o4zZN1DeCDNZ/Lcnl7fq06iTbKUj0fd+13ivfGCB8
JLRbqkO0VMcBj9PF6h/w+ERZbu4d6qtfa5ebhwQp+H3sYn316D7/a+J4KncLiTar
oyeWnGUB5Uz1zmW9vjljU3NCGvpsbWh7rvvdpyBvac9NtZT4Ua+QPaCWGlcWKjQm
nA+nE0NuXNnESiKZuSxXTZ5DfrDADGQnmf46kDgDou/TegAucVqt44vohMICHXwD
+CIvHI6dgVZ/sawuOnqV5gnfYAyNb1PEFAxyfMWwFQnxLm/J7Sef9I07U1yMv8G0
K3QFW5q6h+q0zwokKzOFJN6XPiw0B9ZUCxRZR8VwDKWozBCFra+EvZG/tfD/DdZQ
FwsboW+fBhp51ACKaH9roOBhBoGyZx+iqR/NfPfchlAnK7Y8ZIkTACsoUw/Ayttn
uFS3RJ3Qr8iqT3U1au7jqBNADQ1948iQEePUIcSxAyc6SkeR0CwGpdD8h3gHetyM
a38RhOkKpzt2jsHdEmjhHO/+xVzfVkpG5L7eaylD++AldhnBjy2RO/Dd+sKVazCI
2caJgjSsryv1vfEASm7gmHApqBL29Oz4i4CBI7x04/y3YIF3cNjYqi14bwpcjzH7
0bqoayOnX6gZSt6NSp4oTEsf5qkK0+kipnuw/Lc7zFzMU7T8Je7fxWiNqYM3FWfk
WHCuuOdiI8ggQMsapDYn9wT1wAKT8EkacpXvqYpyJUAYKNiwdQ5ua9TBcFtXtc4i
OXC4UoisceMBCxzXXzu36CiTCNttspEB7FqfmQdLbbWPwJDRy/89qtTdqEIN7KtJ
349wE0K65sCPJjmh0gTbTJHmCt+E+u1mFV2PMLEu7MRuUBVxsZz7ZzzDwnuUdK+7
CdGJe9Uqzw+6pq19tVUDpqznHPvrAGosRWPInlPzcm15+TuxmHcwi1c6Nl7wyS1u
sEu+3/Ey36Pm87Uw23bKBuEc/Vs3CnhwRsjKgh7SDILna4nBFY8zOObtitKSl4h+
Rwo0AK77bDS7JSCerY9Z6+mWUbGVpRBUkJGQtQ9AY4AqskeuuuJWg7Oo4sF518XV
xcFzklpYprc+yZNwX8jZ2ZR+yZPTU6QptHL//+ESEtExLLXTfAJXGor9yL3ESTit
vBscjbyeVaz1ayqaE3sWqr7waftELn9APtHLcImBuOY1SFu00polj8yvw8+adrxj
oTsKO+Ig3mhIcrAPFPlK8VM4ou++n5gR8TCTc4ODJeG2YtCw6JLkiOcwu3yr1tpE
dEQ54jjDxU9pAMbri4n/kWxq+5LJCJHVntzAnsUWZcKpg3h7+hCirXchT0BoMFrr
1Cjm0lWZ1ic6Hg2XZzudlGB4H5G1eAfHtrDug1DzdbZS8I0I7q3h+5IXA7qC6YqH
3VmeHKnUubsjOcS3NxAExXI7TtDhzI144JxNRIey74XPLvwPaRk8n8aQgbpQ9mn6
hoBWPC6PffI3cfEaWMjNUrv0szHCq/+zwEAmRW38Ue+u1BGec4DSngsykVXe6SH1
T5+s7Llb76xzjvJ8wHIPMCIl/o4295gPdGHDZU33xiDOc2Jgf7B8Uu1yEsIqiJ4h
J7HOEbh21KPpyalfRWdaZpzhMumLHYbvLfe2eW8k11pDl/2F4r/HtcRCvCemU5wn
iBvyc9F5X9DhIK+htjPJKuiEfFR/t9bv5F0DU3c+kf3ZQ04duP7+7DN6ih4hSTg+
kzfnGXdBVQcIA3W9B/pYr4TZqVKch7PnhMinftKjKtprgyBWJiRUNIVmaj/9IVm/
3qpR41saAABwE38LF68EH5EkXV2fO9Py3XS7cVkBOReg5LCJuMLIrXCzFrlXHnFE
bsjSPj3phq/e3uJWkEG7vhq3vZU2yTkdgbP7g8qKIZRWGCVf8Hd0Y1OI3zBFgjcn
T4Toi5ekw0sxusivhog+RxI/hhkkytycTFTaeMJ71xqSSDpb1xjbU6LIBPCDxpqf
yyL9erld+B4+F0gXHhmgagxEz0cG99ChJvPzeys8oo/psVzYe92CVYJAkoabM2yu
o9Xf5Xx/wCrl5yKIbEvNFuC6AuMeVlZz4Vn+VN1okeGZ7oW1VDZ/N3McjWtJ/rOT
fF/wErIB7bE7z4ELWwZ4cwrAJbipP04C90DhxQ9Xa7gw1gWZSzoLKKAN8Y56UFG+
N8JA0FkBWAZIjgAKEY7DnUA32RQ75NXFYtz8fehRdqR8z8N4TjMVAqkRNEikpTc1
QOeAJLf1tqQ8wH19gXzpueVE+tBMhjXoLzUWICBqjoqbrtRnfDKnHgele4AK8PrA
iexXviw1WqFq8B5S4XUJYBNt7gcOy4ulDVzVJ0TjSqukW8lRU60e+svvoRPxur9K
Zo7a9E53+luSKZSkPb30lHB61mnPSDjgHl9Id76FYuW6Gr6kUT7x6VmBIQHk/x32
lgYILddWq3c8WdpyA9TKm+D7xsV0BYrLXWkeljzjUFJH8rgW4SYqfQ+iI5JZlf7s
V7EK64j71317kmseu/6M1FkIYRsbfDEO9N8geEaIulm+GB55KoOG8K26kiIZ43XK
Xt07q5kCSO27CHX7AKjlqmzp+gs/ZnbdlNZQKjllu4lUS5d3roPNPZbCJO8Vloru
B3/z+b0oKmGhwIDzIDe92rSIlp5Eh5YpShd1Uc6uA5qw/IEqxZ22JIgrmglZFWqY
bh5ah0jp9sU+ZZACt0FJFsSOjBy6kJJAy0uLmhybUV/VRshiCbkSOuwUKcY8M+Hl
JEk5q/XwqBxH66fYDTvkxYfqYxKyw6X1AEwqHrijexVLH1yphkPkJEo8nfv3hqAl
y9H7ROx3et9hAzRiY5AiDw0zeqVvYTjqSlaB5u5d+BqtA7mS14X2OTkiC/Ss9/9x
eCP7+9kvJcM0ihyicqXuxDJWmr3mCrh7/06IAx23nxyFEfzi8W8pJYxuRrDrHyvE
OMpbYTqathUVGMu4XIbVmKxuDKYmNufAO4X+7Px6csosHhNeMaPJbz2nyCVJ7wvG
3yakCG1uidELt0UDLOJNcj4Z8qoFNzqKDuP7Wr9P0AIUvoeFlzGbBQmjqsWmONm9
SfYH4gViZ/ioAVN0Nkf4QguKQsSoPI8pSQCAN9wqLuxMxG2zl/X/5b76+pmUkobi
gzYHm4SOd72EOV+VL5EBDM38icTnMq0Pib2gTGX3rNYYHGWYk2G0DSYu8BR+kX0Y
hej4mudqi6eWPaRQzYfcAXhLuSLH25nJ0hYSFQCLniA4ZLy1j1ix5+Go/6gleDCt
MkNMUhDgwkzkBAw0gNpsZnQ7zRokLvEHfkEVLw+SxuiUeZhURRkKSFnASUh2SLL3
2PqIxXYhpd7kZ8BdRAvw914UHQ5EApeYqeXuVsS7uJsdlTSc7whuLST+N8MurxYy
jdRNsUWLShggVLSGAi7SB6E0A/yLWdSkVssw7lwcMKyQyApK6NOGWrgwnXl9ODcR
C1Fbt3ewMu0iNwtQZH1SPsaT4uSil6LaJtbAVSz8ge4e7b2rc3LzX92e9NULabJl
J5KHSmT2oW3SEdSbs+jmI2S9wyjByvdK5RWZ6qyzKHxev3xBGkAa+Zh4uUEhBpLS
5O2XDXtMA55gcLYLdq8r0EmTPL/Yaim+3OfUQr7LOVycO1S7KmEFUcWa2ESJOPNZ
1AVEAK7JyW0hvJHyr2Giz6+m+f6NiI4iuGTo5M1HMdkMy5OLM9TLKw7+KzJ2Zegh
mThDWyEo668OnGRQa+TtoY9liY79A0ge98nQnoLS0Y/WBLDOWkRWuTBzGkTCYekt
58g8lCwVV84vAImIaWVRa+aRlag/i5MFBO66MUn1NtGYLDTzpyNpJ2FawWtTD7Pg
wPd0cMH8NNMae+Qf71/fwiU+a7i8wxik2JEK546eESc/tzOAUZc1eftdquSwi2ZB
TqHAcPbxOL/pyC3Fkfsh/aDuILQOMVXMjps0c+hMwYG6ZSXPxTttHqMcewUJa6Zz
gK0kENiMdjJ3hzBE3a1/sXzZ658p53PG+O7aZQkLa0iqdwvFm7OFAalCOpajfBSK
w1GLRtL3dITVBwaVuVoB+jR/cUjwgbDsvjOmCXZAoUGR8WoX55W0vU2CNDks+yiM
jmR0uslLb7qkyRP/a27UX7ObGItUwVUTvAZUXn+EgLBEIDmST/akQikMqhC6Oqsh
EOuXjQEwjI8Q1bk3FZtx/yaUexyUt74JQQcGxZ7UyxU+eKN/oc+aa4GJEysmZePc
COo5LQh4NaYF7i1iwx+84LFaJGI/J5L0LtCKGRyl59snQT3PUxSWSYt2WgXpiLIH
aRmmcCPJvg3jytB0/nBH3TExASAScT6hFEZgPP5QRrfsIrT75LQ1UaQNwS+yDD5d
wcIJzvqjcZFYhKhRPmErIX+j4ESzCG9p5urYkC7PQRjzqpFJVdBljUdGAKpugGhE
voFqeOcVwt1r5vqGy57UYWTI7itAJuGBbpHEpIkqtYvlwDv6voLAcgxGnG51ZALM
ihs20rprXUyC2M0bUautz+ag2aahnZdjCRfKlxKNkWAKi7B/v/2kgXSeIxO8Rybp
5hFtJHpmEXk4ynZlM6bO+O3YEjf6u8xrfqoFIMfGODRNvK1s0anqRUXO62Ro9LLE
gMb9G7V+omsN++m8rgsPtIV3Yym1s3I59LBspa2esloOnL7pyopj+FdxZZX2Fnpo
k5a5+utojKjk6KkUTPj4u2L5mxkZR9qOxfwlQO4SFFRikgVK7UizW6hga0vShl7J
b2TLT1EQ4DeRh+3RO7C7z3SoAiKUot6UA0pm0Kl2w/DPDD8bRP3+zXqYxEYdnLAa
OX0bYfmIBWJmEzy1eUv0SRTBJIm7uTdvuEJOpPvBIcXRXCW0LwCh0cheBBeRBiVK
DIrUWMwEKRlUdg+oPcF1oKiF8QTGxIq8U8TaI8WmnJrKm6SKqfyh43xfZHoSAOwO
YPIFrnsYHfo+Jj7acy+MSPzjUJG6EtZQ08z1Prc+1Bbn1NZ3hSmaKrO63WFlEO4p
71fvjUOQc9WHe0CIOWfGveKZlTaIhPGg6izc7tMhT4QSdMRaF71dwFkpK67BDRnM
XuSFSccMjoYm2ErRSayFru2aDRp+h0bjJ0DCKrXhtwIXny8AGCFsmHYNKo2i+zfx
2E2sZDDLUHdP/5WQzRjYBjOj8ePQfkz07XPT8lC8/imI9PXZsb/WFk2GHfrwtHqc
HIg4o/D9BwapeZb0CoMrXQ74sA/g+poxqk6oZHijwFwnF5P7tQHruOcBuuIRrKGX
Vkf4IxvMWmM/LogkJv9eWU1SWYAj7Zg0mxCbNNAplN0GpP1sDeKxMup9MCl5t9FA
Y48qIvgVDf1OjDSUkm6fuLjSJii25aCuIIbhdL0LwaP5fgVI2Qun40oQDJMkj4fI
x5YPe/PUp6tebRleW0nZjI5B19e5K5/grGSNfKJsRI2WLNdmfFyUgPndEd/cXvW6
9aAxm6yAZ5bQUC7lz7+eutoZK2esKQ61DhIttmpfCY/jeiWCiz+Va/Mk3Lr+WYEx
QJQ5LcFySLNAsLmerHryJyJSRZy8IOq/w24VIULAJxjzRnLOqNhxDdNeNvqv+tMp
Ntzxi4WRQo8m5wVhRbW5ukexoaIlVUuWqSMlzn+EOlZOeHnGm0o1RAsmiGUqqHwC
kVM3gmhpnkvwE0vwt53s2qOpTYvteDCCRGG9GdBiaTuaY9chG6GOTzpGWmcKM4UQ
F+lUke/VG0ZcweIKM8OqjbiAh+QchYzLk52a6hMyrSFnKx2bITbx+11Wl/2FJodZ
WuhMDgVPb8l8TN8THatni4xYGTslX/0B+UBVQYXOgq5fIXdU7YwLcQNi18AR3mDL
kDusSEL1pLoj70JzcgtMP0Up99NDruGC097tzdlsNRRmOGXTFOAbpXiWtUtI/LnS
kPaS49JJLVuKvLozAn0cooqx6GcfsEYwoJLuOgNPvRG9NqgXVQhHymjxQuwshuKU
ksbhhDsmA0pP4Jtc1xU7RySVhvZHGjri++wymCP5pCJnCq1zSLO1dYEwgAHmfV34
oBi/y0dxpl+m7JFy/giLJazI5O+nli3sJWf4citBUdgaP+2rbJguXq59+PRk1Avc
AA6WiVoHxqTIOLCl9R56x2xxPvSTPHfO7LemWRdxXt3HPDeqW7cGFJ8wmdqZUTje
zxCZ5LQ6+qQeMYXNQ5BrtjxsTG6OIQY1R42QTFl49+ceFYh8HpRBKOe/UYmFJySH
7nQtA6+3nHm6Dvl+DAhXS1iDWf/rREyH133QK1rPHaW6E5XAXHU81GC4W3yI18FT
M7waOZAqi5Kg8Q4SN92orP4/h4QT8nYTP+ShrYHJArrRLqWaVJzIJttDp1ZKwNKP
cRr8/Rh4AEOc+W4sf6M48WRFkV6C7xNolkA0f535R1//DMzGNsXU3tnymod0m1Lh
9JikQoJd2U9is5NVcbxSe0vyYq1fLHkOJU92iRSDvv3fiDT/wO0d/QCtNc5ILIa7
`protect end_protected