`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
7A96dmSgV4zZrliWlafzzaTDzeFZFv1M7QoxhQ+R5NFQHZTHgmFSxUxpt/91Yg7w
/RBqDvh/nVmDYUsvj0AupN64D/1lTb4PTB4M5bDsHCogPRj79ESWsgcIhpPgikgB
MrD9hW9fu03cahZRLJh2dL3okQnCvtHSIQt3dR35bDfiDQc68pZdKoSvlygTh1CF
zNM0qbTQnuGcIbicUQbl3ljMSHHY+OzaXVaRYbQPI3kL2fQuzxirQVXCflaubxN5
AKq4NT7PXaRlWEE2vw3Q7LJyOeQTT1cjyYOrkV2n+dpv1uZlvImChw8SDj7zCK0V
ykCb7kL6AhBjbI0OQs2iznxBJlTpLiYrSwsrjP7czSUvZbzQL7+0mNo9pH08XQef
UBRwkFg124pDbq/aBW+yYzLmGfyom6QpGv+SCCiSl/SrxUiavyjSxTNirPZeaRNL
Cujpjc9Gqo2/ua1VwJ0NnrdeZuE/52uCNgl3k2qUjWtvwZp7MMF/c4vEU1DcxYXd
ORVrmMRTVbBKb0fn3ymA1vOGUiYJhFlRxeXI9LD6Yt6byexV5m348bVUxhe9nDAm
EI0WHlcTjoYn5IVLOrrzw22MUQ1rcZKcCscXI/u+RaJVsD2UoD5Xl5I0Zt7TfJ3M
nkqyhNPrknFLjJDSZfvDsdt5r4n0hOHMKYBi3CHCfRAqLnuEvcb/zQAHXpTmqx5E
JLi4W/DWChE1PDE97sLtlUrFE6t31wwH9WpIAmVI/itl0nUxdP6EiZR5z2s1lYP2
QDMdpoeaHD+lDRwiYT2p3np4EoiTpkTB7KzePEZ5drbnRm/Lil6cekThpZHglPxO
c1PozkEgR3uiGG9XdcEbFwfD00gVWhQbOQGK26kT4mFWUOBAyrffUTIJLrZL72LE
F2SrzY4g7J2/sPnaKfThVoQq+EPQVua8zJfqgj/GjPZ05RO8eBaJb9KFaUT0OHkE
ncdAgMnv5T6OdU71zXNidfh8K44SQ+N5kB5l6RHSCF+CtPE/MSpzJglv1YrbhXzQ
/uEDA60dOjpUvAaH3HCtM/UUYBRjam6At5GnDwY74b0SY+N/frmEmwRLma4vMz/f
O80EXnEV9N2Q4t9HBHsGoyLSC1a25ANvKvu/18c76UtKP78ca8TZDnAgu+BOaXxL
3jNIoKk7uhOB7isH7YyKjFKbShb/XkLniJLZXzQqJV2bYzdXXXFaYdyfnG+O5qL/
wZOGW/PyeqhhY+Dnyu5II2UKZk4c+3O39BxdElzJ5h/+INSc/sxI0yPdk6HR7fSM
NHqlQkkIzYGK7kgVTJ+iF8n/tJ0s2Xxa5DQU8gaNMlRA8XjdcO1IdvbH92vNKYZf
QrBFF9Xau7ugOESD9Ee24iCwh8typPGyGMAt8j7E9j66EzI7CXnbVvRCh86BBseV
1Cpj/k/soU2ZqLEo2mDedhf7uj+wjqOOkWzTR6k6x2ECs1wnTKzysruJs/95ib3P
Z+LPd5V3Zm+AYfs2e/W0gy+oL3Y4TIXv29531kJVvPqaLVJxDOpjMAawJwLT/gDW
lzSm2ryyAggWr2qLs45U4Isw2bEST8DCNYVkjTMkwVZvsFwM0gkZCujaJpY+QiVX
LZK2ib9UhQu/zpLytlXx2rT3Iog4R4cw7SWOKddQS7p9VKiARxVryKpCcU98p7Yp
0EGv5ZNvnkFdZOwX4I/O0tOo+mOs1avy7/yBVosBtixB4JlpxHRNlGlm7awdQAZZ
6eQQ8fxaMWFmjj+YIVlJzVNygClaIsSOFZrsAIQNGnCaoRffhQI9xcA1JPj2KJpV
K9vR2EfbGDBMnbfiWZP8oqJxC72dndMsmPHxmbPT6z0SJzFYgv/CZSdIPuKtvRA0
NcT2fClCBn+VOQ0a018AwSOBFSFyjWxxPbdkUlxVpEW55uT8LC4o1e3/0O6QmT8H
N2ZtWu9GZj7l9BCxLVa8jaRSi1baeA+uGWKbqgPKsKS9rrEz0vY7BmnjmLJD+Oou
ilyYMSQJDS8E1ZmWzKcaD6SaHbwJLrV3mHP/Tjxf0hnq/g0FQ3wsyhG2nyl9w6ht
1fySp5WVe0m6F2wIY+hZXYfk/F7cha1CZmQP4ZGN/3Wz4OEYKwcVAntvoL3arNxu
Kpuaij5hO+QmEXphCMzqxHBCaqRATqNgPplklYtUlbTZrcE3HzxJ+0EIW3DxEHYg
6Z4VrSbBOwXcEEnEz7Jk+jGdFaHLzQ2P5orT4q8pB0QXIaIscfqMv3gf8lWn6r+l
sTTxoXlxDC7mtqRysnN+KOHwvPd8aRwBKjA9cQjpEYw5w7FAE0L8ulNOuNGsk0f1
LTZWObIYGiyEYzdFzeDC0YHmkMbgaLOy1nvUwo3txqw6pzyhz0yiAAFoulYwkMr3
6um95361YtCS0LUXWqWB/EHA5cPvXra/oKEQekmOGHTBSbr5Dahk/E+wSpMk4tMf
PW+eJRwu+9FqoNPX5ufjT9D2wyryT80gcrm+6+i2A0S70AgSyuwxLUq+Os8EMCSj
KhLQ2u7OR+REP8SfR82m1wg3qqigtUSFX++9Nlt+cV/DfYOjNjjFKGG8a3hLD2rF
ZnxZ4yV0ZwkJU7E9x8BgcL0Vav35OX33Gzo2d0zOXPrJybcTKY6GZkO78TGVHU/Y
9gHWRSq9I1isjJcbJ6OpL4pE+PZLKIqg1igvG5tktlsaOtSndEpVGpQltDvdrkIY
zkAVYpGXggfXadzsLlhgZstBJICUgxjzHWvVdMQB9N1iVPYprNE3I6qhxSVnIzAn
BNR4nAoeTWaHSsV5KQdq0ZHvZJs+aVkly2/Ht7gwuGf5enOWii9fH4xkY3T9iDkA
Mra6+UXszGogg9fwlSqG6mGYK8KSWEMGJ6rsoR3drF8/dMGil97/dqYv+Tny0INs
JtPurUMQPMSn8H48OI7ktncJYt17nuJtPWq3k6bpRMSSbl11WgzudR46/xvRpmX4
Xbjg+ddks5mStE6PzNtSqhakXgZ1oLgeagLej5m/DdAD+IRZTZ0B6N8mrl1Whf8S
6kyNQxFITfeQZIbTGmIwzMJzeM3cDdYqEkdqr0CbUS0OzBlGC+v8ibcmVa2lJR4x
bzG5LQ1fs/bJLq0M0NJKE7MMqsVkzLGP5iimKpPlAqr2WoF/MeN4z9bZGxSWIGk3
ZBLacY66e0WOLYYfiOVPW8aQ0U5K8vjRUW/tTNUEkdwk6G/nwAOfZFJhKi3F6m/k
bZmjZcHyr2QUCJOznEp/wOpnmlM3mF2fKHFbcbPF6bBqHBzQ4XNTWaLJf2alqtRq
WUWwlTOBE5+z5zx0HCf6CvcJNy73aiynNmhg4zylybNZoQen11nSDh6l7/LqrfaL
K7c38vlS6WRJQz3wBV+Hk0GEGEnC64G6Jkwd8iuWKU/FjXmxxHRhMFmZe/mmeeuJ
LhsXJzh1npobvwFwCz0PxZNag9ce9JKEbZaBSpG6CkzzpjlAwIh0npC1aRwggocG
6Iq2+BYgwIOBZl/lJC0so3H2MGrZStozu/DOQ8GBJzG7dVuZB5twmL8jVEA2dwSj
EViJkiHfV71awMJy7YkfgJ2iif47mcO0BkHHnrv4s0fRhXcOdT882I5MneZcwuEl
QHBnH63W8ZhiyljtCHL145CrEUABCQUqHPlxaanMGT34MQnn/rbS5GqXDke+iklz
oYqZacW2EklpouPqGjPhXvJpbvNgwPFDdeFxmje7tS/Z8Yetho/Js5rhxuXvbMkg
j/dwRDibiKNQkRjl5H69GbxK4h+1cCliwdpYZxk2DGV/pw8Rwn9vC00wq8tm0qT8
brOUNJUfqmpEGA20iQhm2dFpTAQ0xhxzAC5gpGIWUW6cp7CTTkhJ1AsSIumBlD9y
tfrdL34XEhG9C4r1LWiRORzEgbBECdVixclJMOM1zYMeAGA1mG4kH/iK8Vw6+oqZ
6+6T+9GWC2oHfClXYO7fkBu7zhj06F+Wbp/ZfzAcW1TeSwObAM6kA6NWILC1vzce
7w4g+AZ7FFrvNSmx0wwmVM+0OhMBcPL3YE576NAM58RefJ3Cb5Lrdam6YK9fpG1x
x/BH3mtzpIvfjU/GQMnEZ6JYhnVvh3C8/E48dx+jPGQwkS5ix931L85W/IIB05ai
ZEZ4pONAbeaMC5ewHFvYLEzEKE1T1ZVKFGvfGCsSYN+6m9Kjspn80F2omSx1ds5J
HO/otcuKUBRtOug82V1gqWKsCqGHpRwYJm/qumrjlOS+luS5Fksno63dRQ85tXjO
txOPHO7JaCeor2cG/S3Y3elAoXL7TfG/hZlbYAO9RmBualyeddYMNkLlUGCBDzew
qBuCXzWbb6OC6dln4N9E88q2nJSQhvYWXz0+TmT1SYT0RugUqbRyJ9Phw4xhCdhy
zO/Yo0iLPaT2IY77p1oMu9UA0ysNfZ0yZMXP+QMM30epuPVoxO2r2WinqDZOOQOp
0XAfV6kG2sViPhQXd+u5YBaG4QJsESZGcFRBC0NryV7miyShJ8HR9KHzlYrxp3y9
X/+Q3hBke/w9385h4qrKO2EmAb6MuzdpsLdbiuYriPSg8lCCtk8HcabqCdc+fTGl
bRiBL8052TYgAInYLuq1t+g2FZrr9ofRG/rngbyY08p/M+Xjx7pEJVGNEvaSHBiU
psrqofVeEws3UV36tBniaFeou2aTNZnlZubejPM/+/VdUStq7muLDdInGjencqzN
hO2sHJKKxWRfM9UW8bd2YALs2HBOJQjnqRQtz81ka6LlbUuXfTUfqPgkGKI/hcod
5yu74F4hDVtnwcvDfFW1BBnwbnNHNau5hBf/vWLnqX22wnWMJ0SR3qm+guFwLtwd
eqNVQzgPSrNpD7dninvme+SsCGc1uxKDLSew/6+a4Wr01MtahOlLF5G0kZ3OKJAl
piJYcHndDOd9yndhYLgnJWPSgFXMQ79s3BBDiNL4LeEs/tMH6g0FR3tbWefjHyEp
HBexpZ8CtndejsLh1TlBrpjQx6IxuZNsqXbxsh5UIg8jLQmJBWn5KibVva1W55Gq
jhboHUQmTEs9vda2imjYidBu30BrrnPBtaQIYTl9QUrgFQFeOoORK3VScYfHIwPg
LNLgZlaz68XIDm4iRFS/FPf3s1DbVX6W/i0QVU0u4IXrEfHCaktuF+vwqNoZ9Tdv
xfLWuWzjPONoSZwOY2x/illjYs0Z304Hsx0RHQ0Nk6s6QNJt/kl7b8ykxVZPmHkh
43T99PHJltRZwNJpPVwHDJCMzsVfTPBkHd/e5w0hiXBxofM/3R9HTAe9+eL9iswH
a4bJ0xH7fWt+gXOZXZp1lHnlsCrh0BE363K0c4t+dqN/yLb36DwUEs34T2442nGH
cjbL3USwq6qcRNKo+ile68FQSiRT/JFI2rBdYQuZu9JKx2HbzfWzJ9pDueePBaJX
YArWcsL6BzvoNCHTAUps/x5oHvTonqm7DTznxdjRjypmZvXJti5XdrCSNnn/Fljh
cRHkEML+kd/UaX9UqaRZOC7ANdyro/0fr2KhE4q1KQ9fxPtWzctnpQpDtEV58qcz
b4zedKPUlrI3jPFSx5FdBOLwH8b3AHvc9QA76vkzd/3Kre2K/7IMYSnn2CbRd80B
NMRbMWY/Otyv8etaQ7jUPFyXj40u3Zk1iMmIM56ofvt69S+zT0L4MNXk+DQ5bRJI
6nqd/T7z86RVWTlfzNAoxzsFSB/D3uo4s1MgqK2yR4lB2LNunTU3mZ7U3rcbHKrX
fWynRu+Kk5TjQd+T/mYfGrEhTHnioGKQ0lFq6zV/g7z23Z3La1MgIm52kxgYm8jS
jC6sJ1aFQJkvfMpiZi7lycxux3wcb587ZWbJhnv03ZpnBLsaKypsu2Vo2GbzXBLt
wxxGGaklYpECSkUklk+qvcxKx+vGZKHdOjs3pbkfxoAASwiRaGsPGhGE4PnEa8c0
CzSO1C2GRP5tIpwv+3B1W6EF8ITrAubGaawnwdLYOpR9biduznyXdYhG6EM3X276
rn2CSGraEdwTWGHxeebcyT/GdvNroCD41hm0iEbctYjW5i7l5RXT33M6RxMCCvh1
1eAdltQkZIM7Z0vVOsJtRbNfbkjFK31436r2zWp+Io4X1ZMDnDn8PoMG58xsSNJR
fog9YRKTrMnasmx8iF6AArj3vbhcyb2ENKLI40jfS6AD+RiOnKrhY0P0tG6Z5b7X
m4eNuz/ojg7A0wuYvYG6L8VhEUiy3x+ETZX74fstq8sWSaa/Trp/jETh81huD3VS
7IMvirO86zgJM9EhA706gxe8JBW+B9S4cOS3SOphmDOPAq7jtb0qxje/VkFpsukf
zoq71jpAif/apBTG1+G4kdI5+eLInFptW0geg3jRh9c3AScUw747h8bENH8dI/UJ
jzN8ppp0GclBrx8sBXZpqiSae2Ry/LFqi831xZAim90bZkMAQ6pDYgxvu/fToyf/
gnfIkDtuV9SIE48AeGdHLeZxacvKPYNFTEnuG6RsShASFikoWiVLs76NyWrkD9HX
6cUouu+6ejS+jVFmp3e6NElSGYeRCgUZWdtchhQEB0AzBeTCr3tCRLOLeiU3H/pK
OBLRPZ9M8R82pyErTUlQOm1uA9aThRMtzuGMpu98cVaf8+tJkk9ifVydpo837OXN
X/pNeN4xjho1RUizKjkN0fBfwbK0Y6ljVGRK0CxNL89No0mJhYPH0gOliwsi9ZGs
pxCqx0EyPp3S3aVEUXZMJWrd3MW6VYyEbUJhxn2XNqc8baNIVn1WKfGAiukn3D/W
D189NJVZRMFF91aECY1TgJD2g1UkKY30+p9twE+RyB3iyFuVCM8g6cUTaDQGPFkp
cM2uITGthrZmNssjTyGrwd5PEuQUXuJLuDMWKXiqNL7lbjbVfT4S4BI3et5x5BRZ
QT0iUXxDtcj1Ogd06VjfLcDbcbAilQ3AVm9/h2zFJdAlVGW1TJHKWBraurecJEtR
tWPDpiwbmh3UA6iTeCI8oHHzeMip8T2JAAK7dOwvMtFKjMIpnPjJPO5lour5ZHav
kd8dhRpbU/fcO4wKUq6vpR4O9p/K++y4PpSPcfwugID5usGnOW4w607KJ6X0UkuJ
nRF+kHmLcdxl0zbtZz5KfBbalwjVSJYWjTfGjkq1+HUh63f0k5r4Si9FRSGU7wXP
YlwYl/uhWs4sTKwM2/W/G589V/aWWK32/kJuzdO1Fs3NgajyqK8TyyRj8+umJZnx
yS7mSsNvhZGvZKRMp8ozKSfH7Aju//i3Ke8efK9dlwjkl5fy/dqVKUfYwyE2hbGu
lrDymrh9nNBFiXWYVCgpISkq9Zm9D5kacr4hS4+yx4KPU78pqRZlm+s/qnso1sFj
SORRwMSPpg/ON4xnJS/lqJEY8ABiYQGizlYC3jIHxScHMBINFQEgA6XgRuFD5x1r
yukHCDZGORsKF2JR347hB0TYMdfg++6CKUQK14M8DwxSy85MUR5pb+RTkk0gWHkb
//+mfIxYyqK4yKr8VJN5aYtYdpSgQH1P2zuyeNOnN0MVx86Z44gSuAXpO8jUixyA
u2drzJccqBs31AHpDvZjkxDWUkanaBRggE/yCRYfBZ8tf7lzSTs05U52gktj+TyP
kNwRdZxAWMAFndjctIJzj2GZ9WhJ7HFlktB+tXEaRj7svJMJO45/Sdj3IhG0ilHT
U+o7dU9pguP67Th3r25rI2zhUQncSm3X4QWofYzFb3wAyAjzNWXFedlUfmcOcU6r
q815wqz+DPPGp7h3wJoUpJBPMM3SGAkGQPP/NAsiaM0AHD0iDXMcualiMR70nEGC
qWYQ+Ildwsx0sNJZmjFZMhOnNQTGzOjpkweKiwAM+T5kkNMuVcOB1k2pMzxdxIYh
kD6wizlY1Hjm+1RB0VJ9FfkIQLg1V7lH5V+/OlFIesBwBjdOEN5g3LlDe4rIELl3
aErD9+dXJqYUE6hkJ5GI+78H7HIvxXCqhUyt6Njf2GNOOY404kio/nh82PhrEi+Q
+V6ImIQ/5A6bki9CK3XhGKF5/gVisVsWZuCaCt2gBWBkMzCAcdKfqZwhC7FVHgWJ
v7+zJdHxxhiADwnbDerz66vKi+1F2LECG3gBqj/aEX3cr8FfrBZkYnpZSmRrtmgn
vbOtpDw4ibh6VF4H1yVbUabPpFVeatve/a9R9C9Os/uFqaoeGcfgGjNEcMdOebPW
kLrbY/JHCyxfDf0V/CsYaSZVh+A8WEJOiVS+NhFbmihfJqvxYyx2h1GtNllWDNV8
aCUzrHpw99gLJB15RKc46+QmRqvgswoWWQ1v8DW00uWywRGKht6ROv7h6RBq3skb
ofoYg4EyKM7JH0xFjbXBDeyeK0hYRh+XB58DakuPAdUZOPk+3tIrY9AP8XFenNLQ
iuZV9+aMeyJot/9N8E3M3/xLOwYDAhUP0slpLL5GzmL2ka4v+e0FSQzBzOVX22ao
hi0elZ7icYZX311WK/3OcjCCpdpCAd+YqZFjcHv3n8wmkhzZS8o4MEHXLa7fUwwb
dGQJgi8Zhj/q+AWpOTvS6Q1y4YZsGphud4HvfLKPxUTLrHiEZIa3wH18dETDxIkD
dKANp/GsKdz3TVm1oyd1vwN/1BJriDivEMkRDXz1P/ugrhl1Ha7gS26xF2VbIRCS
5HyYhjUcj0s/+YSUKCrzv3fVPpfrQ3hG7jeOMgLMfoPNbhsc5aWBDV5CNKsHP6pU
Ov++nlMoOXEmL5f7DEW1+V4gBh/01Gfty6VnK4TSemjYGILSI1D+aVD4ZvbO9kt6
PmbgF//ty/ufTC6Y1W9dIB/Eb/AD1z87AA8hJugGtcDP5LVc5eK8VQHViTXz1LPa
Y8mp7a+dql+ptFAqqDqMSJF3lW9DVnYgJ2ByWgI5gzGWHYUQaKzWPsU/E+fnNSeQ
9k5nZFuKLlgdRqi/a+KGxyZS0+JkZKZ8m5Xwl8KRJ2ZB2qmZFlBCCwowZgu01Ulu
icGUxdjvsx5XaKsDLi9Yksr8sD7/JvIcjv4KLKfWFFebe+hjPiOtH0Ubd/O7NhPL
i96s0daFA6n/CMDssKQokPP3jQgQs3lJScq9n8onw7Y=
`protect end_protected