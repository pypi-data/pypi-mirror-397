`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH7L1XaajYgXpVXTbYSRXTaYLp8fuWX3O1Qow6GgetLV4
Y5t4mcgSyZqWVqOz2JJU4dim5v80Ksgw6ZBPPGTihbKORTdagdU+CFEHVssk1NwS
CM8Gqa7mg/20pMwWnJl7TnjPcCIfr/WiY1Dld/VGRVY52NWL7HYUrjigVW+zlkQN
RU4ygonyzoo30t2kdOVI3m88NZPkYDaDBjg+m/e2RXoN9CNAqpRsUQ8AAEe0eYee
MsXfgRSQuCerk1RB0B2599eV0fRITOLbnMNKTZ4k64znfpU8jGwgB4qBbLq/TrME
Uq3X/KihoLzjn5wVLdq9AH+eQEvpuP/F/peEHny6UhgFmpxlQOuLlppWTXbXeF2x
p7PKTgLU6Wi51syMPOgcLguuOIAF4YRImAdgmQaGpSAsX7b3PnGIoyIZg85apMF8
/D+L/D61cKPSrFqdTqBV0ZzCVlRHug2E9fmcKTdOVAgTs/w1N2N7fSqRbogY+pKK
L0CT6+BVlySAe9Vjhx6tCOxldyayQiW9QMfKAEf6I6aGsW8n+QPbT89HJnmnnQAf
GJlSwB0Ex49M1jbNSRCX4NeKXBSiQOK2pHPfWwhdzc4CoWgXJNGSy+KAaeRPS7Yt
xrglPs0m8WLitcT4WHw+Wi9KtHXXXGcvrO/wphmpDPDZu/zYK1wXL9TQ/IUdpcbV
44Rm5wY5KWodBpfnJJwFmsWIekogOukwewUkbQUlN50AflYMfe0t456Z3k3BG675
pcxRtB8MoA8oOd2tb6x/oDICLJnx2magF3fpp2NckiSZaYwxvGHY9wtJ1xXuZwnd
XOTahCI5GmpZ019rlUhQu9taTMdRrx+m5KlGjWNdh1hXbJlzPyXJhyO1ldYL2vss
9VN0Ukdln72SqaOfKdnyXuZM8O42CHTMOswZkYBPmo7JIN/eOKqjWmShIWxmAvNw
Y7Kg9BdGtFg/QCzzcD71C6iXQoDwVjJ3BpMyzK64SGka3quNqHH7eOwzWmk9dj0a
Fohj/wIVq2BoJL2U3BCvmshHty/Sl1YI6qsH9woxRhKfAMNy499HfvXQ8m4X/r6w
nAKypn1JAEoR0PxBWOBzMXpQvk/OkZgZXJdhugvWKacf1z0/xslNTwGJQWGWbm2b
N2n4kUdaYQnT6V4U2LO2Zl4jBiGLUB8hJKfv66w5TvsOKzzj9NzeA2/ucAVfEHjg
c3qkLY0lR7ACOHHJRAJWOzry4MZuAULyD0q06ffd3jJ029X7nSIIumiITcSppHNl
BoRw+cEVlyQ/pO5CKYE6Ca/6l0+9DTF76NE2KRmevrbd7YTv+hy9lVfd5AlQ8vHS
E/uoOR2pBIzlxlKlxdbs9J331dOOjXmWigOB99PYgEW3ZwpKUgvAQVk15lIPks+H
0yS9a0/G4dkJUfYbMKYZWok6p1++on4GHzm3mwNnD75HmxmnR4t6Eq6EbDwK6bhv
Y1ocxhX/oPhcB5u5KEcAJ6JwOTzPavzmlzwhFcsiUHso9mQecwNgq7hGUYtUBpi7
BTIv2NHpW1+a8XGUsteYrSzp33aX0qeVuP7M0ccijFnir/nIP6PlB0j35rxuSTiP
0B6lZRUrKMuMHkXSweI9WhvNGkYMvMT/xzsN8n6ZPOD81etS4V8s3ddCnt7EVLel
e9QDMY7pr906HBPb9zetdrptFgx+QIraiR/d+wTAqTGPrxRxR3xN3g4rhH+cKBUN
cQG+MDLokhVvvRm9gmH3CW3qRLgR7TNVbT8W0unlgQO4lG2GYexoHqvUHlERf8G/
sOeo3C2Ejg2GzB+Ilxz6XxcgqkwPF7mxaY7PXejUWY5TNvvoXGp8jTguxwXnDLVB
qiVuDHiRhWjThbwJJ4DjIpsiqJrj6SqAPTQNSPUBsuGES2F8Qpa+Z+eNGrtnIC1Y
AvozXgaXSU3nvTxqLeAk+TfmN+gnGQ0fNQhykbA9cuZi8DnFizM4kdd2OGhwmZ8B
sqSRiGLk+G0jEC7rzlnnZt/D/Qb/W+paTqRfXUgaXcDHntf1Q1R5kzvwpUGeqEI2
Ffqm07ZlfOjUAJMgnbnIA1HufdsPyHriE9FvhAjkaMqfHH1lvmZkMR52eQrPfJMG
0MeUdfnixK5KY6gzZEDzvE/3/PcFqecgKkbJ5xBKbVwuXma88sgeTbUEbRD0x7vk
oSfWfmc0OITdI9+aEuc7WJWOLhnsL9WWYyqE537jsFblh1UHRMz+9ixicEayFopu
vwuI+M8puYI9d+yqyXPNzZVVFKCiFIMrS90bXSjbZ0yZSkD961zLdW2t3RDbWT+9
iakFJnakaKjOPgJVGq7T5Z6bpf/jHfGjYSrTTTKpahA9N2VQns0b00JYm63o9QhT
PtoPNXmmM+4LTn2hXjzpu8htF60MM5gHFEkE+5mZzVwvbJFm2OemBwJfEWEHXhdd
QJ28CLZrikcmUdcdWficVwExRv8+tEKDUE+mcP2+QRFtQG/YcI5SjI1Xno9vNlyT
9AKF75NgI3SlWRKlbHS2VwlkI42oCyv8qSICBG29COlSZJQVhOdiG10ia5h4nWQD
LSrwxBhIetOvzB09B+fx7aHdRo/ofZp5kibnJm8sOnOON+/Boh2Yh+JquNXmq01t
eq9CttSZxQKieM4wOWqcgUguNHk2tGyzWFa9aqBrNjWF66D0ZagLEOL3AhsJkzM9
5JwRXG8Ic94fqCuhwdjLBGLiequiwNf/CsCvOuwjA2lifIxslQ8SGIXRBMcvUz/0
MDd9VwX83V6KEExoUR0eDNsmfrXJIR7a0w3lsa0mJB0JCH7ecwPfNhBBRIfR61Z0
ZXnsOo76laiDilVVfvcBHx7ksnrKfsIuCuV1pj+UXqH3TB/Ek6wBo1E/aT8X5XCB
mGUm17gJwRF3r3SC58BMx3MTUKMgSxBLVVmDtmNhOq90MzhbAkkMPZU6cyt7OHqB
ufHm9woioSIkQ3FKgMboyDrQUYP5XGA4xd6HH+ohyTEMc0uWJZ463j2tXJnGQO2i
SWWWJSw8c3BYvE0wSF/QU0dMRE96dQXJgInJCr1wknUaRcVCyZaOfafLnM9iauVV
B11uh0t7jr2I96WCbwIJUoqg09Lnyeaa5UCdWwLLE1Q5B3NsZtYbQJrQcOn13rIk
iYaWp4QKtNOvJlEcrunUiyj/Wm1Y6hU8zLW8GsoKYLnQruBA1kdBa2njUDuAFiTy
GQklebY44rd3/AcY3tX3dg45QfdRQanuROJ0S5UU1jq2bKxIKvlizPBDHhXzRsCV
HKzqrLfwi0+X/V6qVqr8eQTThZGYBCSCRYDuoAYTu/+hM8ELWnVHxBRy4bTzehz6
rOZ/Ief7ZHjcku/xRghA86uK3CPveFqykySgpEBEWM2vZVBSpjCh1AiI0h6+Fvzn
UmbHhOMd0LQkk6/eVh8tJW61Ikc4xiGVIQOyDT8W/WNg1DqFFWjW0reebL4IyoRC
wTs1WzNGf05L9ZLpgVXYnlqzwtZZru5oluMZz5Ol8lzX9eLmJbDLWRZu78KObf17
U5ip/nReg47qRtDURWTlbJ/j1ZpcRygvx3oWqTSXVqD5RmN+S2Xy6QFZQ00iFt4b
+InUcIei4VXto6cF+D4A2hPxUQiPvRu5gdwDVnRVEp1iycsRDb9ssW3pDMghG9iX
OvV6g6g0pej/7ArizqjTwcN7aO3SjgRaxpfj7N2HGDGG/V2yIbeAzii1hyW+0P/R
Ytgk5yiuRIBl+3Fw0DPVR7fSddJNx6dlrUtTkl0vshZZvdybrrLsOVn6EDBgZkSs
wFsVbdNLox/PERUJS8BJftpEX5ClFkow3FB6wwkIt0n/s3HtzviWr8bak6BO7Bl6
HtaVpJinZyMhijQi4OicsZmbBvg+WthZF+Ia0lLtKRozIlY8tu/murLt4rwdrtsW
FJA+cUBYyH2Y+fnQjyOO+QUkSHP1gxpDypkIx+K5wpeHY0bqAsE7b7R0TD+lY5+B
76gONGIK3LILplJ/o2uCP6ca5Fu6AlTxhTs87MB2nkAbleASJ2EyHRqgegGTvIwh
a8geEguDhmmKbo3ypVwB9ibQQoavF4lA02jrdTk040+BtU0Js6xL1+YpzKlwKylD
P/+X3GUTcxMFhVvuTfwTbA40Gzky4QkD79z/GUG/RbZWA54Gn26VsB7ycWBhjn02
95jTz6Xr8OTsgKs89MVSUWvJ5299JxfAnotk7CBZvfuQEHgQPoUz9u/hRUrl4msh
l4ytgUX5KMopVr3s7KvuvgeQC7eU+P/4FdeLgbKdLbdci2BZBve2O1gqkudZxxiq
PgVg3zlq/y+8uDGoTOTO8LT2XPmCWkTv3gr0ntFai60U3mGR59E1cMWL1XRhnhu4
gnS6E1gF8QFRoAuHbhEU3I+ojuSPzd4j4RCR71/t8sVFi5i+Y8CrfeXkx9Uso0BE
1xAlhwvUoP161SsshgT5T6gmwSnRSSjV/ychES6EU9gG0+jdO1woTtq9sYDDA3hM
rdRbsvAiN3S2QAGXusRnDUiL+uCVZhiyoxVu+B2ifsFMtS9FnmrgHU4sGEO5TBHz
5FWwG1vmycP/9R0VcNXOucYsSArgLWpK/bfUsNZvjoyo7RlfmTpzyfGE/E5H0A5z
jP82i7W6R9FBeSXF+KJl+uWzPZ81j+1uhr9ve/Zs9g/4wUIj/zzqogSmqfyFQG1u
KVAueL3U929bEf3X3movBv6+IkbElL4JXV5Fhl+QEBmjgkBzPmfOFd4oeeexBqSw
+ojR2gke0qEMGe6uw7vjNcnZ2VT9o+6IhxERQUvQumhukru0NwAazadKSb2Cf2wO
KXgZvRnkH9FadugapYOno5NHr3uWC+HRviZuh3l174OiLg0uqILthugFp49T/G3D
mUyWplydrvdO91SII0hmCpwJFAjNkXfPu/FoqGOlhTk67t40H+cfMEHCYxci+gyI
NX+HmuHBuSrM96vQVKvWUxHJlYr7ewD+/5+q8aJwpaihPDAaSK/0Xc5WbTYVd0K7
1w1IQ4BOHaoRGKjS50/25kTdT5voVHmMZHXNI/M6zviYUG/y7p4vch8hP2ape6P0
dK610GloYS5O7qqnY/qwBQb0PiDQxBDFbbjzRdyrnHapTEugvx7k9SWDSLJOfuxi
O425eZvb4HnoKboS26Z/aVf5ziYyl9q9t5V7vh2JNJVbt/yRKP/8uRLow6kBIiYR
XamxpV6ugmj85bNuVZ1nWsEQ/+QwMF6gWmciQMJm8bxQYiHoCdUEvdWMog+vDTVb
dxHL1SazphN0kJOntyv1u38eM7ctELu/CdPh1FMxRlP3wS+S3UMiTulaSrwnTLYY
my0+aOg++Zr6nPhiDQOUd4ZqDlIDgklHR/RGZoubDOgoSzjShHOE6WsRIIaQLdCU
kENmO9EUwOw53bJnl30v/7u1CetvRkZqs+0emtP7oSjnDR2zin0qDxlXd7/3Ia7d
yNusAAXrJU4BQkGy0mLodE/DpKYK5n9GyyDbs4McnGVPe+r5KHJ3GJh+PuVx7xjC
oFrDQtlDpv1/K25/GTZu2elgUhGcAh7pU72zyXYfaWKVlrwQGQb5SC39l1jqTYGM
gD+XwdxF0vONM9ac1ZaW72JbqCIcr+dtXNorgbc8EO4hcVb5vf9ThMXBX1E+pB7c
6FradKmxJShwdcuI19ZWwH6wwfuCqOSs0GsHWR9nyY+wk2S9738SNjXYU8DZpKe/
4ll135tXjrHl79nw5ta2v7yjZMr01B7jBM/kSM3GjCy4vvvKZmQnuNKerJGmFoA6
N5RhT75nQw/Zyi8PvAAWtFONw07vHh1lu9C1t86k2PSr7SoW+FgHVTZt1T1oRY60
HxfgvLxDaDenWQ1W/D+6mYXGO9UF1cgJx80XsFBolUtHVGSX/0gJImXOGRlzKqH2
q2ZVfF6wISYfWGj1Rg6m9i4SHiCLdMkJgFVVTJqOHEvtggxAyh87KhyZsaWvo2ej
2To9w7MdUQ2LbJazkwu7lA/IpYbAKvI45uROvXc6GPLjsu8cNJd4i2s+M23Mpy4h
izYBk0ykBaYrSrl3IEMor7VDZcIXZSPy+dBS7QyT/Gix3jBHH6uIEhVK24LEjboW
rOktYStnEjvDgqFz4qfuU1uqO9z4y7utwbrveavb6VU3tZtcdY66FG1GjeoURdGY
Ihmdrc0qRd9uYTtW5YtAwbP3u/6Kk0oSjLqtdI2FOqfB0dWZSQ+L8yOaZ1/JbddI
jqx7CSMkOJ6AUznTBeWwrjfidMMosSKIsrstE5Ml3xr/gLX/arNdx1ns6HlY4tVp
6WW1t9bqPDpgA4TeMd1Th03iUZn0M3QkeaCmPntZ/6CJv8/G969x8g+Frk03m/ix
SYfTiElRWB98FeNsTsINJykCOeNDXKw87Qjf087Qm8UdVLdSdx9GHvmqDGmHUMT2
sLJiHLRKmA9OdEhmiSvwRIqIJD/5XZZUam+RQRwxdbIZ2JY7K3sT+64uRO+f0d7i
blMGVi0LFl6S2m3+ci8vdg+dU6EALWvjf29CmZUD1aoeKdebFZp1wdr5yeWw8G5J
w9mGnm/JjY9WlNoz3iyfwU9fhST4TuFGNAu8Devw+dMjs8JJMRqza1XzTzVJi7a2
t4D+gMPb62vQOdxkZOp3KN204r2jBYCbsC0412V4p1Yp4pZtWhVVCcGq8MZQGeZd
CwVN9ibU3kU7Mjj8rkOHwUhlLHWUPBcfQJW4KTZCjnYlg8FWBBOLtKM/x1rpPZCd
RUiqlGyjGcoPgHvUBziQfxDhDj8nll1Xy4rNvRgvuJbKTiYWwwyGhXIoAlSD7IuO
Y0zMpGzJZStmKq4i1P5Q7u2qGMsiPRtY3aURiwrZPT7m9ecd7eLIwkhbQV9eZ25n
o6iZgfu9Frn1OrwwxpA0JGN6KfwarK7TYVnVgVBpWlrsg1oU7AY0z5N2XLYtwEjC
K1rPqoSf/cGBfO9ETV4eAML2yg2jjixPQGdyQ76oCVg51913BKqVFnZfn+AagxmK
e1KJjjuxmiFX3V+KhUqCkqCVGPEOQLzkVGGlw95rtQz4xspQAWsOw52eLKddul+x
AqeHVgEYZgliw9yKQeJM6F3lVpGEvjwdn2ldfS1qsnvDgJvltEAWHn4UkDgCVK52
N+5pN8xv4ps0UdIzs3fIiqivjl+T3POY5+S2bpYeudlyorYYTZj8COHf7lK+/ngE
UldKg63DTFXqdJCk6kTdAsHJk5hQyUIkIwr8YmfkNHPuzGyjujUFwE3ZIK2u0lrP
CWm5XTl9+k2ead688WVf9V6tUcdpGfdWVz7MB5612vNobMJdJaORRR2rNqlU2wjv
q0raVLN5hgIWWsftK2GGFJa0fyge2sJZYCL7nKtKEmyZ0jzmU9om9FA20l7NsBkO
usRhCdZodZCbcshwPcU1bmsc8H/YY4GEByNHvrfonnVLi8RFdL+UbQjFUE8ewHn1
6ypUdSJ+stA/vlbxxvWAoVL+H+iLjth/aMzAqcrKCDBosYRkWTNJbLgAg/ySKMXN
AJ9Os1hGyuqpEUmpoCEk87cc88rg7pt2EgEA+lSLPnE=
`protect end_protected