`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOHyGRRDN0qFmB+KtrwkHg1FP8OV+u9sBvdYzWnFhDedFe
/eHCnfmM8DPMw8GJRWw6xvIESOY0NTetZhw3QrLWXNFCiQFXHI+h3G+I6tOjahP6
5StNFh9bRgRHSFJqT14vSoOr3lwMoAcEIfOUmBB3himJBNUAN/JKCpImp2lj0jSf
YfR3qIagpyLIkmtyQ21o4Bb8TskYByReT1KnL6n7KaT2yTljZ6BnMin7X6iN494r
3RC/dXW8sFzo78LMe3irt2e4ZYMR6MK1biNMNyehwG9ZrJjRw+0EMCMEC8egfIcC
tdo40Vrf5CIpIgTLQLtQQb0RJ35jO5hIxzZntXYoj5/cSitFA4Hes1tgRefk0ub2
yMdSDMT3wbIfdePXbleaSbsmLXinE4Vdj2j8AFMH7c+eaLLtOoDXGJ72xZ7Teeku
Cj/wzc6R0XUDOC3X42JwcOe6123XwstaUI1mXkwIKbPvCwcMLEXUjroGN/sV0XUS
SQ6S7LvFYJZItZk4ABpRLOraPbQK2s8V8i3ri6a3lgeHJQyfHr0CJGOAjLUT4Gmi
8fDeJjqL2CbqSJhBeklrXc6y0uZQNci3GURIDQB35ow53o9mTFYtdTEJP7VZgvOc
8BFJ/27mv+8O+m6POE0wynWmVFrT4eX2V5t0aPz+tcN/Jr/wFhlNAfyvs719TjBm
pKjKzcFMalsDW0Garpk0QVNqt2o91lAM51+wVWaUSkL8loIhLqcLHo45zuSj+nI8
oo3+fb+kGjjOzZXEzYq3Hx1ymwPiV1qD+3eQZwJ1HgKYDCSS3NASwYbkHvG6MjCA
AwHfFTWNhbGa1LmpKfdDfbnjMEakwXFwZRtjSiG/s9uMDerC1feswKNSz6idd04w
5EvPudaGX01MfdL7opG/dNOekwhZpNt7aZHQUq2GXrAZ21V/32sg9Wd8H5t+Mg/E
8dDQ5ZUnWgaFnan5HOIIGgVqSXuKjvEOCs7BBXrk4Gb8MLLTKHK9ALEsw56++40b
5dDhhXtLhv67TqcO1uuHiEM7sjGW+Dern5lfS1pqBQp683sCc2+Q2IbtsTgpj27e
RDTBn8u7gVoY4dmouCGa7foCUW2rcNbIGcQluoOnW4FwKFQeCduhYndh5kdkIm0g
+BVAnWNXShe7hQlokGjm5WmGueVl5MnMiJ52XharRP3nGiGmc9YuiSK3ALtSkWVB
CfFcxFAVwE9ONp3BJAbkP6Qf6bzamv5f6klTYHV3TY/p7+Ifkn5VQvZwDdpz04Mg
tHfyQvPbNB5mY64HNuwLBsoiFq+tvlbtCp1TSYLSTgXu9t92CygPYXwBPHLs+m+W
I0ma5rb7cES3ZodCUjEXmPlX26M+zyFSzzyA4E6aoz9W+Cjhg4Sh0yyKcz1xwS1V
Qzjk/YY5ECBGW+IlWasrrz6hQH0VYKqWKKVMcINDxKCtA3SAm/4HgapaxMd/aW5L
WDoqDw16zttZVIwLFe/yDqLztHv/V6wDQWY9MDfRHDjEvy/EYnEmyUbL78/uObby
Ofx8HRzSHQ3CHNifkaUqJclH4TOzbV/eEZBDkOOAfxbrc39WjSCdz6cFIrnB9S0e
zh5cfrdD5x+9k02xAHWaS7DE//lyDZkqAj0dN+NH0+MCLurnKJ2SnXL8M5Wy2mk8
OjWWdk6biYX5MGxWhbyaLesN8zmN76oslxK3bkg8PHaBK3K0q5fW0g6fu8hZccH5
RQqstD75aKIkqE15//Jeys7eRsGl+FOJNCJjHbmXLpE8IH+IgPVyFbG73+O6ylQH
M559Eg15gyf7DF/1c0KhxcPYjVn0alneTfrSJN9LOCJKUf8Sanx/nxkHICZaDdSe
MCdO65VL4XsCsoIXdVN2RhKsfCTAx+d5mRFzF3NiSNPdaZPnntf7e11l0ndOzTB4
TDGKdHIZ7UAR9udpfByb6gbmcpM1Ulzss0Zr1Lhuv/PyHm3ryNITsxlkWm3LQCjD
WChcwCVRpubz38eoyFJCqS8lbJc7QfSCjcuTkrCEZOTpMLL+NXmdaDQIGkGKKOdw
V7j18jXmh8itICKgonDM1GBiz5hxwyMxYEpjrOkHPivoVr4As9qOr/qncg4Bf6F8
x1LoOqbTVxEQ329QCm0N+nu50nEzNM9cEHqnIolxDNq/qEDzg2XhUgLsUjDFm8ib
D8Z8WWta5V0wGL5vszG93GJoJsNPp083KeVRONitjnj5i7pm0CZcIk2ZBJubn/UX
JQjstC9p/sUee3ktjQmXZm2MRQ2Yxd7pPA932Bxn9TJRF3JhllU1qvEY7tKc/SSj
2yakmxQ6ZoyLFFckQhVOvrLzrtJ3nZLyktdCaZEQJUbHvZ05EF0p3xfxSgwyKgu7
1VCIfje/wkzE7ATDKtdC00dgF+M3JiFmlJByRH8li+HsmmqRhqESdOO1Kwr8A+UP
7IrGdtWYfQHYrWikhfVaqAABgCr62pkAPxbYORjGTvZyxcH03OJnQVkPe+MNpL5Q
BZ7WGqWKGZa2FtjrZ6vW7wjDGlbrJbsr+r+7pfFFdXVzUS0C5w/skKlolUsXjZPs
okRpLI94udyZxUWxyViQ1e+u0RpxiNQy5ZOhTznUZuR96F76b/jbrm/jl5S34MIZ
3qv35Ch1D3J6RlDNtEGHLtK+/G9bO9jF28lqaqHfrKvP6omlIqyKjd2G9S+8Y8th
mCeQ0qqKsKQS9B5q3tBl70u/xluwYyZNfndE0aZ5tIcZ8wi6+IHE2RqYVKgfNHMg
8QreSzDFgePXTZ+rI2Wsxxcl7HQPAsZb9dT1nvfXylkizMgWBkDo1WDI/M4rPvnB
dCym8RTtvuB1zG76WkqotHg7YxUDESI36HKnmMP1UPdkTWdCfe783cZcP8l22C/D
e2LFmyjb0KTj5UEf1NC1hTW19Esa0rdk1RDtQ2EpmNNVkOjksGyCtGqo+tXK8eiI
/5ztZaNVs71xv9JG9E2+gD5NIAFs/A9aQDeWUnnmA2XsCauqtEFD13zc3qQ96HBo
5a8k4u6V2P6Mg+IYbNMOmwDK/Zkj2CfF/IjqHeOd6qGz8BEkBM9y0sHcZzgtPzBl
OpgJb+wjzlYtBECQLFKx3JuWsdGPbu7o4PsesvkzB2zU5OCn8tE4Z0SYzxjjyLqg
kQ/5HoX3I5bSwaswLm1VDESVS4loFFoo24CPUxNYMi9SXBbO/mvanjiNTf5IJCr1
FyROMcZMuJUupzYgeUDaLoKv1wQz86xiDPtH572kWanz+1IzWHbjv4kCayLQnNnq
hC2cWrO0eCKnA4BHgzk0pN2yx+RPCVsxrgCE1OkE7VqGv93ZG6o8EuqOvXbbrsKh
zMau+8UkzRw+2PsQF1qdF8ISQKm1qpaX6X9U1ilUM1G451BBErrcO9JdiFGxF+yd
GfKT7AA6xZtH16J/D92EIFD6/AW0ygs1a2/FcB99V5+P6uSVaQ3BZIZigX9nVMz7
OP8+oQyZiM1YIQTwpvXP2c1oWt/0ZO7GVtHtLZ/qTaVMIuu6I4r89Pk7H7JOVYgo
tdQvkawsdViMIEb5gZgBvwbXC03HJl/KTRMuCpJYSjfRHe8LUxZAhadGUE4URAI1
XIMBNBjAWZng6dzdNHb5rsq43mkcOIo+UiAG6LGglrCyqxNcbI/QK78BSWDEvU74
K95DdQtWPaStJ98Diku37p7VhV1G5buApVDdOhALKx4KomAqyX/sg17J4sEubJzx
Itk9vwLXfbH7MhA9JebynwAJ76t3qrnpZliY+C5DFzwctiT1bikAbZvUd5Dwa5bI
C9wOEgjdz2kiT8FKEuSUGOAYYUisbSG0v27wxTzNf3Phink0gpQmKw3Ri6x3IybF
HJQyUE/okhm7hrxhSAr+WrKHHWHu4SRwBxd4TLZztQwXBOq6I7hq4i/auvKZh01+
TNjBifs6VJ728tvyIEMAaXcjWscp07zhznqIj5iySafLM2cE4yxoJG26uQS32dIb
64KdYO0B1EMlcLA3L1K4s0CN6O9l7d9xNGWtMMZ5ngecr32On+zmmmpKuZm7UtVO
kmlQ35i/qcDjRxLG++6TN1Pm/B+O99f4iI5FHUgS2j62ZY/FIliNE4ZI5VGFV0z+
Awzku9WXGYJZ21pADC6cypxreYlOX7j7z3b1ewF9MIV52dI/7Fvb3lcqRIRp11H8
5ZYCKr4Hqt23vA7II1CsQnZAcDCKeumT5x6jx2J0uCiQ3eHEFUvL315cPivR/pSC
BDhTwM8f4BZAlwHObRRM5+UCuDqJ3pQCEgpep5wemQ4IC9GHlE8T52slEgq8n4dZ
Hz6kHTnb7ul/7VmhJWQ9D/eamT9RYXhhVlCrYD1P8oj3152c2Rhdu0IPWeHs61PA
BBf1TaK39J+ymRZLtQ0Yr4wOMU2m9fvHYFUvFMh+5I6KgsA9c1TA62/ta6Wri9se
ejP1lB/F0xSdSd9r8mDEMCtF9MwVIvbP0fqufSA5MHVzNUIxz52/P58FJ99MXC8f
z1uYV5y7aXh+FybGWM6lR/KQ3zxoadiXhOiSwYdVJoGYZy7l/BeTpa2EI8PmPCLB
OnLMB5QcnTq55qjsBGt543xzFKFk6StVM2gnJmw55ssV/WvMTfPO+7IuBkr7YFx0
/Gqqo5MPurLdssZeNt08P+l44jmlz4zE3dBiLZytI/H98aK0kOjbUlUVlDD3bT7q
xd7hWOKVdZsEbTy8duHxMTFyLODNSM6MwJ6eycmZNLgncv9EM/dLtu2l/UaMWdat
NCr0y/QoDkxF7cEzK/VKCEDr997RZrPhAnmn2siHzhwkdCrdhECPD398ZAgJvsh/
UcA3EapPg0F1UbhPlYF2oeccJG8jPiWPuhsAaSBKc/dDXhE8ehBJF2PRfoOcyjpZ
ANKJNiZwwCIkzt9GwXDWj3TTr6z5/vTh9XKQ3DhtjeYbu8piceTy/byFcFtpJLYf
sNoRfKVIfb9zw7pOMiIaPt8OCKzdWmY8ZJunzkQglA09HWr9THA6jjUA4VtlEF/l
S8AgteysxvPDhsj4BzBt7EKkgaQ09fkOD/hcfjlrIXwLum1aVHIIMxUgA2ZWkTG9
8JKzFj0Cn9tlPprUPKX896ZGSNbUnuBdgFDN0zMZfsT3OjMXtwOq7zfToOsXa1qE
m7Pk/QcV3s85P6+dk/DDUfixqn7eIqHk0YAB/TqzLHrPnHEDBAiU9M3d7U04Ew8L
xT0MxTg3Lihz9lWEQwPefvNTVEkwDSj1h7xQ94COso64n1z03gAou7Uo6JjfEHq5
LSQ1FXuFeQrDGa2KcsbD/3zOb5z7Hi2PP4IyhCFZWNoPYtB7D1DYDQQLigAv4xus
GS0cAp2Sva3HKoCB9YOJqSgC+pwGi/kEpZrXeHOQMx+aoKGoCjlip4vcRnWMTNJM
KW7AaY0GjmoU7uhFyka72pj4r/yrLzi+hdewSRj4r5LbNTgZRv3I6+aCMxC6YHjL
HsWhkUmqIAJIYd0xOBTIA1VoUVLOZmbnqKO8K9rG/J/MxQFaxJnmbQVPzEbuf/vH
xXaYxbMjwYqNDLkF93dTtfTXp7/sWTja6p3AlpZ2wODxZ4yeWUFpK50ENYiinfOw
t3Qt/9OMX8QN3eq92MqhxWiJM4RNkGR0iH+L8W9Kj2RWpCMT4rnQXUK6YTY3HReO
SjLFbboO2h7uBnGrvals93gQyhYApawBSdT6qLPvc8PP9zlmwFFk9wujLeDW49YP
LU0hun//sDREQcJmO1WRABmwyKyOaaI/0/SvvrTuiU/1JHxXZAMjRFCisR5MvETK
3unQ5V8lOEDyBtZEBr1E4X42hfZfLkoEu2QOAFb2vPkjcEUYWOqoxyjTv42kC0za
PN2j2F2snewjugzS350NiTvVvUosWQ2iMGToTNMju82SMlpLjuDqwlbQrdoZFZQ/
JBGpJxazf1TKo86NnvnGqzlDSYj5WQ/EwjBPKTp/4uu3ZYw2/2mo644ahWju1PdI
7kTFD1Oe6NYEQFVXNP+HTEME4VGdFuP7v48weFJB2E0yGMgFnpiOflPa4URWMK/a
7QClX6dcKfzPcvLdzO4AWmpPeQ4wmx2mx4FLHqn/dH9OfMtfxyleb0eaPsZsQHwb
tGZUYv1n4e5Tzqgtj1tCTFhIXzoI2FmM7lkrDwGe73GsjREqmzIILlMkYtA5zrwt
/Lrle53/093HrGkcjkelywOcs7mW5BIMbXGtbrnL5s+/DSqSTgZG6CTpctP+f5A7
fdVoD2mCPevmIbUsOpY/qGany0cze5e//AxNPAewndkii5IvAv/Bzf7Gqz7ivLn8
k4pkJWnP/YiWMZpqiEIKa0qxN92FNQ0vifpx0UF7iAiqJ2q3TG8dO18OoXhyl2gL
BPpYmdKdaALy2hl0OB1hxfa0yYdA0kNlN5hv1mg7kdeM6RKLBA2MLhKz+BSkGESg
ATUj8f3XPcjaE/N5bEN+7VXwx+suGzNOqjWodo63BsnDgF+sJvgkXjnVr/j1sXFz
FoSvl/wOEj21zX4zfUtyL2cCIj14ReZFISg8UnyA/f6IKw/QShJyJqL8NOdA+plr
9etihzSa9qUHix4r9C2BXIagflMVCsabwmpa/eidcmvpAI8Rc2tJH87roK+v2IyN
eBlQ/ZhZGBhWFvDslbT0bwkQAVYxx6pjkJU85bOVfY7ylr7HI1lHz420eIpDtLB9
sxpGdGDUzoWsUm4rTq2fAjWk+ijVmOVfDbAJmXcSkdQfVigLb9EzCp7S0Q54nS8T
Ft4ONrgNRr3rFteta21m8bbDFxqIaLEEJYwM5hzmDtt4H6JCHDgJ58zFtrg3YKOv
+lriiBtuYy0EBL65eaHtNUl8ddm4sC9ZVFfq7/S5eBX+BNlFyYeNPXeicEb9gfF5
v/2JMTeMfC7wEvFGI/dKs0VZTFbkvscYcWt/EYI2qX1vbTRltq1G4AWJ+gFHZxNA
BQs0VJQsxlMBzKagK/qQbtoBksJ0ZES6AdRY9eieEw8IefLkSTld4WELe6iLMPEo
Z7jeqpfybk1UPbOCPd63K0O1+j06KgjVmkCl5ca4J6OOPVF5/Rfe81qJprjbTNO8
U7nuY3qyz2VE6+07ZVntsGN85KDMTg6Ns70DNiqcUYNsdTbCrvWDLgSHLSm0OpWc
8H50Covo8dpmW3ewMHUJ85QSk/iAnQwjK+MYe2usrBTzBW02OlVrkUMkbm9DMXUK
4BZX8IrWIpIigH+3iucN2TlUv7AX45sHnWfhK8t2mspGeGmt7PqRtj7Hn709FuOa
ZChUE6zhf9W6lvY+vW3SfC02Q8tjw53O15IeEo7Oop/A75u4YWHA8EYd97Rdb59H
/Ha0LITUbZ0mV5ueGRj4UkRziu2VNhLV8ooPU+tVdvK45Qcv4upP6jgs6uhh115+
wvjPG1QUKPDfccdFfItFVfiGChNJ/TD0U6lBkFvvbYx48sfinHeiAx4Na4vSZ8MT
boq1cuB1i/4g/MCK4YyPtWL+x/lMBYq8DHWDj5eCtAry30051UQMXbtPdc7L/LWF
WXUsJ6UfunRk01SZDXhHQdXL5IJOkQ7z1lFdqigZikINZ7IQ/v6DBQMg+TqzRiXu
nFBpdEdYaIosjONZSyvzB50Ws0eSZ4SVkRUTqohKTEF3exqAl1wNkgY29MSvlA23
QyIfgAvLYY4bPScaNcHORaZsZeacEdfYlCVVzRx4cui29kH6gT4o9V3tmrtiQsjc
JpSkIYvCNTXc/3QfphYCzn5X04U2dlKFDUa6Oicr1/UbzrXh2ZHq877AR5F+59a8
497+EZAC5v4MZGpMtAFECZ327NbZTFiOetfYk4HuKwhUs8XLAjSM8PBCkBNoXGOu
TRECGppjbQZQb8uIfhusDEKCmKq57+FjFAwylbFi5sjOQBC2LZo/VyBL7aERHO8K
nQUDmvkLVd4K5otdtBr8TgnmVPt1QF6LYFXt/QOY+V48GBf31YkVLoPKv58cPrGK
GO3crFe7B5S0wB21KJvKkhhHXqYteEmd8WPgkkk0brRCZEtfKsg5jlXDnzT2O2Bz
i4rLybteMGcx3JheV85ZkmPnKzyxBW0aJrw/N6e0ryR4WeeMDGLwkTCqSN6gWy3G
0gUOWXLt/lTCzrwHCiPTrAAb3vv4GNLlhf6Cjh/lXSbkhpY1kSPfNeAKrpyOzcZ+
GH2WCMgvllgQmywDy4ESUKBgly/1Y/JN/4s9hriYpJ7/jATPpWTm7ZZmfNgETBs9
qkm/hKuRZuESAZGDsblCFjar8HZitvX96HAsYcLCMtAhZAiVLgWQPWqRYf040pMO
i2D/ZCufHSFnHJb7wHb/LO8Zw6bHc0CGgDP4CvprZyQ4aYIoEsyt9+MqqIdQ3H2v
BJkmG9ncYHhoSUDJtGC+Iu5QWWPsc8Liaa9wB5BLEVB6R+oSTfwInDFRvnZQ0d1E
J8vyl5Sd2pLfarqPXa5ajx/jpTQOH0fVjFma4piOcjyKEQCZccqeIXN3UXbTffLb
5TD/r61XNmI6CjRa5wg1llzflpVEUAxwiUmZxicSSHIKnVt30K1MkyvtSxJyz2UR
YFBBAfgqcDRIWsO6cR8RHm2ihgJK8BkGwMJabTPNCbPwA5fAF7ZtJ/bf4aZI0fFS
LRh1MLi/P+9LTMCp3XPTiWGnyo2PFg8VerLLfhNi64zC75G3N5GHKgii+2khL6te
E9HdASLqINCU6RJpfPJW3gkxiU9Q+s6UvKVgyEZhSVxRg+UhS8RXZkgZ0DV0ZG3V
PQUK+2D7WzSnYdaSh/P63AMa2FXSj/3iZJOHxSoVU3dONHtH/goyKkmRd35f+Thj
YAonTlNe2X2LyLR0NPp5ytgd3+G2C7Xi1qDK/Pku5EAj93zhluig9sTNGTeXt9n+
phSSkRINEdbdSBGVPfofRpprgQvdColagCd4t3Lj3hCaRsjp87zYbrf5IdKsBegL
zP5VmIbbfKz6fAy7O6frb4u1H6TZu0B5L4Mn1Meir29WUsn4EoD4nSkkEYp0txS8
x3QPFKjP0OWsYcIex6YE9De9hKqjg1w8y5EUtoE+jnqDNpoa9VlDIYynfBjX1HrO
ajHRO4tFIr9T+kpB/CbosYeZAS5D5mUcvmW+gmJTUf5TQzGMqMaNJtXjdz/teVp/
q4ZEs2NgOxYJJ7r04xtFz+rtohmeMOpqpqqlYvDQCqDsZ2HI+7YsiMS+JwOlMGXE
c9IgDH/wpvHvRUu5zeRQW4h5e54HXpIF0+9uniAYmplSxZVK2o6VNHUQIENF8DkI
herB1vRZXcXHSfiE9cQES/zhH+h+JU2Fv7o5tJmUxJaNNRhHmfiMByc4Zs734GEG
zuwP+NnT/VVEU1+R5vEXCrf7pVmEhKA/bfcle81W+akwr168oJ3L8RMdYrrKdCd9
LCUjbSjxynz51Dd+Zp08Ycm2DjigDpbfu4axfTH32F8m0nnxnf1xrUlin7XzY0Wa
M6eJY8ZqldQljpyYuwvuBHmwncHs128WHOySOKv3J6nUpvoD+wOQIJ6YaMjkRacg
VBIoHCvxVXZLgXGsbSDQMTBSEMaFwnJ/EZLUWSdiXy59HeWCv5uA7iilSaLyD1U+
rYgTNcrlyR1k1kdB/kh+nz9fltBYDv7BCxa3FseqXcDvxUq7RtIxHSmAurM9kPhC
EoumxQWNGuX116NLhkNjH7ZHYGSmjK3bnD/TKw4nCcqscvgffkqoXkd42qbnJwum
mpsxHur8gPrtYiEtokRtFWh1Mh0/+tsXrXoyBaGlNKI5RiAeyDou3yVYHqXA2u74
UZCXsrB27IqLR+pW332rAgjrcGBCZ15nBo62pQclkzvmmh3ZQFUHdg/Ptl7Gq10s
jtWB5jt6KxM6I32CMFJBiF5bTCTiy7nkzrqclNJsCOm9msof3oZwKhG5xlG4JLQK
n9SDvcELXBbOXTmZB3kgR0x2DairDLXsRdx0VFx5w67PMPHLqjZx04VY5SNC+WJO
WFx0TYwF4ogMBUglI9hEtPoiWVf21krR4gKhnttbyF17o59TeFsH3D8U94ovjx5/
WNYU+zXcyqPKvvCRCLWqDsG5OxSuvKACH0czxzIEYepM8lmw+U+LmtK7MetgYjIp
nhp4BCgqx12hx0J/CR7GauZ0cTLdc8BMAEGFt60lrQ065sQld8Uw/B6oy1uMDyB5
imZtVzxBWEOKDVgZ/d31zwm7aiySsTg7kc/yVktfERaAKzUf2f86PlGKkt63RbqB
f9M7Ru/FiHW1TInaKX+T87Ha1BiRjwBlIY6YADU37jW5lyfYMgSncns2wlserMoG
0CXAfmXOBEjGrTOwTbl2MXw9ZURUsrv430wL5Ls+RRk7tD5FgqqJYCExNXD8h8TX
KCPakaOKRHwX4yWv3VFipvzPM+wcL7jxm9oI7dvW8orYWTycs0033hoxcOiGi+L8
hGgGzlUOEVG0FhC94c9O3FK9aPvD1fEznNqWPC/a6UJSiMsyDWe3tVNBjrYJ/z/2
zjwNFgrB/5mrTPVenU9Ybya9OAPA6b7KizsN0ERUlEBO2I43fT2S6GctN8WGB370
0k50hv4MEtcf76RNZ3VX8rQKv6veK121o7Rp9pAKlogBnkAU3t+W3fq25yEKOOVN
Yl/6ZT2kVgDkTJLB232eYAyfUvd3l69Qpjf1Jy2rzwpgXwJkvTqupNfV2r/2mkne
RWUu8X+pCZAFmGU9lYplkq1N7wMnLXug1rxdAosJfPQml39TdlUNCWSMfHn3QSF3
yk/AggKKm7+EUipB2jRBpkb2qZbtqwLqdWpTxEYNPa9GMKGJog0yoMVpFGpW+TKz
qu4ulF0FrKMAN06hLhr4IxYWBnJM2okaqevDxcMNenq5BUoW/ksUECxHh3U4VzHA
TxEwYgEgFOoLW1ThYlfYxGS4gACsMEvRCS7sMo58NFxmq+TyR1kt9rpwTrgnljAe
7Z9xk4ZYWyFp3VdsPgQLeRcMTrWzaqmpwewqrzCKWt59bTSHO/AXolvovdrzw9sy
CTrFs1Nw6l07C5TMyuwFj0w+N3JvKt8HI26z0stJxVz+9WGB5tOF9nOXKRGYH3pg
Lk2lUoOPCyxIhi/3xY8LmM17WGVB1qRyQitKl7RCx1TRmcOdGJIb6mfj9M0VQerS
4LhXoa5N18VfcTi0QTAmi7zYrDCYCHrLLO0LvT57Rn4/qYPBAPzpgBsjTrQLrKdn
8w5GXSLVcAve3XkIv0d1WUilvYlRycbp2+Y75keX2sn/gb1nAECjkzb3PY6WTacP
IhOErysE2rWXU0ZU9Um3pQT94oe1JQ6GxM98QINcb1IGinApSdD0oSvd/BjtT4JB
TuHey1dvlTrGILClBj+UBVjyHEUC+Chrt8eJcJl6fo+ELM36kgQ+hnlyrZKj0YsH
zINP5mN/C+SHtX1hyY83UxYfxyYyf3QCZByHpWK1rlgN58U7MxwcGopC4PCBdLJY
cBUlIZYzLP/fnSjUAzHYCO51yhgc6PL+A/4ls3vJt9C8TK0gNiixGY4xuzKCMzEP
NqgDltNOqxWAdaSTq84d3tIjzjIVRnovT2DK07SpOlxj6IXrr06fBETiZ1aGvFk9
Sv8vKRpXZt68dARH9OtjGhoFgxlVtAw0VL0r+dp72DfZM6tRHXcGmElByvnxfcfE
KILMktN10iCBEvihyeJbRkFg4w0RxPES8HsgLEo+5Uz9EKkVcPaNZrLnHb/oYy0w
8bdwtkJSuiwysezHyVLEvsZXwnKLSBG4boTqbNZ5BoX2pAbBEq4QesCPb7tcheW3
98ozshdk6kTYZerOGARNA7y+4hyeVw1KNplkcNU/HtBtyd4QJ7+CSWU+qY/bh9gU
jlRx523Q1t0HMrGs2tejky+zPIOeioHg1u8skfo/ox/HHNbS4RdYvpvef0NiKEuY
v4GDxvssUdAzugMeqUnG+apYUjIQS91BS5BvxEN5PGamrDuQU9jMC09StTgZRrI8
CRlrr/+kp61M7RaO08gB4vJ+UOMEo5nYrQZh28TqNB9qXVhSCtLn1sOyvjbYIKW4
hSfz1CShvtnPnrU+WxD0uCiJ1GPUTb1Gqyvz1DrHMMcG0yvN8jQneQJB3P5r9JLE
uTCj2P3knwRppqeWj4SGBmFFr42NIPaWI5EqQvckzuhV74Aaz4O9KSTpSn8GIE1E
P8BX2HoY5kPR+9wjCQo+hGYK3OXYXwgqLOy2d/RJ6dGUewC7afY6XcNdKNR0i/6l
UIJdZ/y3v+mEKQBB7hwLYZevMdyos5cOYohvbNl3SSalhTmbF0cr29M1RqQw96jH
HROeGWkDpFDOi1b0XgRrC5kRh2WWvyinK5UP6oCWmUxPYduv/mnf4eVhPbwcYAjz
3JSijR4e334aS742nYZIZS0wCjy2PG0SMQ9msAOWr02PPW1bYhJf6b0acl8XpV9m
6MwUrjRzgQ6ogO0urtd8Gzxj/FdD3jynQOuC2WIbV1HPHbcNTAsexgVwDMND17IO
6yvu1TN8SPi6W7IgicP09Ap0cKpazkff9M7ualsqZamX5oUf/PM7lzVhpavA1VkY
bEv9iph7QB387lULbSNxKCMCqZrgiyNQVfUf1bLKC6BpxTUi7MzCBy379Gw5WQcz
9YDgL+Ih4dE62y3Wsdf0UINO0b4szhrVFRwyUmK2fmZL9VfjUDuqep7FmI/ZpcDA
X0L8hEzbZqE5+40zsk6rHD4MoHeuO45trLvIIX9L6Wn2hJ69MA+5ZYPE8RvBZ7+S
yYtrBoxYftAFIVNa8VdP9zrQUMGa1YJCP7kcdOv3rr6gyelw2ul5eg2iZ22Poft5
kU/a5gRmiDu061mhiGSW5s0k3IM/Xwzf3faBSbgc7/C9OLsWETdwrqyuslfLh/R8
rWxI1oh5wnUXJ3lLpDf7V4Af3SrWSCR8RqLSwyY8dSvuYx6ZRr31uZPfPy8WQM/m
VHBrDIhzExqViWbvwU4J2xEW9q2wP9ZoSorZqMi9jGcND7a0/+sRLZH0jHYBfcyn
P6fI+WOD17JCAjjTw3WStw5Xh8RHFCy2R625T2W5/O9pij7z44cbb7zntAbc9vHy
RB84dYXxLNzk1ojTZJGEc2vn8XywKfV89MEAx7YSUFPKd00iGUbF/9DoyMqTffKM
aFBqFtcSQzS6jGiVanSPNlvtcPfzyZ4aeFkhndbEpJOIwpfjlpx0phkeq+mIdt4/
LOD3Dq/RS8gBET1cLmC/8x58mHSHQxlZI7SM6uu/6Hn1bl2qhTZOW165byZexue0
8yHZLaB1L1s1loGMD3KdJLcT2GtY6NNdAlJuCS0kN5zVfzD7Ea6yWJ3hp30i+0bK
VDUz4l6RoCBaVMHp2oLol9mIHyRqEk1sBJgzyctnJH9XOWIzX7E8JLRB7ehTbHWn
U073rLGgS6uN++Vdgfxua8J3NistROeLCSN79mrSD39hHUOoPOR2B5Z9wX1cA4Px
hUY1vltt/dSsmwebOiLDp1EEHGshMdiBEjAQTM/MUl+tkQyjHfhX8nDSE7VdvklI
X42kCSXo1B11dSzZMnAGz1aO+zX1sQe8s8sjoP7Qn0LZRFaose4tX4pmKa/Bmomh
AZyhG/cU7qwYmM/0nJgfmcbpVZ/QqPo7awo5wQgxDF6JZc/pHml2GZ0R0cKmW/6A
y1KqsWDwMEG9Diw9zYjYI60zDX762wMt3QEYAQKUtODS4HZkKbU1x0mFWnB+TL3X
2O0uEmiEXzbYpxxb4skERkFKDJl3C+1FxyKRVJdNTthLyZI/pQsCOxTjNVJzVV4G
CBTs5LW0TCpEtos6uKd8prJH1AIzVvvDX0PodETwYgDHZ0fpWc7bzhB0ZByu4TQD
FjjyQpxBJCbqhD9ahXHqd20dS1TBZPShI+z6Q+wVvtQdiArzqarMsOEyz8Xtr1DQ
hr94zNacZA4WSO2/U2ubOgKc0X1XnoLjzMYnMyrabSlHkeYaD2cRF7cYAJ+aTgqT
cSb8x5qm5MU3U0bdtw59hODP6TVutYWWL8mv/xV4Gf91r5GXXhIWcavEfjB/xrk2
XGJ5bdPoLOevBSluJ4OtCor41i++FJGo+478GkP8otRfPww1C5MJbNJaaLROrL2s
2rEuio0KRj4aWfJeLrMHSPrzcgx+dZLsmtbBXGzeZAS9gVbOhJWZVYldqWEaVDLG
QkHFHxUP29y8jpFNpq/Bj+e+j00Kk997FVee8M+HZXyJ/ZxGjdk/W4OwfrK1+9Dj
wqyR/F3gatqQ87ppr7YCd4H8PAxwHCr7ovqAdYOO+VjgPabjFJnLPZGJPqf7wr3I
ZJ+B64pXbCDRoDGufvg5bWhwPMm0Y8CBR6UW0Iv/PmwjOCKajj9qpQqvMSLYi8XB
bQN5u0B806sldDWPMJt2gNJQlQg9D2HaAAXF3PEzt7PlthmfBuftXrF/EEAVWpJ+
+VDzkf9D9nK8wANfHVoNTHlAjRrRR8x/6gF2UVZlokLS5oH0I/J9LWdqbOCye6B9
Pem/Vy4/eNubCdCKTbZlO7+rUcUHz7gbQDvKrF0t/Eti+VSuTXjsL3Ebccn06FmD
pbVF2MHlDVKVQVIZvfNvIr8pRXu5hyakbB1ez2FJuK1pGqs3P8IDgYyY//vEsUOz
PQDgIbuMbBPAuBscjM45z18ZxHR2oQI5nHVeCvtKCSYtNHlLUzMpK3v0nB5Qgw1B
XWcOBrKq0y3lVhLLFa8BqXUlt2HuPxdzcKcyPple/8DWxkF19F/Jc4jyJ3kHn4Gq
H5pAS+gTLKXz1U4Bp7jIFPYMVoOWbSADyrUiAfxLTYSzlAamyYY+kVdqiFfI2MIj
j88jYNHr8TzeAlGQm8Wm4GktrBQE23x6Pi2Efl1plA9ACFjg4xTRswMh93twfppd
OxwYlUTeOyEdWcNDE5CIdnTvijZxhTEGVtwa6YJQI1MP6wkqd40gySXM23PSf0VI
2oduejq4F7kcNqCSshYCTtOOW1kFFUSxsQQeTBcJbQrQLTccx82Vthh/twLHMzAK
8Akk9kO4wjc+TrDG4Tz+TcJkKnbhrRkZw5dEAiqzJetjI9u14hrziQwBfUhe59H0
vLESoOvpqLMkkmfvjrri3yq2NRH6hIoF/VBioz6C4y/7j3HGVomMTTrADAjZBoCI
oziRvYSTA20oXdRwA/HF+iFFtDbsH/GQSxu9LhUVsNiUb5oENsbmfEvLsqe3PARu
O1MQqfirTMqJYv9uV/3vCgsJf22u+vbe4tcIJx+pjMu8p7INM/lumrjGCzgTqBZ7
kzNK5BJOGx83LxQ3hDh8HQRrBIDN7h3hRh2hH3KJ2RUFgg9/YaPU/fenHGqnbDNX
aRCVN7u45c/aRQ2fStPApSYEl33ugec/WaCcvZKAB73UnhgeDXA+L3htXvFxgGSQ
nbelbn9sNy2clcFr/jbyaxjX9l1kR4bDIHIDrsEHkQgTscbTbOFTQ8OaJ782nfs+
YqgCHoGhb3UwJNqaJK8f5sZFJiojDusr9V56s8OMQdQ1Vxm6nE+9ihf1VmAWWIfQ
sktf93oaoQuB7aEwgENOT0Z5E9IeGwmmoefMLjlIN4nA3IzfBOmPsAC7w2Jsu12M
h0e8YdUi+ImNNbD/w8oZIYHIYhX4UTeCVY2NaGN1/GlnXF3kFeSzsQA6Z55/YyNp
mBNI/QcrXNFbSwZ/CFj0dQz0ALKRmuJMMxIKFj9vz9h3Ynxzbwl2iEqpozwda4YN
uIJZ0k5Vtjf3UCBsUqIPkFI5TPL4HDdtANnC9wJNvz6ITdv9cQifCWZyQHrNlmCL
MRdAU2zFKBNHsEljSYdf1wUp0tqFJ+dNmnt4CQSqs8RLzy/0SC0a91kbziUThFSr
jn6b/X144iyDmspL/zXhltLS8AZA5wz9rmRAGzzB1YnQOkgRioAr3Mh7hLs3qLeF
nqW5UKpn+z/vigyD0Cv1xEImIY5M/1vuytrVr8OeqfmKU7aHuXbzVQBbUxePcplm
QEcC8de2eq/V7KmX39m7QMcWrlB07yi5QlHt7NoaoLROAlB6JF77F2eAE9Z8E8ok
u1NrYjGyVjzZbSvIBXxpxAJKrRX/R8LqjLY/Lx4+S2T1XrA1/7VMDKTxei01gJXJ
MrZMKp7vQ6uRARVkW8Mk248auwT+rQqwNZM6mMyXacaLsjXfLFTL1l5ISnOTQsxf
pmBA10dkkQuJh4vTBmykIXOVoCs9qWxAS6MNxzYDbv3zET3O2J6riSXVdWexsm15
UnjxghegPyuJE/VvOz4QAs3dKUo+gWhLl5iE225MLbmmyQ7l4EYAzc8qZIZcPLQ4
6FQfL7gxZNhUOR46blFbiMXPeVfbevPHbtB8B5aeOY1FFps1VtK4gaApsjKVUuJJ
UtwjOPXnMUO62qtPjJMi+mv8s4/4oE3Ug8DCT01CSO/yZ95snuNSsIZ+IOroFW8U
fJYuUyxOAgGtrcJtSIcjSI8OTf6FdtnSl4ocXc6+RjJdACdZ6eDfKoypKte5apj3
xAuI4k7PohCnLQY7gNg+vJ37dH3AxxC+Zd5xA2Gduk5q+UB+n2xI3u9kWJmXJSQV
gS0P9I660PklK6HZLU7B75sGR5bABCjWj+570ER4GwpkLMfYj9KPP5dFANlLFZ0Q
KoNgVpbc2gD4l7MhwxITklsPKjZWAmgqt5RcclaYW10frjQ0TNjxuK92ksCHS0l6
qGIbivvBa9zYTJP2K19G96Yc5ysdxsFTuaVgTB6bg+u4VzOZxDsfcjcvyJh0ZET6
1xdZ/1eYmIDI60TI+3y17G2+1ZpM+5UK/FsamquEBZKtJywo7Dp9Mwhm5EZpP5EH
xxHhN+LD5jZspxDWXwE0WRTW5V8H8uKi/IPqa8Nv91fZ6ZDVw5wVTQ8MlbpsUK+V
0FpKmKGZ0FNIV3ui+mGkLMMgD9GDW5hRlWtuUxji5Aq63UfrMg8lz1+LTTkRhZVE
x8Y+uLkeLQpt/KmCfyPeyz26/vQVWBUqR9eyX3v/YsI76qBpmg3N0ZppM3viNstz
kPKdHfi1b7sNvBxI3JTdkkQV7owCh23JkqGXYLqZmkHIu4+K3trmo5P7gc/paU3f
gT2iIQqE5n8sDdAwb1Tj9hzYpr5lp9z4hSMxaMRsw2Buz7iTYb864IOPFI3nzNmM
Gn9AWrKUD6QDy9VOgypq0UeE79dtys2+OSpQneTyEIgZ7N5UESJfkpBh7eJw3nc3
vI3faGP0l1amgLCadzF1y6LtoaAjBYOkiX4Rdp63vIL4aqCR0ozbP/3oZIBZ234P
6CgrbtnO02QzLXUGZOdfQnMXtdAimjzPbUkQCU3949JB2yYBUzHg7kEaG1v6R+3j
Ro6KOjMnYqyqT+zBa6+O6JjFQSm9w7C22j7RzMoutHKYbsnSrlStoZF0GCH05C1t
iDgYdY181pktUwfIWhX9UcYeptTyUmkA72Yfu1s4yyYvn7d8Mg4lIsoiNGGxCG7C
yMNxv4gM5QBYwg8OwivDCNCYUKKJdvx2sZcywaLC0vFXr2XlN1gqGgprGLwK/7/T
nzPmFI11/QP6kza3DS09irIx0wAYLiCaHUprYWsMRJqFTXMtdMXBFyliripdBsOE
aK1hCreBLqT66TVLO7RYjj6IHdTf4s6U53Zh9VqEaJYJuxpufyEKDL9szRbFGu0F
lLctn1xhfDv9tOmtnw0DyMCrE07ZrYYuWKQpouR7HwAQkEo0Jn5HlBTHcu7yHHBe
/f2iXVLheouUw8KObR3qVTpX3F1dTUVh4VLqfAS2IrwNXN1rwibGN1AC2uHNQ5Rj
m6THozviniOVXu4keSj+KWmqgXQ38mSpv4++7/vrU05Gdotsw78N48r1kEXFlrIf
dsfLj3juDT/jnKmGfygHz4bu6u/tDl/AO/haBw8NvdkZaWuuWvo/tgy2o93dIaJ4
DLY1SOSUX+1WeL7b2e9VBu/kHVwreOYd6wOtqYylvDwQjXzgv39btHRmR48KlAHS
JsbLbwogrACI9SWKKrP5HRj3gQLBw/mag4PadJyeRQTu1tLV8VBUlSaP9K719W6B
LaD239qm/CXZ5OS5IzH21R52b/elMaARhbcPw70ZutoicaGmOInR4gY4mQ3T7Inm
kSJm7HiibS1RrMCVSAGnQELVilEAIiHkxSjMw4lhsO+mSkI5dZOcIUoW8vvii+j5
aLPC5u6+0dZyYPcl+lOM4X7JtOU39E+96a5cvlMUcrvSRYfu11Zqw3PDeZIDmZ2N
R3731QpR/xFIF+Kllsr0QdWtNfXRDFuBFWJub5SdFuUwY4C4vTQkRHYE60n0Vrcc
5mzB0ggQvOz1o0J7n3qhtTjdrG3d5txD+2/tuZCUlyQlIpIhchA9DTJiuDkw/vpf
tJAOksaUWpy7uUFZbe7ULoYeIkcOdBR82zM0ZeN/LspaF3q8fGEDJPpf4lDI+iXA
xTqdQoNy295Ag3VrxTGHlQQnuGefzyRCTagLBBTtNpk6e64DP0P4bFAdiTTnCusO
mMEqYZRMQYYD/G/nNXZc4J3rZkrD6fMsMb8+YG2oaFrWuRzkGsiIyP4vgpmqvGb1
IuTJN0hgTh1HqB2RZZ6hYtvwIBvYFvbUrEmIQmvO7la/JUd45be5JOLFTu4MFAez
iGAcgepLI84udWkQOu5A+P6ueHzToTh4QxAaqVEJ8ozOYBadHrhYWNjzk+oV3edy
cVAsQBwvwCfyeOveBl8Ko/KcydTb2RDiI5cpeDrXuztOy03RTOC/VXHU/h4KdCb5
N3IgEXMKuDhSjTi75BxLttvwRkRmHombXtjMs39dGaBURoPcfDuvKiDmSEKCLws4
EQcZBce8KrQdLDdzOLpdxc6W8leJj/NEX8v2ctE9KA6NQGsUz4S5SbRKTGJQ3Dcg
F3ZKKayy26IrjEk+MGiYbSZA3mjaJw6ZDjM0wsWrKITgBRvgfOreIIQimmOy0NkI
Dz6HS9FKuMv7aGIjfm5iEghrPjKc9CdEgJ5tJDfHFwfh5wzFukyJkdTykNIcIVrm
nKa8F9o9cZRkM3YC/i+WhfC7+QcSS09gpaeJ3WZHPf9wlo+4ZUpjR3+xIFZADjIO
MlczNb+9WOs7vsO1mbLAfzWGUHoszOyILJldad3mpHy6Us1ah5ZnMM5AcxylRynM
q3+K4pZgIlnQfEkmtlOi1hOOB5CoD7H3rlmREZ1X5hUxaqOqufE9s9FfPzL2V3XW
wDXdB2pOKSUeVJQWwyMENaSiT/SDmhkLZpxTVBSA+ayUWYH3WST6Vgh62wbRuXGR
2F4QN1LC3cRhFZd5kY5CgLWjqfhsdO0OriVzgVDWf7wrSLC0NxlI/3Sgf0S8SEy3
4UkQJi84XgiDD3VmNcUXzraxDI+FMFuloE0XULuHNnloUqSq1Ot+LayJDRe5aHTP
BwNgjpFDJLH7PE8ENzdZVDCJdkyDHDAvDOQmay1JV1ec8xK1fUa2leLKpeHMwDIk
5xw/V1AG9Wz6B0Vevsn4laKh9A+zQo0KL01lRXlNhbKcJMlP8p1B/v4lY1eh8UtH
bPKDrrjY3FKaTw+gNSLN9p7ZZkOuCT0jB1u96+LwJqexHehcriJvE4UIp4X8BmsS
rqlpegLVIx9NP89rW+rSpKTzX6oDCGiXs3ilh/CwSfIxnNKaT5hPFm1jAO38sz/h
dcQpC22FMZOzCKx748l5FsmQgh+B/r8uZKlRd9EiVBLi8sied+f4z5ZfexOL711g
e17PPwYfb/JG1QYT1DDHjqVPQtL8KkkNmc1zFroEp6VhFCVtc1CkqxBngRuzoIx9
ByjN6J3ez5o6d8P/dH5lgRffu8R9MDPYPWj2xF4NYkWVu+rtnZDnB0IBWg5ayWaa
eyCktDKULoxx7t7FvJmP6tp3qMIhhsjhrbLK5ZjD2JSgnBQJr3cwCKezWWrq8/1W
eod+SlEBu+xh35I1YK/KiL9eTfcQ+VEOWjq/Dy4DtpUsxAO6K+Rzv+X9ot31TTWY
DDs0fHK0TSOq4OW8TOjajUSwOtKCbvdsk21wBnxJWAv704V6Br8F++8FxafObXuR
5ppQBRT9bbyRYdyQJ3pr0qL42DPK2kFJQWBEa5J8xKA8C9XUH2v3W7BEQCRyRzJl
1Qrwp1LOvN1x9ds61icrHFMAhDjILN+XKFgh5UZo8mgMhqoVr3uZVwE6REFvNLnp
dJZK6znr/Fiem+Hlq9bQs1V4KOpMYLETKh67RN9+Mczvu2fpgbBIB+/bzqO+eN4W
uzY3aZ7JpI//+yivh5m5jHrsTWHuzlcL1fT7B2QSwNk7YwPSADy+5sojJ2oF4Rip
WZD8m9leYECBqWeaIJWtQWnenGDZNYY4qmyYqBDUSa0ihPX/1FLLlmWBv6Lyua7c
KFLLeqAsEBEO7P7Z9ZfqsYjfayiW8iU5LWpFlwzYgPy5WaromMDWQIbM/DCwTf3u
7fkWe8kRor9TrQDAOpA92DVtQW0DBI2hNF+8zDsRAxHWtZFa3bpf/RXk0zYGWOQI
mO2xdujf+x023SZi5OzrehiJzkkUPKg02aWM996haDZLNVlJWgE9yNfkljVSG2qh
3byF3oNSG+o3HnQI7Dg5OA5wxSTY+gJVTm4q1lSaXc+9bKVYASnZIf9WiY5Fw2y/
n0HAkBlx3etvLr1v/NpG4RpCTqkTh8pLFxZxmmNZwTjE+7thUcjpkkM/DRPBeEZc
J5GxDZsQkxkiMqlQngFOTGiXJ2FGr1RCdnc513pNgVh823jDGXnxASGyx/Kj6kBi
wBjlIw3BYd8MWce+qV09AUQK0fIQkWRi4Ec2eTODtomSQ9vn9WqIxZOZuXh4kahw
dibaFtp/icgj/wj9m1YwNqJZhWnbTsCo3opDPYwwKdpEPPwtOBkv3xTQXHCYGzOO
Iyomz6YuRg7W+WLV3/SgWAgUOUlc6g97IcJbq1b1s9IDShMjLOGuQbdkNKgnZw4W
ZN0QiYkDAW+KqMDbrXQqse5ptLyo4gaZWGyfVrF7cZA54UJwqqlbNpnuOl1YtKY7
zzjFUtFj1y4PeKIXlFVwEt/cU/oBmj/yonE+wEiICHPkxpvHWxXbgPzK8n+bL8ZC
NA1g88AHrQx4hcpxO9KIUU/i+Efv3hdLvo9sqURikaAyKlbb4qdI+4IbZyBUiqh7
VgKvWJ5N6cHwLVgdWuuob+EzktV/Vd1XH6ETjX47JTZkqyA3qEf/fTR8gElCyCI/
u88/VdUNzH5x0kCYDz8EWml8xAQAPWr06qIPi+3BLBD2AGrjtaCIOHrFsgngwb9A
4d6R5waa+RPmxoARUmLuk4trXkXxKL0Bsbtaw96CQksWczvQFMajaKICzqdQLVGi
P1lFSme1IFuK0SuMS4suWPNnjZLhtLtNJtWky5PUaSIEk91h7AqQQAxyAeb1kbCd
c6jBm7hG4Vz2+g+YHpWJS3to1XXvyzdJLRThvvaRaQutAPHEvOO43+3/F+Q5Ui7V
6ZqNKnNZY+V2I61fDE9GyyA3yzoTp20/fi/MqQ3kb3ykuoyivbH6BrdTOJkqBt+F
T99WiJMg58DGtn0Mbrxo1+Np3g9wZikHx9sAmX6c7BgDJgbTKlp3bvehRi8W5wkP
T4xgilGyZ8jxKQ11E4CaWxLDS+lsJtUdP1kVq/e33VnkzKwJgwQmK6Trn/kPf7xC
9fx+oH1Xd+B+nXWr9uMpbhkrJEF/bN9UJKEvxHGHJLYff7kTXV+6EPlNztqItLya
tO9ZG27sP+Y5VPEziygbljE85HKBZzC/EYb8Ec8Edywe9EX0qK3cik2XQfze7vxl
jLo3EvKJCKOtJnme6MVYyTixlqg5EIYeG2LdxSMXLrEbHps7LUNClAq5TTl0a2JL
8BVJDj1epEYmJBLtjaOuOWw9kdfE0oZwFBcOl5bVIpZiPr/v8FJXoPxmA5jMdieW
v0ZfBqcVJLNchWouqpXnYX+Sppfy75m+vIeB/Ql1tt+oE6MBxk1wqdaRighHsNpY
nErxCZdZO52aZPObIQU54K43F9x7pyW1LFRiauWyY6tRE95iaEcSkfQGLqEhmA1L
nEXbCtR5sPvFo9llLM7aaRhuz8eEuu6HnOhaAaua4eXeu7Zbmn9/lqapji8/pi2V
Gk3CbSYbqSxcHtZ+G15K/C1O4Z6KTGv+feHpGdd0v2RICcUXLeUrfvQuE5HlHCQZ
Gx6gQIFNOnK3SvGwHRRcoaq/V1QmNnnKTaBEA4ONVN9dyzCGiwK2eXRfIiroMBXn
Gc9uemLzLjXzQ57XjuneF5xTEya9+0Kmk51xynxKjTDArLRYUkx2bvvWjcQY539w
/mT5CsAXeMhXolNpg2bZ8F6CBmWM9izUU0pg6RZsgjFD/iXyiK2uBEDtwfuUbjaS
wFUCPZeHKVS1P3dwSeWs3maEo88v8lgSw4nlpO4ZHk/fDfhJdHerqKiGW3m8tjm7
R3eoi6BCRYea1cQUy55uXHXt29YNUTJH6nZhsdQz9Lbcizt50gHBQLtMQTsky1DI
1NLQNO5p5yOzzFrjLDq2gyH0Fxjm5sz92DfgMbGmvxTSU5e8Cq543QqZkXzlTgFd
rJuG0j6IzU78FbjTNVxg42JjriGjMhHrTBF0KQF/SHgN/ASMdsMJimpWHxHTEckH
5sUDiLOgGeOY2GJQ4BeQB9CAUYeDGBfRwLYemMRnouAqHxmVx0BOozhfwJ5ponk8
dq+grknMD6vUflBTT6jjXicIwkJ/6SZuKcvXYZDkANeueg3XOynFQi6KA7WBVpV0
OjYrdMV6l05EHfMaCv8wrKHiSaVTehZGLt3YMeUiMSq62z7P3bjvF1B0pdPwAxwM
KK4PJLw13VQVn+tdR1CCkm9/hs2z3zFIEuKb/nt9cUVvLj0xfta0gA+SjjSZfM/z
s0aYDExl9GXPe9oLI7Dj8BHfegq4jXMTzzTtsxOCaSJdo7f4XK/QFh7f9Zp6pkeB
R5vSnTyaY4B8FkAJ3e9SJk97XTSzDv/m3TuCby6+YCafIrsNgzWCPLbuT5Yi8lxq
WB1b2ktKiN8WW/wD322UDqPPVa9cFm1nFf2uxndv6hFsIJXIBsI0uCIV7gwo/WSy
UylozLhVQSGhzli5zBahH3iVMYMlvEfkp0VVl1KdPU77ksCwFuxcpE99VBhenrjV
npIhnjZUSBUzSbjKGeEbZA4JoCebI4LAnjrjIlI6rMVgoaKSzq1g+g+iy+FLkKfT
hxcZwWB9qXoQj5Iy48//G4/0qIPRJzHhCXIjlUNE5Q/FeQUh0QVqTrOwiIr2SL5G
coR6+XNkZ+PIfEu8SpIymFGR0Odj3Vnn/SUJLOhCevV/9kRjuNT2ns+FEv5yl7iG
9MeEo/kLyaIfzZiZAlxWLOOHxlSYT1C9/gFczdbFWYekyus77bABZfP1hfiAkbqu
0bYlgkGWtRZn8lCf/tko6M/UdQ3lmzS0R0/NtBNUacC6L3CA9bqYo+KHJeIVoGPz
s9aHgMu0h/Ppy1LXXJUBl5YF5pSvoRcuwnUfNhboHpce+Yyqe3aL76f0XFb4Ryo3
iGzIVJCm0MZlc5UVnJncPZsolbM4/68VXK9djYhKGCihvYiDGc+TqnVIaD+tHI4w
B0bmvjd6HW3BU/PiLPWq6mM5Aq8uRu62XSYw1XFw67w8V1+U9WitaGZhSUNS3Y44
jfub6+dAraE4Sz81B4G//dg8KAq03EOySuovOOt2Ggzu+1JRW41qcdFwPwYLwNKx
TC6zdKXWMimlw2RcBOSmHMRx5ESYOoZJG8FcsmRYXApo+YTEJcsJBRAC0e2GTpGv
j2nqPXMkdEqlE/ZYJ8/PGaDOBfi9LkYxiXyXykns5D5b6Ga3CBAk5zYO2EKQleE3
r/7TkOnaoAMGBcuHsNo0Srb4CiaXxnJ23NkiM8Bn7sPbDnGr8iREqPs56I7rDJiF
1b2YdaSnqqsp/4eSWOKdex6B/eEKI2YBgaWhuWiGFEUsE4y+O6OPQDqnxJ+a7qAa
df7BZS51APnAkK+MDGRj5xF4xgam1pxT4+Sj2XsdljLU9b44KBPnZtebYVl+Vzl0
8bSr11m/46Bov52V+lx3MhTwg/YMN+RhDsMF92TdBVEtLIjP01c3dWvbjOShGFTX
Li3yHO8SJzLpOBVtffsi8ygSZuFbWHKgML6QLQrx8/ohkZQLKbHoxbE7cYFtLdnj
rVUQDK5WXx31qvJbv5AdVnfD+h2hUmvbfX69753Ze3NBHytguBO3vSiXLpBHsMmN
BD7Czd4L3eXre27x8ePxuj04uxNIn3I9/5foS+NYf9ydW0GY0U7q1RF8uQuUiFLg
yEr9C6a6kBXfOrQkNtqmMYf4Dv1KjU+S5bO+0HJxkFp5mXlZUi5g+sU5V+KJUHlc
wgguyZ1p0BcG7sfYVFQaHN988QLfUDPitgyZvqO7M9cnyLAwuE1y6fCkNLJYhgYa
/J8f23ZXCpFDKVSJ4TqnvX8Nm0Pd1+/blM7vS2v7Exg3b7QKWZxMO2CU2+OEdnbe
ht+6Wj4Pq5kc2ko+OfE9YEdmx/B/Ue0WjD4xKjhTHibAJEZX7mR9f3nxQGPzO+M9
a3bhAO01J155iNJPaqhOm0f+YfPsNpZCNUYLdDjaNbGK5eSyb7YamJlushbTOO2O
yUU6Z72kOiFoxp29Zqmdx/Yn6hdmy144yNPGF4QP/l2lyBi8gubA4DNcyr4s/4qh
I+nsJ+sJqcQF0aIczqoSi24ei8WfiUIu/Rvtwv+Hr6F6IlNVN0Zrz/uRzgALaPoQ
c5iU+beW/h4PRmS95nc7Tl93E9gxiRtLDniGDLSV5QMnS8enKXTEEx4iIxlS9jPa
Tmwjx08gWU+Ge+yRV2u++2xvTNf5A/x7SG4BP6nNLPX2/tpijMx7juidR29Gy0na
CfowHHBUD3at1S5g4yt5F5AFmoE+p81uPzYHRq7Yia/atCPPIGBqf/422rlDsbKo
ysp8fdY7LmKgxnEzT7BzdFCtNbuFr5iMTf06/Pzbbhm2/JllMxncSqE2dQvqwdDo
Bh/8xCOfpgJk6D88AWFXT/DAGGJrCERRMGQXfoDugKcGVIjUsYu6E3qgO6ugelP5
j1ffasTxh7IW8s0KWMqk+blG97nNHqVBKceoYiYpbhnKBJv13PTUwDKd/Mz0N80D
Qm7Nfkp5QfodectKEFhJGp589D0w5oGs9kdK8e14JM9ey15VkuR26bN6iJxbS+Sb
Iod0PK9tf5i85xc+Kr53dFh35IJSuYRDHbLtXvBXE5OuBpgbYC87NP5nyUfQWn+2
bE3dF0S53hT6DaW/M/ek6x+oPshTQ8mnsKtFODpFoxRDAMuzghiU9wYeB8DWok7h
NMG4HLZnHBpCg0A9MNKCTJB/jR6nxTvnQWy9uPuEeAY7bh0c+K7BgoTRc2mKB3VK
iylRagcaHr0puNZW8bZkKrBLY9nbj1l9OLR1/sWVJ9SPqMfNLQVXWo8XymmThZ5U
0i0qfwWmg85aOQRDiXMjT2SYv+WMvwiBX7mAclJaMTIuzE6YVlNKnDqcDLr4Dbqg
lduQH1LtlRLiwRAdfQVFUpKCEVCxWTOZJP589Nkn7Q9gX1xGth+/nUjRXPd6Axcv
B9V1dzkG8Jkm+VmDsODmsJTtQOwc42yjZvgwzDWzN1JWxy0QeIABGfqie6HFyyTV
DtOx5X+q6M3b/ZGUvcSyoSZUCR7VfMXvJUenz8Zwg+2u3ElnUIQqPQ6nyhWIn7BD
cwoWHjEnUigD2QrpdQWi8aLi8DnDZjQ+jxa0ViOzBIc2UFwDz62DI075C8vIbYIp
vruM0rv5DocuSgV3LV7j9mGx58ZoNd7LKuAO/VTizhCJ+VvmgjfvFBwV0hvmTx68
H528kabZe0/JzUsCqD30XmqnUlWEav18NYHM7yklq91PyWw1BM6eSfvE8LRHMTRY
g+aeX+zROvx1uaMmiy+AeWQP1+cGIAVMi3oXDN9GOEtwrMsYDDxkUbIGPfxszJkC
KqwZObWQJCOTos7NiioLeB8QJUyPe/h4CVY2toVKjyJKeMHM22S89oh6V7paR9bu
gNf6xzeQxJT4t6pAdv2QS71Abl9tbB/5oMKYV8/9TtCH67SAoNq7/XiUi7WXHRCv
DABNRJfIgjIcTBn4rMwERgwUitR3IyyZpxisUiPJN+AAQOW5N6iMRPdRcJchWjvt
6oufaVO/CWf2zSUFSzfxBBfHS6n/EsebaixQLPbIlmvL8Ayb9BFKAunQv3Ifnj5/
6aIK2kK24JAGaPu4cOIRns3tLVQEvY/i7dyIGL5dlojKB7L8QBbXA8lZxOooDOSG
B59bKlv/aJnZkyhfoEy065Rypy7hUAlDHrP1IoHmWV5bJQpvFBT4+ctns4q3HlJf
2vB/ArnsPZIZ4FP3dEvZxPSOE1wE4nttK7xGROWws7WRgeVnGMjmwDZDTh2TYeiK
SCVZeBvKzprfs1awY4QOFW854w0qrNU6YZL2Jen8PxnZdkUfIK+HG7HIl3MLstrl
CgvZPJFxlpL8BU7FqKw/Nt8ZoQkaleN9LtjtpSpopRqgbNIDyR0akLby1RvKfjMG
ELJEPoJQT8zCob+hJwJnZsO+7bDAfcJzJsVZvJ5Za4rCP9/K1F+ViOr1Tbgd86ek
8wXXj9slRtchClG35YHcUhOfQYSEIdT/JV5FxPhyaQUbIcSRIugEykqPqukvGxVe
/CPztQ/2HWWI49hSNasThPl+rxhvJ6mWwqfURmg+x3g71mHyvu1t7U0VQ6vDy0ig
qXuWeWjEyig33l7RwuKOxYcUy2ILuNynWdMHzNenHKQUPiVqQRnyl0FF8RRdhuvC
7vOC2w+NRBjbgX8/T9kNi/Awk20YUUZhE9tfkK2WAf5OVhthFZhpkOaytODAAtEl
zE3kISQXB0nM6P9E7J9HfMFR4v/v5gmejFxo6wUg2F7dt61w1BhQA/pQNRraCQgM
DXRcO0zT0Jh064+sxqrxqsltfB6XmR1faBKVS/hdLzpMlYStD75nHLrncABxyaT7
Dpmjn7HdtkarlLEfxwRYMScMtRrFiuN5RSXYmerFItSgcOWrPMppKI+NUWtlyunZ
bamESZcEt/mLI/pqLEyrFYFYLLt22cTN2tc9DAlKsi4yjAG/RZMwsB3c4258Weuo
dD2RT60tOUxBbSLwXQcr9A==
`protect end_protected