`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH4AluBmKIeSqQeUSJMIf4raXR6jmt0cwr66mxCVxDQZb
esnfmk2FWl+zGYLFlcMsYTDAr6K23CeQlEUkFUjrO0XIpsAPPwJL7xS4PEvbRX5W
5deft5hcpTC3nabzR4Oa3YSSc1XyZH6p7TBHiTLomXbTFIyUG6UkTR2baGwZVDLH
/KLq55WCu/hx9zrgrnRwC1bmV+GvdYWiI1jOyo3ygMzLcz2te4Dz6HQ/gwUDcMXB
uifjH7ibdAfSxGSsA3q4l/LCS5tenWhLv8lpmN+j0iiBtXK6bTsCj8wOwou/FbgV
q3iGWTifc2qxftk7Ei9SjCeMcQypAWN9mW2r9oovbQncTKMHCRiDSH/hxrm5FIti
noUOyovYmJ2awRu9+1fJ+cTeN2uGbBapDfYVNoX4mYX7kMSjQkaX9yIzAuApTJ/2
8ufPbZD9xTmfgbbfnOQVIHsu6/1zpYgcNtLoDHPNE6HDyErt95IKPWiysiK64ib9
4lq/ZZ/iscuTj9o+u3rQURzD5rxpxO4fa8Q8t+BcVEjVbhTnhg7cI3x/mGpkEKDV
9fCcgviXs/H/aIvqCWHmHpMe4loTRrwGWRwxTOCBoLs5V5hDpPC5lOxYMCTShqnC
ahQWq8DSRMExH84S4OJpZ/R+rmAxYEm8rao8Jlwy0n3T9ANQBLSwP/teHIL/1lGC
4/ptib2Y4hDbD7aUI8HPm0IsjZH6IgObmAfdeGskLsqjUD7LrfSMe3k9c3N+3xI+
WIE88b72dBWOfprk56WOl/wpcMAQUxYVRxmGmoZhzRbKcQSlFgvjTAFggddK0Nwc
9R+r1CzcLaanfy5zhIbpkP7Dqi+0Zl8JpyQhPJhpOPFBblThAum7blnbrxgUfKBW
PJaVXB6UC0SlL6Nm6FywYb5c5vxIuFlO+xjAX2VjB0zK6Dlp5Z/QcQob8EC60ulX
IHlQ9JiWyGTGMIrUty8QZH7z2T3pEFDvRoWCJ8DajcbC8CtpkmaO5p4XsijgwOj0
XlJLrpY8laskKWZL5/Y1uYlX64/R9QS6zZEB/5DqzcNhqPTQ9yX8ZK0QTLBF0rQP
Agq8GTuCENls9+Lha4f3YdKXnGLApywugsWmeyNuPhqMq5YwQw0dfT/mmj/9oL36
Tj9zKAAIyvqUVsqZ/1CeqfixXhVW72nFWRNjTR+Uf+0x0c15XWrRY7kHNPgoOazq
todKrqGKqGoYUQMhU2XEMnTpTVoh4Ns2+pRC/My7GSxjWVYsJWSnCpVF+GZm3EAZ
4c+EoqJjsApE112/xuYJ+XA2TUJ7NAfPf0XP6nl1IHCn7cM/iOo9xOT7+pFtjSLZ
WI4W/1JAohTGmt3P5XCNc8F5vxnkfvdT6/8S6utguBdV2YzcB4JdD2H3eJFgZ4tD
11pa24jASDZ+zFGThh72RccI3ME7UbPFoeYcWQoL6ll8mMbGYvA+8yA9dsuYJwAF
l9Sd9fGAC6RfGhUAJ9ijRqxr32fOQ625eaVlCqanzt4mQi+G5usqZN/A7JutKNgZ
1mhds+9KuPBUjinPBmk7vfEAw4LQU3127IIFqKLeLayIqNVY71XdI1XwTBqv6nt+
XKZSpo4OZRBeaWScS3yiiIdCz8pzLDxzvIrwvpXi5q8JdnCIBAI6uuDO8n7RMxo3
phUp7CrcFqJZeVMnSd7A8JLeA10GhoWTtN6HaHoksmXnuWieDMIURO787cY0oxJ7
jmGepr3AGJxVD9tryyokg7KJ49jhjlMKPt2mWj4eNUm1RWztJAbnvXXOGoeNDZEE
mHvDHxqm7oYt3aHHh4zgedP1VyrR+LY4Aa4K07Y2iddk84bAKbjUBJ/9juT5qWPh
+FLE+UmCqyPB2vlZeOWNv8wrDOAoB++Vm9PqBZHSB7yd9OtAXGsvbEs4O4BirZ55
vJJnUULQIgC4EbIPDM4NI/NguNofXCbZQTIwch/jrmQp1HLggv/6PyK2QnskWY18
c+DCidzYlRMq4ATA/XO/Uw/uZuT46KteS+VD2TeE32OzrnFxhSwOj8Hcn6McD8gJ
pJRQgxUPfm92kIISjzwytFvS76bMcF/Uf+SGsIfXnFjP6Oizh/8Jv+F3qoVCdJSc
Tb2p0AmGgX+sUlqHht5H6BaI9Wu2w3sfna8SSWMgGZfIT8fc+kqS56wHgkT3EUfg
/L6Qtt8ly9zEU3uGGSBl33AZpbwNCFH7T3bi6GfehCtpmWYdoMS6PntbRe1ZqsRm
FS3K1f4SquoN9PJeJSdbSdUXLEQ13Dj+Q02KgkSDB9s5SfTtpY/4z6hmKwq+xfLy
LkmxLMpboJwMcQEKGyMg7vB42hIfrydvtTh7Sy7OfeINwdyGQQdRQAlyRBa/vcXw
rMI048VX1fOBCHuGmXL659p7livb959Hx0BFmG6AlKYjk1qw2ZHdSkMt8WaaD0Nq
g/3t/1TdHlIKTlYJQA+WZQWLaBtAOE79XSqouTRWlpKv1g0Msqs9apW4AVf5u9Ap
fQ1yGg9tz1Iw8i0TibO7/7pQGqWS+VggOxAOSL6p7Fc1SVSR+mCK0Ktr2N6qmpsG
DstzjWcCPrzR3HznwGHPAmMDk3UBJkYMyk3vM5iStUPqK1wQTZCu1Dds5Ht1Yz4h
rRqpx4S3GjsLQH3bnUue3hjJhDqok5Wd+VtT1NzPbYK+VAi7ytWond2mUpU1/5J9
oDrW8V9U8x1LEGyiFD8G/K4HTBLvDqlRlKr4jSxnErbgNS9lJ71SL+YfPbDUAT1R
8XU7x0OOFH9p1gf8c4Vg2FyXHu8yNlDKjoGZx89zGC/+nwpo01jtDcs7vDKDz8D2
E4FZ0rhonwH+6O7rZ2uD/IWeCnH4/OjtVBvl69u+4jqE95wKdmLR99z/t4sg/kTB
p60Zn+UZvuvBONeKA4lEcvSVLAOAkRxX2RtRbTMMZmKrdZeXiRGI8ou2vHnm1OZN
xj//xlEgV3+PzPckCcZ6BS+pC9JeoAapXW08fhkVAuIEAjyI1G/a73nAmndL21rS
SxLo7dNyynNZKkwZRL48BGqV66/sxx1tl0omrgpO7NH1nTWUsCAGW3uaPAjxP05o
6k4el/XDQchq5wj7k1maG+i6YfdGZLHI/Q2Vh5DbRNItRLQcgALoH3G3speYsKCg
W+BpW+G0JQjXrSmpiEvk5Kq1VibS8zpeqa1JZoBtcRHqr+uENJk+25MXmCApNXhe
ulB+KZ4q4lwVDtATjpIDD1aW+IAg95es/PF49g6Bobt6uP4wARyZU6QL/QYCWIVb
Zv/gpPVIp/Ml6ji8SRJMr7rDBKJyz/75/Ry94ImRRbdvmTZtZWOu7Wz5ewRKcpmP
fFSYvDT3Bp6QxkHYWktESg6bELPKu8EqD+vZGJP3b8sdb3AMkwXBCCLwcw4Jie/1
thyl1P0QOaV7L6mzWlqh+r4MQZ4SYvZ3vhIbLDhqDc5HbYhtCzTCBza+GXBfrKrd
ZTPAGzRpWLCERc6Y6YA+NQlmtaBG5Aj/Ot7DZ2ZjxRrOKLgxgWr4i1CNDZMFbXXX
62/rgP92Nj7tuuvRCvKnEylWJDMGzV65fWGcX3VTyXx1TvfHcoweAoU/5eTyWrD6
r0EHcE0ARC7IT8B0lTjQOO+byC0AailN3tGyuF93Gan1VEwqdBqKoRBoMMjHvvI0
9KVB7knpMUnlokp8r2ehWtugt6RtITSOsK9njujehfiP09hIOW/L/aTbqrdn0vcR
Ya5eZstpOoeirnqqN3xCZCx5tQNxOBDFVrz633raQKoLMbprMfLkJiLIKicXDmz0
4lmdZddRvfvJ/aGdCuAEfMun7MS0pgzHxq2YNO40rjZGux6MhZM3cPSieDPETMvb
mLS0q3/ENbYUb5rpe30zqzSF2QzGrtzrG6MdVJHJI5yV0T5VcGAeYF3VUalgj6vX
LZ/mn9ZdsylT4IqpHontffJNLBSnCXhpOtYmE/qZO2TB9GTyDcxmzfP30kFGq0Ph
l8j1F+9pV+lca/9XYcHZ8fGVzCPl5AmfmutbohPNOt+8QT6PFwXIEWAqKXxrQkau
PDmk4ivySoBOmyS2QM4d2s2AeYeWvNAlc8kOYlhWpzRqrhpJ7JMtm25bAg0jZQOG
H6KpLNSafFQW9NdMu6nuyIEY9q/ZqYngpQ/ozMRUKSBUvXA6adZBJ3zxPdSRumUn
lySw8c8rtLfcPeaeQRzPodief+dz1ags+NeaFtv9W2Ij+XfnQHQ8mGNV+osFs+Zc
1SQcP8YLZiahxXJcPBPPFiQ3g8McaFuAsCBSlhe2ya1vGDVoHBfv7/4mB/ZTLnfF
5Us0/s/Dv8fx5EQMFI6m8MThv5oGT/rdCntq4wkLUocWfAt2+PFyVThWBJZqhkbb
tiQQEoHLxyRSGqtY92BW36P3ho1+vLAQbtqcsQs4TlyEoPPvXCMidDM+94epuid2
lsERt1hwYT0rMIWf9qt8yAr6yvYu5/f39tXm0v9PVvcXDU2gnrzB4kmQSk0n8i0t
RPlbkHFHi14AR5FtLCYSLcMfizqkOx+djCGD2ay6AkLXPQkqoi1Nc/gB40ZzTHrF
iVSADQRW+gRHrnV+2syvR0sEsjcdP6raViwWRp83nlAoiYG4WZvpV7/7IvDMcfbm
qeIX5vf1tXS6rv2yP/uFWnovPGXD6KjiETsGcVfMWk2EITy04Qe+v0QY6Zx1kpir
dGUWf5U64QHB/LEdBvy7ERD6TNDKTIzbFe4iWnZ5IQ604oiDhTnaxLlpaZn6jGos
1gskDvRJc82JdT5TIcsNbGRbYfXQte0YLGqsmU2E6HOglZvdHV6AfHS26gEVZEOj
I32jt2YNvjSY5aNaU48VxzJ+yeqF8P/A2eBNsc3j3ACAbm9fC2UZu4uXGwcPu/gx
MNeVxwZ5JsvOAlIyhWmkoN+ppMLhSdB/FDYbVhcpbvZtHBNzZKRHGiXeCsdxiC8u
exlhyolLWUWFxTzcxP/Dtr3JH28Iv/uxKCUHB/YUghfsyqS6vffqipsKc1rX4Iy8
fcY5/vIP+MBypGd5m702udWRnQCp7VwwTIiEzbyzS/10bZ+kaFg/+zkEiKvZvKfm
ay8XIvRjNn4d/xm7Tg64+ERIoa5bVyDFuWH1jCbxoX0q+fmq4Bvr+W1T1Y27lXbr
1eXVbOZ4e8Kmd9bDzJ9B085VXqwEwc+fi7WsluwLiB6RUTr+PjXYYrd5+VSl6P49
038ijmRKfcPZVLrBpBzMpnUWAexyY4uyOqxW0Vq5l13wRrsW9qf7VLZ5TmR0RIEW
928Riw7u86WoIatV8dMMSIpZA3cnZnEFpgU4OaLgA4I/PYVRIcV8MXmmH/yB4O9i
V2UpkMnwvTyuuqpUjKazPo1GCya+ZFYpM/PyNuAuy1qSzV5hs/LefL/txENgTozR
dZUs0PV2omi3I8ISRW+B0dhK7JJvS9NwTvc20JFbeSVqebNPXmXxR/wTYrXmu+8c
bYlrpAV+P+WgRsxMjJtOkapmb0g/ZVDwjAu+Tw9cHUbaeKi3f63O7m+8BYxuaGp3
XqzmCnuORlXFW2jOtO4P8qh0bbM6pijCTANUIEMG7/TzTAo5KdUeHAWU0uDa4LWn
4PdaimP4RNAArWKn1IGo7hbz+8/ZqGrKRXAJvWFIZWAqIzApQpw0QCwRCUPo0KVc
8YF7BdED7Gu4CbXZJNokkhZCL/ue6sRPmVeNM5q0Z4CWIEKhyvNezdn1yW4Vh43N
J0FSK0riCETs2i+VXAGgTSvV7vwX4dXG2Bs+ZoD1XF32zyggkCH6LzaaLi9lRGnS
BQwRXlSdmTeUEPB3ni2lpKR0HHGxD/akPLmbuP7GiYuucJdovFJquuSsxshjnJBL
wIldvBFs2EcLJnc2lLAD34tDg8eybfJ3oOvnnNLoC1WddDiejBPfY0O/8tp3LHFC
E5ZcfnnGJf9c4tM2CMmeYz/UqBYyD7eKXLU/Kl3BFH+BH0BHtECsRHcLgHibDGRU
qFVlN+H3najwTX38vvCPCoOvjgYUqSzrfg/AkzdJJgMZqp12UEZL8HXXm1w2Ofol
ry2HyLQ/QlWKfpMVRZciyEt5rz3geYPao0onSJ+PVYMHrgTDbyVCRIdII3sgnoEk
PTV3q5Hv/pVOk8Geamq/aKOVop877VvqZCtu0vIhcFsDJbXEWm3WSju1PF4f1Lfy
oWinjPZHuZKvDy/o196iR2MRs0o1HJPqjG1C5sGeMojowyrC3u7j/FoKQcx2QxzI
yTeMqnANvCvrW9D/5uIJ0MG9NLOkRRDo4n3HStLvd48gIyhygXhw3k5DXG+EUubJ
ab5i9XX5QFgkgsdZQcTC28Sjf5+3L6/cGGloycV9mmMaiG/gG4mOX7tTtLDEt99D
7w3LsZHev1jins0T/M4MQNKEEBot1ZN3nq7R6rEE869Aarb0NpZH+kvsQIuqTiF+
bG9xiE3gPZT+BgmkgpGKWE9Rba07zJh/HKK0IqEPX1OKa4a6r5ZG3Y6nG9y34/lf
jYRa5mAe/LXFb18B+EuQgVv2gCN9Wx+yOhRAyts1vjjO26v9LCnNGJiylvO2fRiV
XAYC6ekZYiCr63FFmMK0rIR1JybmNf0iQefXNspZIkgdyMUeq2Y6psnRCHpHF6Fe
+uyL+KJjyg2r/A0ibBwHpLaMuX1sB6xfyil9GmRPfPlKiC28/aCnyZPV20dy1g9M
Zag2UkZYl2Tl4Id4J///Vu3ZF3owySFLjRsQD/GI4kkQ3fd0Ip+5fI9kD04WlCuO
9QG3qTJLEsgbjy0e2OVCs6dUWKaXgfSdDKpCUkbbOZ2uXI4Y65Ki9rjAFYnCZ7FS
6KLnFy/xRl8HKQNzEzieHLSnozAASQb6poBbQRvsRnVFAKpa8Y9B6lDGBLE1TH9T
lENrgaCh0++cd8zO6ufRL6tpTI3Nm4Zh+aMcpuqeHRrBK1nWnl1kt5dw6AlTWSvp
I599I4OKSh9w7W9yU8x9dJgdCitFe7k99lcVmobfCISj2pRGR66o2VjmxwuqmuZe
ZzdKMWKoCERmtRHjKcC5wxFQQzTdup/JGb/kJhWaaPbYhjiMxgcnJJs7ZTO+Mubs
nGzhzWnA3YIfgEe2tgBkYRA3O/wEYwgEiRJhR7XmoIztwQl5ztuDJBY+Ad1laCRX
1tK/30N1SuW+BZ9/FsK6tAdG1shreJKRkRk5nAFVTZEdwdu/aOQuROut1Q7dFHXw
2ftIgK1T/4HS1U906YBJ8XPWpls5hd4qUfHxbJC1vrA7goV+lOSmQztsavnmE0FR
LrwT6wV17Bf5CdcVzcLWqIlqYUttwCsGpWHhYdDnQEklV1fBs/QZo43Mj8seve/r
RO2RZfrql7C86uccjakMoZETHf9+fJ7EDKmVi0Uc3eMuJDBM0O6Me90DRX38tiPo
39mZVKxhpw1wQHsDtQJIlOnOpLhru9EWeEWvv+cyDZOMYeiPlXN/miDKP0Rfs1KU
0xb4Rvtyf1OPyHWOdoFm6b3Z/cE1BYiq/fvmJTOfz5tVpIK0kZ+0kPfKtMoTQd+G
qJ0t8N1W7AC+jZ7mHdEiM5xWPBfjlB6tWjOpnv3/eVTkiO1OjUkpZluqlQ4oACsP
2Fi5SEeelGZdf6qBfOgKpSZ6wwSynR3Xv3oUhnDQplRIq8ExlNASaaUgXZdDBqmh
FoSkov5Op/qOAxazohnfj6kyzkNTDk+mjS5AZeOubA7EziQAtX117MRPOse9nvY9
rYJU5ghcDjIt3/01E/qit8eaxxyeam2uAQo1JaEPrOc9WA8SplASVHHjf5vHnEIo
FUhk0PQNbqhLagTYstIvJKwvRHMiC1OgLDeGPJ0d7TrGNJXnXXVErEK+dP9kKqLz
D2Lx6ZfcbLFkoQ5z/0prmtplQBQQuTNP3kagS2nKSlMU4q7WMMFf61le6U9ccQB9
506dW45Sry2ZfCG0yE0qjV48ZlsmRT13I+CJSMsdseuPGYRyIVEx75uwNhYDDlQF
NGrM6nFTK6HE5LU+vupGjXtoCtV4hxZAAd0QyLIFb3NqozAGMkvC2MSxgH7ODGmE
13Ds4wzFHLsALaQljtx8kxjb8cBuIrlc8ZIkUGxf6OQW+RoUb8p3c8+Bi6RSY3A6
xzV0ZWBkd2xQS1aQ+NPqxslzJzoOALA/glvYc2yYDqDseCrLIL8eUu3by6aKecL/
jcdVJcFcEhMywXxGrBtrlQFmD0xTBXSAag//JLc8W/peGD2acvQD3knYWxSBn921
foS4QInrj/KDaVwU155qb0tjmH/35nEAnkzlo0IDDKAtitcMn0Vg6u/DZlabE2nw
NhDTqNn5SDO/UO4KJL1NfpbZTYBOuB9sGbOSa+86r51eu7f5QktLsjlX41+7wlpn
Z1pEDWytdkdnmc6/O8eAT04mBWKu5/hU2Mw3JAQx02uIyCZL479ZgBX7RIE87D+W
GC9vxt/jEkcx1WXvayqghQYJWNsn6VjWeL3LF2BGgId7fFY0jPEVOn/FLIDudpJd
F7OT5eOBCNE6rpXU1FBWGabvgNruggieLYGpjrQLAeE7KUobFDwlbt7XAQ2ozqyk
S1cdaLiInfIHzyBUlWqney0Oz0/XD/Yv5lRN84mch27K8IvzrFm7JkxlDJqyRZ3I
BB0JudxoQHRMuFuo3jrZimujFU/Q6zfuwrc5d7qvouLv9BladlGUtZzp1n8iGv2b
R+l7ryC4W/QL19e5f8kcPJidxXrBMZLRkx61VDN4+Pthba83rzcwSVq3fYuNu7W7
qRPivkSpaIiWZWjtO/YYczg08Ah/CxhmGhZl1x66qe8C7s9xI7IHDAS2fdX+LQ6N
rudKlLj8ecqpdJVGHu4XlH0jb9MKmuvB4kv8NUOnAeLfeXU2scbKcLTbiKlvn435
/qCsBELH45WyuDOqE/H3kPVkCtWyZBVq56RMUG0M4swMBR2zg6+x3TWeOvhVFUQu
vDZi+SyiyPoY7WhOhQqxNV+eVW2tiZup+Qzd7hTGhBL5TFaPzcUkAGp2Cm9cEmUb
Sl651JychkWcrpUcNAXs2U0T5cMP65aBoERMmVcdNm0QDBH+8pl+rcQIs8w7fsp3
GfNRIrG9lnmE3p/pdSDqNgDyhE7SUlVOhbERTwVfIYNut06vdugpIL1/ZPbB2GYU
72QCv1u0F8iP3K8bL69pDSxm1/YFjJZJ9OHUdqfW/jqCi5JCnS1T0Ic3o2JbwOMi
94kCQPWvYD8L0D6UwzHmL3JGjiYgkBhvqPI4Sg12PpwTZiSA1Ltdbrl15hroJhp6
2sAjkOqYmXFSj9/6pVOrXFQH6xm3iUnb4Y5T3Ok5dtL6EAUwkstzPYzt19cGgK+V
Zmxqg+V4Vkl0YakIDAYmhzCuQQwCOeCLgrHGD9jc5zlaZfHjEvOEzHHB9QMaEVN/
4wBhU43WpwWruYvt4esXN/VTE0HphPg+ZK6b0oLyi9ZgcYYQS9113qn+zzP5FNP6
tehCdwhaxxzudUiXSukOOMnTSCFv5vMImC4rByKgtiF6Q2qJKfo+s8hn+OGvW/h8
FPHtyLvtPeTYGN94yNcB9nivztxgoidRGM4lwnJ4ce3BFXQ4FI4zSJJFECZYzvKS
b2MZo20ekHRkN/6SBnvy00uRm48B64fwABku/KZ8V78OLhv5H4BT+8v6EObwvZ8i
KW39TM2ujr0I5mjUTA2DQ2zq2zEXmh06B5a/V2HtXc7yIpGB8p+PBLldtkPIbUAH
DFHDB1gMC2nE1JVpehqLjLXWhcpWakH9iElzTC1nh1PQXIWEPggufZv0eVZ0bah2
oTm3caqCnAYQ0I1JHomQO499LTk8NTaAFjlamw7725buKSRZE0jrn3iHSgcNFE2R
KN0XSg0M7vtoklYBnS9OB619UoPHdVzglhhP7rQgmpRcgrTus0ns0azQjnsq+MQk
/WUckK6bq8z37u5i1yYhh1g7UtNxVgor9/TqKUHCLoHCIvegVE52mAGQastWxNVk
x1wMM6ZJUHBbmn2Pa1MNweT0MjgwFT1GtkhXAudnE+Yc8aN+Y3aZOGAfoMezoqzk
dT97hbySMmV4zdyisJdAUhfhU5ytGsePU+Vjt85KOPFZUDpyQn07Dd9J1rE9iz/b
nasz+2vUutn3JJItwQZsixCslWc4vr0vktaxFvAn0BMFo9fAYHGMIyQqxEHFo+cn
0U6gjEV1NuSYOsFN6zUpE52t+Vpprj4NXTH7TgPQv9HqYintt8HKft5eqYypkF05
jgQAzoGd31CFaSb+A2tSyE1k582Ylt9tvZsJESXLRT22fwZfC8M+HqILoc9wMneX
NRn2gTjcRMyVvyEw6yrrpQsyne0EelWOiBd0urFfAgKt7RC2YCjciseuY8gXA45H
cFfyzubGv/T0YYBFSl/k/0FRDbPe4H1q/GlVncdeh3NJLnEzokrfyLQf/kGXs+tG
egdvi2aJDOADpOqPNpmMLQTnMOqjUoL7MdUHd96Uu415bl7+WXAbdPtB9BoEdQ4+
yCZchlNZN60zAw/qnU+dOJtiixxpLZgjBlXvC4QDsbakElr3N61p90oso01ZC4W8
srnlzw7NXsQKqJOxEoPTPwAWjgTpTvCm0eSbzCtrQGoFSNTRmLtt9x5coigXkePd
Q2hbZfz9sU9euFUG1sZ5sW/VWLp0CEqC1Eke3lCqIHe4btG0Mvr41WBKYjnK7/hT
IDtYbo0OxdVRW0zS4qGY3QvFw+mQ+gs7l36oGdefK6ROptkkpnEKpC2EPWbp89QZ
tW4kgrLmbZ65lvB6MrkwArYde6nveqTHLWJw6vKaWaHWdB4eXfFcXXQkvB4q2M5y
/n77HpOfCbsNSE9a9twvtsmLtJh1ZtIr18esABzsAJT4GEp4gwltxW3q2t8TDdUL
nEGCBB+qJw+gqpF4SAaed9YioVrVvjFxEX7+75/Efyh1ff/kJb0NN3FgtHyun++r
NbFb0X2M2SF58+f5Vym5K0HX2wzqDRd/A4YJZvo6o6rXSZdhBa6X3d50kSIjcRFU
dhvN1Cf8gwIbIcBDh3mrkNxdWNkSQyyy8JuV87YJdcmA3EXtvMLB0VSoPICx+6Kx
xeKMaKZmGGgXSbHqS+m1rjOBXBEo+7L/D5FWJk0+WWWZc/wFiyZqRG+HQI+sWwsF
7kHHrYKXIczGPh09IFmlMJePC2fC1LkriFLbmRvt30gzfOoEHVEI0pvu1JxRs6lQ
XwKaDVwsbkY3S4m64WEIfqkBd8SG3KoxL1j88OmxB1CxxiCW8aZGirk0GfaMPmN4
/zrVX6FsxxFZWqPblVi9e+j8/VNppbXIK5y3lDYFHJLgkq61HaKUE/JVXsIHnWwh
mcdaxeYqqG6MX0VMufYVHzfLpzmttlMOWazMo5Rchx3qL32TDo9GUQnNhVw5cldD
2gqsR5RIHRDt+6t2/40ZUrgRz5MeCYznc90ajyEtneNsdjEx/i8nJKW53ht0ktvS
qexrb9f1kunuE5njlZXx14gKenVnqeVVZvL8ZqwsP7MZjxXF4EhNktB0fA/rnSnj
U4T8WJ5wTIFqk0FYWEfaghP7p+2UNOyw4uEKSnmNtjALfRgAiF2kV/XNKiJ402I0
CPgkhoIMvejYmfmsBedJ6zc2QChd4u4TcMYPy6IYgP8xSr5psk8+HrxTgFnfwjrq
KO3FP1PFjm8o0zcKMkTN7Hgl6Usub5+suL5gdZdaW1YWzdErqAZP0TJeZ3ElaNS+
2OVtvKrzFbwIJqSEimu7S6dXQa/otQDBcGkExbaYKK7x5EzyabeklZeQZxYvOt0F
6iJ/rtWY0BfBrxEb1Y5w2DQpbpGmSLCffSVb+0qKmJHiw/b4Q5H4prPHPtFCsw0O
kS+K3TMsPqV33aaNf1LxgyowT/Qc1z1jqu6MaQ7Jf6r6SVdIwhtLJIT9AIJDOPyI
JD5RO8A/3wBiEEMNq+vTyHvK1hPybQONIILKxkB9yPU0Yt6QnungBjts4A3YH5FS
6dZI/PspRgeHcg3KR4NfrkE8QW7JJKc5q6pB48bMcHLsBXItL+A9b1uglxDwByFL
l6ld7SRB6kRq1YSkGSngQCY1t6kcmmB5pJ69ejmqzNS42Gbdi/idZHeSmZt4aTAi
8vnIlIYQYlSSFqyeLAwtC6KoKXzr77K7bmmUTnCEe0Xx9AKtezLwAXkJvRjL6eS2
2qj3aMd8os803emgKuqwktMo1Rbojf0WxA36zL4cdMta8OtMM0WpmgyrtsCvRFji
L7j7q3UNzWvJhE3sXYZxCWttkO2ne1pXjRmQLzoUYbMY8EBVxk0YUe3zkbrk7BxR
rlT5IAa9BTsn8C3diJKRae67Z7iMiIUVNo4xGrXFP4gKjX/dBEystFrG5oqWOAAI
95nVJSgSL412nUF0fk5wcN0qfWtv+OtlbJ9/AQUFGxia8oCgT+KSgqgadbG6SUqy
NePlKs45fNJ2+iad71VQYMPWhWwmNFyiE+0m8GCCxUkKIFcYcQNarHAe1N0kVHRp
kqKHK/mhuyqWe4qfmSD4qji3b+/F+HIMQgMdao+bA1HCcxCLPiXogHD4CSzsSIds
hmf8csJgin6hiWMgcMfP1NXFvWAJR5eJ1nKlW94196SUZUlfD6Kz75TanFYCqS/H
/b+lIgMVBxqQBner1MSUB0CKPhk6yb4EI6l66hMSxYonsmdz7sb5QXxVVdYmNi5z
pg+cr2GxbP+JBYHpoqFgcXEvHx5WJr891vOIk7s86nuF8hKChO6HnP2yee5eelSp
ZdU331pyh4bdx4eYt4kf1NhkoSFNBQgQXIEM+ctyJGpFL0NC+gAa7+aH2OiC+tLD
D+iT71tL7x8ETNnN5AzpxXXzi+AmrJ6u6HztHcWhmM8O+2UNQ6tZk4QArQzWRC8s
y3BBpft/GMdJJ3D0FVE8kZCq3iV0ps+kItZ3DOrL5LZG59FsA5Oz0kAVz2KxFHhl
tL6xksd7ChKlnZ1qntSVDsR1PgFf3tn/bZH97OHYhkM8BcTMVNYCTFCnaCRaMagh
DVLdME1DZYLYqSMAlfbNE4g7wk6gM9dVOKP6Fw/C/ntltm3LeczSuGeFtN8snXhL
RtzKmwZzyu0UpYkRRzWaOOdWvoz/1oGJW6qFooDONvfu35s8RNfgaDJjCvrXhADA
5gDfRN3I/Cjn55N/CublwFvN/rZJsIDDnZRUmNnxLTdfMCiB1y+0w/EUcLlJGlz8
kzNxfjTilfRxgOWVmTDpWZunGYCTPOnGbwE0R7UXMfC20JNVUlnUoumGA7rkUOhd
hvxJPRyrPuU5Fk/QeP0W49bqbzO8QHKYFebdgcyITGMkYELvsNTZ2lBLlAs4ukwq
ABGIZdBXAlpNbMW1/gXfr6Ko+R6hoSSyYWSaQHV9l3fiIpTJaY4bVhNvFI+tiTZ2
oOo9OetPvYNuQ8iO19TgZrhj3j6MZC7zdpq5uPtMwrPxGMw11G7EY/YnGjZ4fASA
G/mkoWanAcTFnJkVFqpWEgNHdAwncZ2q6j8eP985RwM0I/3tkD0rX3QtYH77S+O4
dmJlfiom4e4UJwltlNhBi3zB7P1Ojm8vbV5pCdV2vkVdmXGd6Svmct+HJNzoN7U9
wqNsltmSwFJ/BhyYsGdPzVvbyEl93pGOkU9ei/OWCwfl2pK9PnQ7DMZoe8dwdQKE
TQ/wpSVmdrA7y2QkisaRbTsJRHqJLMj99bFw2MOUS6TU6mlVIxoVnXZn3wMqeEHR
8Ib5J7N12z39JTAVVIrxu/N0JSHXKPQhp+z8C5P9xmuFTK0xD3eQ38l246LnVIl2
JVuN7OWKdQ7CEV2zoZUALJbugunqLfNqdNAA7D3V6xq4xVXFxWce08ROR1x0Xsu6
Q6b77DtIfBMBhmpYPLJCA0R9GKGIdKXCC0Yi1EoGE1IvdBIC3uUTUaRIi2yP//EM
wmny9WQViRGy6SAYuqaQDzZvgXk4Bkwa/rH0oCA7TbDAwhGhfoAWuzmGZ1rMtp5x
xPulBs+iL6T0ttDSuOyTv11ChnSDC/D8ZOzqwO2xzpzCZNrtqFJtEMqhyy9ffHKi
SuASXROkYzES5daKLVxlCox29OGAtt6Sx7/cm0yO9I1x+xUlRVl5+aUQyXSNrrPt
Qs/TvR+CTHZmjkVuACBfglfPXRARtmIqHodzrKZR+SHu9JSCa84WjIW/YJ6QXxGd
QOKZukNeYz7JmC8LaBIv5WijrXauayveKBGOHSEGdq1dFtheyHl6OVAuE00dt0bG
XxW7hGmyeado2hCSyu5ot1y6+0QC/54dlHNcaCaX8SZV0I1DdtQW9MI3eQ1+dnGT
t6Cvt2P+1XCVFayBWBm7WWYPMzKXFNVDhDe+hVNL6aBJRsdsoGNypktXHNEU+bVj
Xd6LnNFQiptWZmuH7QGFta6BgzcQ/jDrtVTiW/R3ajMGXqp84mM89aNqFb8Kflzj
TJ6ZV+EKnhqJHz2HVZx1ycmeoHQRx9TKlki+k9kXaT5AlhQivsNK/eaGBK2BGI0H
3NeVTLHTv4gQ7R55jcLsfzxcDvDxV8FOaLvnNy2e6HK0w4CCDn2XudMX1BNdtB0U
h03vyhuozx9MhvRlya7YU1Q3//vw7wymB1buZD3Tpz8p0k3/IA8fA6eKXQfPMWsO
JIvhfEAaWLksExjH2DDQE2MF9F34FWktflLB2h7KplOPIZzjm9VIASa/dI6ZDMl1
Xk+E2Eu0K0Tm5CAfVWuAsOn/N/DAf9X1L7zazDSBt+MLTxOzNqoB3WHMIPatxuHr
ZbPSIh1Wtxuarc9J4yjMZ0hNsdWjpE6BbvPLKDgVZ4dUeM1xo0S7wyStxg1znYJc
5idh1RX4bANOy0jZ8Cp3M7nTKitrNEeZ91RvJOp0PdcWQ4yqS/cglcF+gpsU9Hbj
J24s/a8w/Jy3Nu1kSQGOItJUtfetNlzrUnda3D4E2XxBhtwe1ZGPMKDtDTZk/mDt
fn15AxGRVOQ0IOSfE0rM9xz3RiO+uxlxn+4bMry7+6PUABjFKHiZbEbBaB2PTfIu
A6O3yQ0PlAPLfHkjPB/oL72ZVS+4bVLpfGIV/SHUFQHyH8y//ods/Pf3nDR465au
4urdKGkQ1n/KGEQhxw3WLPfheuH5ZnG7i3QMHPvvoNp6WYSM3H8hc/c9spDQ2E12
ki/i3yxFpvyjOgveFuXBmvdSHd/dnEQfJGs3pzdnY42uUsl85HM/LLvaAA1vsgd7
0H2ytkc+/npcOHqy3YdOSeZduGCHOPvDwbqPUwocw8WUy+4iIw3crdZpe1qxLEoC
yCrPvrmwZqjTixYV4u40PvKYmJ4kBMHVkOswyBKoopSxM2WltZN/EocGCmLB+PNP
8vZsZEwd7IsaWPcemtm1nPl64VUzfrIADlleQARNoo4Ixb2o3qkTh+7x8Gvuug5Z
63KnEPmQ5Co6c38PeZzjyMszETsHry2/DcchA3chZ8rQe6Q9ZT+Im2ndtA0ZKTFR
3/b6J6EyLN0xiXKA5lAfrM6JX/o9ChWWn7GekTXLlpF6qozwJAamd/TQUtDmwqLI
C6Ck1EvoWU6ogVPnEfUq8H3qjoOJBmweOhGYqAcGx5QOhs4SNC4vRUtzMtdEYWad
1SjQdT4RpdJnkSDsAUzRw7oq+CC8Y1+9XbatmROrsfnMs79wldgzE7bAEfVZfXbH
ycRjhwfmeSL7JLbQw6PreMcKwj6PJtikDsXbF1S2FzcaD+cIlCYUkfNDgWV5izhY
+hal1XGwLkYpprVnE+Jr1vsl7/w7+DcetHCF1aY72GbzVH+5yOa8KpGkWl7cQWxt
D5Val/B+AttR2slmAUE//b6LWp1wM4Ml5ioMy+BXxHJzfRb3TTyW/50krG8201Ky
/BeEykLCVaCXMFZVUfS+nSaHRaKgdzsZDyXqGQ4itdf6mpjz0MkmS2RslpeJMg2j
IX8t6BVo+gWkM2Lo7x0mexyFx3s2xVCUq11d3UTxJUMV4ot5nN+zOsXlS+QXWCOi
L+XOi2CPABd3sikYEBzwdnYKW35fNbbUxSQpsC3X0zZWoQY+/J6y7SMUdkd+SKdc
WjXLQ1JVX3Y39qAKUkc686dwevBM07/r+A4pxZ+XPlucjC3R9uZvPQyqp60AZB6y
1eG5QyuDTZqEthvIUEWoRdFWk6cf+A6rnl6NRsDLWEJPK8ar8Zh5qFJsrqU1tX7q
N0O29NNc4AnlCTh4fl82MvnnuayWlG453LhE/CFPzSC7pW/UrPEdSqO8rHYeHHBQ
5/j19dMkti+YS86w9LDPLIROELGAi4wDmTrYhyy4JxJ5jFF08uK3pCAI/POorSMe
UNR1mBwZfYYS8VzatTSHYiDeKQhc6sXpcSAcsDLKm1yRUe07SOc9bJ9xTEAu0eoF
r3l2G3ut0DCuZiA1QNUqK3V05uXVHPAMEsaDSpHD6BqM85LRvPBfTnQ5P4a9VNai
cNwMWDXYr8k/ID9cMbcWau5mtSZ6c/sEXBGeM5NzREXHhlUe8rIHWHml2Ee8Wui1
Ezz6sMInjHwzf+3mK+XWqaPwEe/aa9A+dB/qpVCTyJuG0DVoYJ3qCGAik+q6zcYm
cvLNQI/gbvt9JhvJNSxUVMQyXVty+A8vXZmSjutR3xvssg82nvulD8IIDeqoIN30
dq4dXPn+/25Bn3Jb/nCgi33KgjXmrZ7GOu4o7ZldufYFq0a73hgpIuKRHChNakGN
0+zIxo1XD0Sol+1AIt/utBucMqCEOQsFKNSYIWCPLlnqQHzx0PvWv1BQo/Oq2eIf
Vr+V9yaojU5R3+NL+f69eHvh1g3tlI+OD9VPy6QF6/d8OpCrH7QrHwkscFO6x+2w
Pe+W3SBgkhMhazkm6UegjP8TwvYnsCayJExK1IS8Y7sbI+bmFfViULrSsVm2FCaW
iWikk/uh6PzjYFNGpYAiJzh2U7etx/bfCd0A2o8CPlrJO3CabEUFbz6DPWvIsRmh
dRJjOg4jJEzKSzttIRC+SWpPVMdmOLhl1HxacEjttK09+LdUK4t9gclaOOJc+T5u
oeOH0REfwsQ6ntj36CRVnTpQEKR6Jh2KpRKFMiGpt65VlSms2rgiYH883Ihf9uw9
bqX5J5kvWSp4Fp+7EOSEVoe8xeqkC1znOOMClc2BmO/Isxd0+AtOho7n0/jNTPjS
dh934ZmN+LzFD6dwZpdjWQLxE9RA07T+hEePPUTXj0Jqrjlri8sd+2hxUgTeW07R
dKIApBepPyclZHuEDgimHb0cDhPAuiJkJr9ZcicS4ffyLXnv1p6ID+ydlklJdcsX
PdFU8yYmDOEn4w4DKvbqLtQwX0CINBwTNMcqpsTNpydJAgiploQFx4OOaSaAnhg+
oL93i7CvSn5RUdeteRCm7SrCYRo1yNUEKkotkKZoc/u5khtnENrMGQzmhaSDDL6U
XDHoCWae1Fw6fkm/WZg3dOH5TdMV02jgbk2K5ESdjwdUycJJQbjxTHeWjGuV/Dvb
0i/udMTX9oQLDa/wQwdm/tRAvoZ8sErHH2fi4gi0hNOsFcWE9XwlNVyeiQg6Zvfq
tDlJiYe8fcAyt0cV3BQ8xLZNqvnfylEmW7VTIu0BPJ5CaScygqfpHq+1rMblfN9m
HpgRHiAGFUmVW5mnEB3QZPJpUmfaCAPQzr7H+9QjzWUmsU57wpWYMtcfvQNLFX8R
r5WsAjPwG2ZKZF51g49UkBss55+BdSvRxQa+uTBmvWjWEarCKQFYJa2pILC8WwOQ
99Bo35O4yY/OQ0qpn9b2dNZMrRHwj+J3KK7BiVDJ6HIEFEgqAKfQemucAxuXAZJP
xUfFvLrv+QHZMMi73nYZGQD4QSwgwFmgLQ+bVijdMxd+lEyRU1sUXLVbDyJ1eeil
8RYP0vxh1c2+R+ubRAcPdMjNQOULO3m/UVWkDBK3t+uCFBEfJWdERqm8v253yOS8
rmJ+CB/gURfQSdz/FL9fwRvcbShVHGVqdPY7nBbiKzhNECi1SlgC2zibuT22uu7w
FUNwfuHVGlni3xmbjR0nTqsQPXrLu8/YSuzvrsLTHpam3x7s0cszdJUTuSe3hl2I
aLrLzLCbg7L41MgVhHkvor5azwn/k65Dm8/No0HrqA4EiX7AIvwOwGJSwjD+vhzR
fmgTTfz4ZiCdTQhfqiRTKSseYSSg3Y7fZsVDVH9CCAnVUrOrEu25Db+O/vPTVbbx
sRtZeLDCBztxfSf2eudQcvoTSDT+f9FvpD931iOIXSBfP45pWD+tnR67oFo/fExZ
ul8KrT75a+GbDWYLlK6nuL5JD4QqxEAkFcjQuGxjErNuGdOkMFXL8DzqyT0mrWCi
dEypO48IT9NPj/MrLKq18VTD2LVdlzB8ehM5pPbcAa0vOJCAwh5Jtl7QiKzvlqDA
mPW4lwgWbymbntuwPU51LAUa/jC/SBl03VcwO1bfHK+FwDFTbdPaR19l25Lcvpmz
pGoYNk7BOtuTrBQ2fvacTbowAXFjti8juKreSuanHTdwKHbyb2au8KJYCb3bAcbq
L4xxrOKg09O/VF+AXNs98TQCimpq/15giSBQ5lKe2EqWryLVYglirWDynJqL2Hz7
yNnMQFIP3N47GQhAJSzOYBwTa5MeCWN19J5v0ioXmvvGvY9x1G27ycoiafTxMW0A
65ELOgmhyAULqmep9zPDIwcRRiwIhjrC+ofLd+YuP6JoPdjD9473AXTsrU1GmQsO
3ozro77oXdYKUQyB6/oWT2U8IkJ8M8GeMRItkNf+J5CR+rP+3onA/+dfHO6lbErC
JxSFmdwUlwauHTaiD8L7jzh4r86uLqXJN3Ou3kyQTizS7HwcM7x7BBHmeCFn4Pew
koTz3StSlK+wIVUqJAzrXDwm7UyoPMq9BOxklVtHolyqo2oh9gF6CqQC1G5OFgQr
vSeX5TWRK3YlYi8pqcdTdNnn9RYZr6TN39PFJFKEIAk5tVUFvRVvg1uE7Id+vpex
Eck1HzhTp4idMCOgnVVs3ggylp0PR5f68qf3ry2pn5AXquPRpKea8FpiWAofPvS7
+W87NGN4nj3SJfjkjE2UfcogSktLDm04OqWCScJ8SPAf1j/gWFZguC869EbT1knI
GAQluKoLASNBLkHmUk4gYlvfBCzl05hd/L0HBXIdq9x8UFX3dZU0+ZxpfVAwrjQJ
HuRIA5qkhm6D5OqnqvgT8+l/kWmOdDP6/C/Uq5ZUIh1MCWTChEvtDCIvvnNIj10u
MO8EBZHr5EfqQ8K23IqnNEBVVDsAXtg1dhMJIPbf6uaa6TkUJNTZOVfM00DLk8XM
MbBIOrBxdC9PQcYvxzGZt0Zygf8pbfQkQfa7JfmZmXpCrz/DNq07OHItwL59+4DO
tUDRRH6G96xmGb3dRKBCo87fYxpQ5ehxnR5XrgSL244COdLaUBi02enPF9+sw11Y
1IWAm0z1i8SR0S4ijRHmcR0Gp+CaGpt6HBe7w8Gyaf5N651a6tORT2puxT4wn8TE
OTsH8WCr3+7nS3vkApuhhw6f5+h7tNq0Zjf+0JWP4tqOS/xhCfnUzEyF2pdckVSA
riD5o7CFyzjQ8U/Ca+J6M/Gn6I6BuBkjOKnUXi4a383Y54z/nxkrIrsuUvxuiepG
Pbb0VJMsIN5hcjhXze31+RCj99CgP2de3lR037dAszglv7FBXSe8itPArp2cS1ia
G2TW24c0VkgaIyfoLgndLXiXFMoEYGodLDMSdn1SadJXAoN0nUbzQcjyGNPO7YxM
E4C26Xz0EeZEakz5f5hTOXgpliZjS7n/gpYFYEzUIenQWxeVH+FHVnR+xqa4exAb
r1z+6hXW9Yaqkb1BqjGPJoJJb4MGG8HXKSZoOptsRrHk6ng7HkDtTruq9R1uaq2G
arszOR6snkk6TCrp7v82vuJklHT3uFf+mjfTx5bwnlnWYFtjnro01oMd3+xj8qzA
HfHSRkM0gzeyiiWdSn50dFzcLGpfOMKcvUR/e/zpO561thEcjiT017R6OBaBZZ6U
YrU8JiknFfC3I+xdwsb+5DNlnotsGGNSm64sB6YjJw9k2KbFnjtKyUgHXCZv/SHK
e9aCTINqv5jDFslPwGs6vBVkhjyOFDMIvuKr0xf+TDBg5SuSedp5CmkwCwq8x7cW
raLPUMG1ucVnFhd2OVroGcdyLtAMKd+o9tlI3qLGCaR9vWxhz52IY4L5CVoDHe5P
lCNmNqm/uw4VPWmHImK+hE9R9Uy6kX6zUznlCASYVW4/nYM/yYl5IKymYtXCrAk8
c0O8M99WJJIfyYNyHDqoRNOKV1jWyDocteZQGLl6YF9sQcAeLPdHcqVGLKgvFrUu
23jeDA11FHR5Lzp8K9vFjVcVL0Xu9b4cFwrKzTwFmyX0Zy/ppYP85jJHPs4PuwJo
0ZGFB08r5eufU9Fevmk/Tjk9cHD7TyDuWLfs1qCINa16E8ypCCTZRVs7vVKVgO0w
VQartMBfmnVc76vCR0iaZqBT+99038fzf977B9a5sly6z43X0vS/QRnxfajvdtqQ
AirMuhCIoULIn2C+XY0BdB/5/8g9Qh/vMvo7HQk/vtmnLC3cd1MYABlDpdhUCAXO
WuUieoJv7W9kClJWRE0yvaquDkbwyx/B3LwpfKXKzQN44/KWGl0wXKEmtAhe0XKr
8pyrV62KFrT7zvBGEuoMjGqAa2tAY0cZbkWpSkJYu0SAXDygyW9ptSKRKWfy08tO
G3ktJwb3SOCZSbgVYXwmg26eWbMl9PyfGp3GaJSk0KmzC6n6zzB1OInhoEmS8uoO
S8dH2WZWKiR/P6CWi6v3hqb9M3m0IDsx8ILZCn6UCQQoCc2XvN6Hp26a35JE0sVD
YkuJTuRdVWGCATt9kmeRJWRVYxJjOSr7FLrXA2oClTA64fVeF/tMCXLOWplCfQ+k
dMJGeQ3BpDeakjnzSA2OIiugST3S1bYHAg35hJtjRNbf8lbJkCxoJjMn/ZU44BEW
9+GiAGjD7ZfQNuP9O9oH6zJIfeUJe6TYgqAUpkDsqO3hpn/PjHx0YoiCDfDHy/mu
ue985uWsymErSy0xJ6D3GT2EB+JO4wlsWNPevaiMS07mQwIPHosCUPNLWr9ZCs1i
/4/cZGEcWMKMGa4VD+S7mfU5nhju9HuzjGn6zDXyqUmj3Pwtw+X/edebTiImF08t
JrWXhAfbV4Ex+TVwirDU7gPKCBJW5REODpdfZKe8IZhg1HMO3U7t+wgKPpaY+Arc
IsgTi7W+q7KyqDhhwhYTGkZDoCeaiHyfk5GIcIwnxwss2c4e4RufC5pNZWHoUf8d
tTftRVMh7V0DM8wemYwdEUVvETt8woHO5M10ePcIBYuHARimsuH3H0rI6sSVDzXx
JkWMNWCaULEoSfcM1vp3HwYLH/1uE+Vyy0tS8H64L79roJpuFvzeQc1b/ZmoUh9X
yQpR1umO4U7JA6eygCXWIL4HzyJkUDnUWP1jP5eRElCFZ0OkkcB0/DY/exLHiQuW
TQwrp9T5edqj5HjVXrbbj9z0AOlLczGtYFVnAzy+NjFZg+C9Jr+Wm6hU1gV0yeRm
KAsIxFUonl38oQsAi9hovA1sJTJ+ivnSAhK5xIaIU4WJfiycNepTXgaz1KZ4LuZV
Xc9GU2+ILfXPx7c+/G1MUNvUtZtVWqvShCsTRYh66ivCcB70zFB3GsBugrR6UgNP
OB63s3E9R4hXOn1ANSi61aXxqhylcOiOdffjZsDW7aJm0pVsCV+ncX8E4UVMPEzh
Web1lVjhNrKMeuJlKiad1TuvjNj/JFTdwgMH3/reANExkA6IlaLtX/JzhzG6Sg4P
sDsF0SyId//YtWurbpB2pQxaYbl0ZLhEV24HNV7dBtGy+jlL3Itzuqv/AfT/USmn
4wvXY26EoyrfEe5SCwNJYXKvg4uGmcfwLHQaynH0X3Knrkr6+sux+oI7BHj7vVL0
WfasVKPFoQKIYIZjReUYKLHh2tmlzT/JS+UJUV/1GsMNvcY6VeItNSPRc6zxXjg3
XDqps88/ngJMvWMaMhI8pL6/ly7EeOm5jm8L8/yHtC6YiMVERFpa/jA4gpaHWSf9
B+pbqh3FKCUaBSw+okauwDrUvwmUM57fIZu6wKiQdreYSKk0gZtbTrlCnnKIgY6W
mTJbqHehJRQmbnkp/btoVUiL4xyk1m0KsSAQOazM9QZ0U5MZi9El/atKVySacQrp
mCfw0qR/JCep97ncmuzpNrqk/BsqWoZTCiaNTcyarTAs4rWkokZnv/k88gf8chTO
EQTjOzD4ojf1zgezNo95swRulTbo1E/U5z0zlDH+uOgKHQYVeMAAxRGqUnbpHtfP
QroQUov/KOqATRiVpQggHUs4j9NHMKrbUaHCPM9OYmN0yt3Bh/HrnthuGIbzppxK
eQ77GvyMWE9WoKyeDK7TBeWefP4qttQ1GEyUrI7K6vi/1Lh5AUHIF27AbdVi1dNR
BXYxdsw4tZgrqrBvrc5tgwZU8qW85mV80y9Sj5xKRBm7x3Wl5GhoO4nJRhsdtPBB
sN4O6pf9zh2u0aszr2Arxh59iSUV18UNpTd7SO3Pay8Og5Iv0zJ9Fq65d1JdbgIj
lJA+SfY6M6uoxnRDt8v41R2TWuSKx9ijuizL4O9rxmTa8Y2YAtnqQNp7JCZ7xSPa
Isps3m+BWok1tazth0YBYyq6wxcf699SkZLOB01IvxZsJDuLJNx69S228EOiM7OX
zg0HB/OYYVtwv8F6AqEeFvaFU1GApzJm0Hu4DvuqB9quwS35zqtXrzEwrVn82Mfa
EL61U/FSX19P3GaT2upXx0RMnImb7kUkOaXsVPbp6ijNoR4QfDViJmZ8YmTbMxu0
S70XVPtpR37Myv6Yn5aFXU4D26nK5AokDBjB1R8iFXmWs99Z2Y3aNUrNeAr37VXY
J2GY6TKEa7vmOmKiBieJpKOJoR9c2wyPak9c0hE22bGK2R3wLjn+fG7XS5tW1h7a
NbeWAAHWV/ajajE9L2eLDLkiNc2HHaR/1K4Fw0g9LOb2GHKqOzkXEVn1qa1zFYNo
BpzHmIwVfIvdVSBqAEIUz67FiMMbrMJtKngjjwKImx6rASpXhj/Drq+iHePqzc5P
rBzYKz7rfnCpCoDJWb1YkxTrgLFAGh3wmx0RImr4/ACI3y0IPdixGyW8IkjQNacH
zfaXQpwjGDwdCfpwW2Ogcs0w8pxmu2V6e1TyjwWa+/heezwbtY1mTld486VSaNCi
dPpG85TK4oiwyufQvvpP23Pt6vabJBJi42XOqY76JWbLPYbABSfFlexxBTt2yW3I
YsmS1QQrnxSCTpDSJrhgbqt7uemvMhlWW4iaEj+d4Cnn1pGa22INGG78PDKV1JIY
caDu9ClRQdCLsUW7S5kYYUs8iv+3uQ9Yj4mTxjKmQrTs8CtwvkO0W8QajyW8t0sD
gckqzma3Lok4AmQ6bCW1235StDVwGvAxAc2w/QDg/BrHtRvGewc7tIsHPk/zdHjI
6K/u3QPi/DreLeAeftyNmT6u/qLSCjznEpGaZGgr6X3YQqifwm/b8gLezMAJUtVR
UIiYFFiBdnW2Ggzpn4+hha8cTKX8nXG3aE9EaR8bcgqorziBqdEgl8Zx4XeYNoSV
RkANocCRgB8sNTvIib1HDAyzAa3ryrbV8vXjv1Ryn8A9Y+vnLno8yzlLinMuj9tB
1pvETl9LnuS6mhoYgSwBBvI7h2pOPcCFegO5ANO66LlwVES9v1wrRuNK1wKBuHDf
JsKQz5IKPpn8Gi1k/VcG4K8rn9mX22DY/SLxELVC+XkMPODsovBHwhrJdrwB6/J2
pbnQ++3gPyBoULgvOJ3v1ymK1eyU7eb9hWndoKfToPkYCBlg94nmTH7U064DymJo
Lhwas/VLl+WZFuucWL+s3K5jCdguQiWL9mxnO+nhqlei/iHlR5kcHjV2Y0HpYoin
C0vZJIyxbmO8pnkzKOd6NNQVIR+6rXRh9Ten6k51fd8UTB+bP0/5W1P5k7zSRiJd
XpXZg8oJIfyP9SWELHjJlq4JI+VfsA60l3Co4RTQEf/e6N7MAjorD/XC+6kbizPH
C70vYoWTua387uli80Toozf/FzWDYbfNoOm0xcZ+VBywOWR0QSg2J6P5Vavsa/RN
N51j4+dcpeU4+OuVuQgT8zLIoS1f1/ip2HBoCPu3KaWaorxELDL7EreRb4+tHXFJ
j/7x47Y3TLVzhDuNVebkacb1v3rk+DDZN8bKW95azqyn+E4cJKRnVDfDXU5ulWHA
C+tWGFSe20LWCoc/d9qz9QMsVrSX9SY6tbqhnQJSodWQfCoIW0l9LONoSGSK1rbc
hBH6GzhIX/Caa4CWy8oqhgiUVdJxPNRyHTQq0TFyu+MBQr9oTB3yct8MKNgcfeg2
AAmof4tE/Wou3lTQwGegUau7QLSja3tjiS+bNwi4k60vmFVSfWs+XF4iNg5DpxG8
+nBPP8/Hq94tm5mXpgUPC6i2wxLAUttDGykdDDzfTfpwBrjLeDLQfZPvOUV6Yq5C
UlvZ0eGF1F+0hNwOtFbc3W3BxVh1EJp1sypYvsD2CAxyHNBbbSaQolhz+M8/ffN0
lHtV4JhxcRk09a0bBzeGIa98vrPx54UXjYYDBuv9qOQ7voS/49kfmJn6BrUPT0F9
cm7EkuU7UWj/dO8BpU5rinuIMCO61ruq5c3cYU8yDkMYLNp++E+TI2xomdLn1IBD
e9pnlnkIoeNTHTxl+NM7aRi0p38wHcbSHysmEOeN71AMlb4B/eezfjloagPMSDGS
brSgiGPYAc9C6atw/vnt+CrfbyDXvN5DP9vqR8Bd9YiXcv8OsOL2oLv8WcrMR3h2
R1XB6LK2JYY+LqRXYuZIjhY15RwiIOhm7IfibWrS5SXEgBAXnPdaO9T6iGonBXQn
JoABgprm8kafX8qoiWzHFaI2Sx1aWJxMpCNQV5MG+nevecZ6AZjegXgV23o5SjLQ
bN+H5tr9wHI+5xrtUFyxKyW7GRpgePj3uaFfA4mepWMx1qQdf6ZXuIlKir7R+kqi
YuoS/lv3ZlM05krnv5/rx3hBFp/3w7UI+uiMbnLH6PNeV3fooAO1Hk0R5tBVBK4h
/eWO6ps0TDxAat37EP2sC7az/QzpWOky7bKojo4fs6KCFuD01dXoqV/+ug/D94Bi
FsjHj1y82NPIt5eVYt5FlkHG8RLP+E+VKuLfv3vYzBxqgaUQdT1lgO11nPp/CVlU
r6YNco+30LRZtha263iEYTfKs1tWvMxELjR078OhiDSSnOfrfbcMcsGWy/1EKgar
Bz9AtDJYspxHMW1oyhupSYjnCiKOCuYqjHr8qjyApGr2idnXSzLogfx0UAVyaGae
Wh/JCy2kiQkxJjsih+TapGg+m0yh2gR67Gmyjg/vnYqomjNclP0690JjtTQ/9Vq9
EStsvGU1KyAkXlux79quP61s1D11LXC+3sl9peEeeJ7oDw2Nh2oqtJQvKZmY0sFS
FcOtIG2a2ZdBhtvQWHIee7797/aXpxWYYoHCgYQmx9GZEMkL0o0Z9uj1gK8yThSa
a+Dv2WKkrkg6tLqSKA8b1v4x3qoRMBLOZBW0TguAhJ5u/zApxS1M30tGh+n+r2Wq
pIklF30iTw0ieoN6AM1OXi1TNwnd1hOopENXnmukV6O2isI4UifXOXo4HQoQADxm
KbOGgZkn5maVQjFsRo88W4Wnh1V/CpIRbZe7uD9AMyddV1PakyMJb6GkNrRp0Zex
/SuqqjKPWIHYoIXw641HBvX+/k/WUz/rx12gAgvIO2IvkoorsVUzOSwUCLNG07n8
x3lkufrKWA5NZd/kL0ZWnnjF4fTdJQrRhhyy9YBe1xeH97dM8Z/h/bmp8dZITVVM
r5+x2w5ZpEKewI1+fT/vNWMdF+yomuXzWa/F2u43zdEuXczvBRRGiL5ChG8HqAGS
9Wgv/O6ZFSRswe5jZWRG9PjLRfPPf4lsaziY/9o2Xg0iqYQSODgWimM5x9fC9KtC
9Ir3Auz5M1bIQx+ikahMsJ/Z8TNIg6PxPPPuji9Tx3Rl2CbxlK4IZ5SHMVK/U7jF
6S9UCkDN3yF8wO6ggbYRB6rFVCOPpoAKMVSzbk1+G8qSGQDkgjZ3303/Ej3cFRGi
RxyukgUNZehTcIl8Ov6StDR+41VoIk9weKp4wX+7pcwDiFi/5yPnAVfv6NXH4KCA
Gwx55Ko1nca2cB3Stnus/tJssKh4MXQqVZODS6wmwp/vi5ZSTWigwS214/PCSd44
R0NGPpNpzVWVMZTeey0yJXJ27Og1ugwN/mOhY1JZAcLyAe7X8odODyFyzA6W38v2
EFwy3ARAYZT/rL4rYgKbOOdn9mLDFtqyt4m24liUWOf1u1ZegO+v/Dco2GruP1Wd
6y6M2xCmLk2EiaOZ1u4kD7kalph/6ANuSLbq5Q+vpABbOIPgV9e3EHLzpsx9QbXS
TxWYIH+0QCnxm7ExtAhkNzHY7MTTMG6sOSa94CBobvbaPO3tAcb/dtMaGBBIK9/e
5Xcabo8dS0ZrxgOAh7DDrKmmbWhvhF8RRkRRboM5V2w6+SDJwhhsxZDlT8mHxhlT
kZ9BKxqD5f2G9q72sBqdSDOJ7g+WMs8t3OnJ8xA8PyIwHazOYn2HhHaQOVn08516
rNH5ZENB2uT2rXOGWvj3GZz2OBWospaeuYc98pREC9vynzBCe0ufh0ofizRuslui
1rmE7gweYp86j1GbYW9H/u7FM1HVGrItx2hD9TqnbO+3USQ7x0qt6LGfBNQpzsjg
6Oni9OGlipjfMBpuiCmFmrxLT/P8HJy8fBjQz0NHOMDr0ODh3K0HnYtZWmSiPkbx
4ILXicN7X41xuKJqWbpuxNp9rQICNrTt0ncD5CBt+gl14wF4+8/TySJlVuIsxybo
HF897Qh4t2g1FF+3LExPbubedTq5CoEHurLUXZfJvsulruqAZvcUsgqIKfdXTKLf
d1oM2nArjAHCL7xMlidq8tWQX/nslSqug7NwfFEqle29JZ/pY9DPpCrb48tobwIl
lK4H3EWd5musKcNpFpNpYV/z9kfp+brmTGAI4fsQetB5zZxdiF1VNcjpgfQCK2B3
Z5XsXmbnVWh1+kkmUoDhDXW64bic66lW+Xhxk3D0C4EKkD+RTRJz9zgJNRl/zY7K
1nl9w8t/ZSKxH6jIDYM3v+p83dkHznqezYGUkrbqL8BMQ3Rl5Rdx+csNVr+Aj5L+
WeP8cU3fOxulwFAPMSFaIffBkndXhWfva0Xh6vZACCDIJnyfZi/K+WO8uu6yEc5O
SxR8LZbjrHS4dFYegMtHJk9q+qJ2mBfAZej2Y7TVfbt49XhVxqPHhCbOQiqCib6m
pVd/roqJYu0ZcwVMf32V1FF692aolhyggoyK36c+yJ2CxRffh9kJPhAPY4EiaZXK
McjKbROAB3cETLsH4gnllIZ9gwoFfQNlWqzUQ4dzbOjWFcIjClf4IKYUCByMtsN7
NJeJzg+4pClMYMzqnQ4yBI01mygRlH2bATWvvWwd5QV+bEL/nv1GWGh3LzRF1T+J
9WXnQEM41umANAwT9CLYnVEQptvWQ2LeCIddhQluMGzJtyWg4nX62AgCucXnr5kY
mjWimuMiaFqIcIIh63H4OYiJrMVudxRZ4Zx64clQplkoDNsCKFEccZw6uKh+/Ufv
KWd/5u6SxzoV1CBiad22TpOkU1gt0QRHtRxIUlasYSWHre8evmkhcxM7zVHCIAMH
7e8inDiD2tUY06iWiTPHHlWzP7mBRIrr3QXJH4cn/FCzlHVLhdQ+l9micV4B/ccR
Uu59bPp7RQ4pOsGx5XgUGDDHTEDwyUd9msFl2gC8O1KKkEzts1BOdyvAfVHNAXls
JfGC0F0NgDNs8vkJzQHNbpvxdxeQKB6moud5kC6dfKC5bCUeHtsTZo4NtUzhUnBj
9zLQAFQIs6m0t+1GS0bjS+r6Ry5sIzmkNn0jpDzXC4vU+NIpAMTQJWNUYkwZ73S8
xoyo5VElNCDLkMuqpPOAcP+orCBDPGgy8GuY3asdmIXoL2HALwdJatphKX6KNNnT
YKYbTVgDGTeecARcV6bY7KOXoLySNF5EcOiG4IMyjxP2kDFN5S3dAr7QEhbe5IGV
zER0nFiQ2o1JRkJE2psppBfhn4JIyiNCo4sJ2Xuy+BbpV9asoI16EYxxWz+7NRJ4
GGWRtFReS0BKU+71koQzRP9oU15Tkp7HGGFL6iaxdwB1dWCZuT/KPcGCbrJUeWHm
r5Uvl5MyB3676FA5Nx8Qg7+UrXrMwRKS00rcx4x8vV8HiudXsyrYB+KSRXzFgEBy
JVltOr6BE2vNaKUBASVEAviRcBe1Sz6sXgRfZy1S6ZBv5kXEwSDNrKeIiPYjnuA+
jXRZISwFxfckv5pJ9o1lTqTYFx21cskJi+aOOwE/5tk8FrDsFg3DPM17nuJWrsIj
Gu4wXyTU16Ji6k3RjiHMTOfSD12ledAW9nxzS24LzBk8YjofRda9bCv8bQMLg/Jo
3mMew9fFb9rZWg961oHGh+zD+AZOvDDrPXDocgwEMKBz/mRLQQAd1gfdZ66mPRQC
fXrbFxDXqlTWC0r0jBRs9oRl+ab3etN6QxJ6QMpMxvd0VECrc05887u63wRDLhGp
BPbdiYaLa6BvsIrKjUZxOzXwX/oFdOm0GIzauQDVus3E8kXSuSnLCQzYFKX5s3fV
WeOZ7e0nCDVZuzICzeIP792HWsoIA/sMBwJz7WydLDwccCJh0vMOZpqrOAaL/v5I
P5d2sk30WY1fhjKheKGTmU/W6eQqaURhDoUrQotiH0NRn4McstrMGRppQoPXbc9u
YkASQYJFpUyAHIq065k5ou6XD6E2Z2HUQsjNeuZpO5O0mP+mdI0DK0C7uTm1CWzy
oYYjBLFgRRXtcExDCsPA3SiQ5NCyZeO0t1pp5VhnkDBzoK4SVOlI2Q4OGBNfLjkU
HkxRJVKYzyVMZZ2mxUv9j62hv9dEgpvYqB9rzVlzBMbX0guyXGkAriYhVxrK4XsY
ALuPUtwIGel24Ykyd+ZIkbi/GBeQd9I1WufBRejTrMhvA5A6eWD4NLoWFLhKVho/
PAWJ7rDvM1AYQgVUO2ilhGVfBisOb3dm2sTD+h2hUdAbqlisvbTMlxuSqNx2A1fV
BTmT3UKdDoUkOGrf9sUXDUzEzhu1aXADWBJsRb9yf9OMRvKU2WVFVG8cEgtrKC29
L8M4e0xk+VyvZWtOi44oPpKb9gayv5mEVJSGcCea2VYSmzflizZ/VXJMgWyTMF3D
Kx+YQby4NzaA+IefGEHrlgLC2CMzONgW7eng/ZlJtVehH1Ow1CwOIccUbtWFHZ/I
u00EpZ7N/3LvqmjIwKBGK6n4oJoC7DbfNBQVvcMtiy7qEKoTvlNBwhDu/g4O2xC2
QfpAtEEv+rwlWTS5RIgj787J9AD6NA2m/QB7AqWdekvlUSBSeyDHihpjuHB5O+5y
ImLKkPIqEhpJ8AfnAb2NUpzd2tp45bVp3UAeb+OrxfCYCAPBqHL7FYV4ZhY9c2Nd
boiEEpbk29gmYuFMkcK8aXtka5CojtzpVp5HqBorbO49A50RLQXBmy2jq+aBw4fj
yA50/pH5k0J+5vUvzKV3m+hgdwVMcANqn2FctwsqCCOgJ6fT3hWHjoSSdoPiL/UW
tlYn546F2I5l7ua9aScyeZ9Bw3X+A5nj2yQVkG4Sgng+auVSvcfIyRM0x8ko3W0q
BlscBtcfIOpQgspBJcmlBps69BeLv7ylbqSSJdbtUZ4g/mcB7nhPQ7S6sp/B+SPJ
YeQCveohbdWHABrAXM8SCWxEUjERjvrEWjN+BzmtmqsGMtqNb/wfJfmB/pb7pzUi
zIHjG0pEbBkC6pArIuvltNwXOcBkMPG7JtQ6tOQ30uzXUiM+tZjq6ZXz+QCyXsBo
V86nToFx0m2qwEckJeS6XS7PZlLKaG4vOSqKHHwr00+uJM7r+kiqSCXnA7Gb8SIY
f1cZ8RS4lyvEceK0hOSsCh1GdUBNUlnVSdAD/GByEDN/nZUabe6bwfy/ikL1ZX9/
EVNBvj/tlr/ZekamLSrIPV/iKmV6FasX/0speWzM66MAV/BmWykONdRZrSED48S/
+KAcxmuvJL1dHbqrRuA8d0VaI1hSbN0GWxBaTqQB+zJ7fr7kl0733Q08YzNpmzTS
rWv0kI0vUBAYslK9VPheKdJsYHx9veYRzRCrKWCaWh6tsBqn918e7GEPArGF81Kd
0Oh4Ugcau7MiR9I7Nl2TTthtUyM6UuiIdCmyTbFegjJPtXDQTqJVaTMdVrNz9e1t
aAeQ1udugI7fzMBZfId8vw8eUqqrgAxcKRf1HLas54zxhFVeFPkwUlSnKj+LwYuM
D8asS4mntlGj3C/gBNfWNiSHMQ/XSxveoCi8WEMC0ydr1NUFSc9ITeFk/UJYh/h9
8nJRekwYctieHmDkiEAF7v3EGfJLJlFEg1lrpSbQre4v2jDUQjxtXsSlPzsQFf7F
811io9FQxl9Q5eLMKEzUh5Qv6iyguCOjPe8Ei5XnqpJna3pyXXFVt2NVrH1B68YW
v4dNzB8qqRvsxNr5jB6zmHvoQeX5q50hVM8WCu04a2vLXmgTF6/x70IqfNMaR7u5
gPN5nUGVI71p0URGebQQg1p9dRlHBWQdZ7xd+CJMq+qgPCX5T1XExVF3ITGew9Me
TERNqU2ICIMLVFAN1uIxDo7MUFHmu5BhbfQ//DdYVjn4bU/dtz9u1J961cy2EbpO
iI+Ku+pb/0DAXRa52uUBLxcqfLi3yVVBXThyxmwFNmyBTWgRn0mS9DWSlPPDXqwE
jIhjIhXksRSx1RQDVo/mebUFfB0D1bKCbNvhRTklCU1hfbyVC8j+wK72VN3g4PKb
+5vtifzOQDPxlC+JP/OeumKyWrQ8kV36bDoCXtvwKc58Jj21YzbSxqE5S2O+6SzV
86vCglFjRVR0vuf8v7DGDzTBkZYVYu/jIHhK0hLFQYEt9p9zE+6PWvbo9wouV4M3
JKidn3iuqo+0gBCSa/1XuOYWuX2XG6h2bwtc2e/e0xXjbxkp+6w2DAAnIEuu8zCi
Chr+bu2CQBzgMa1nB0BNWY4u4DYqBrC0/bTsaI13F/reeS/3GSjf/rEApfmPdCFM
/NINcme2QlzE/fEO2ynBAhXnIyjeu5th/Tg3NduajzBN8jBBfA7Lf5rscgSKehv2
reAvhhDAHKTbr6Un4oiKwRAqpvPXu2uaRydbB183eSf+3JxFMKT/WFI6XHCtwg4X
nQ0cx46PwO7togTLtYQGhoGVZSCxZHE3DjNDgPoEUTqsqRuY7gKj1MFX9Of5TXEt
6Io/wQ112j7ZCJGDkmqbskVZatx2w14ZTriIrI7UYp2jP0DAGeSq/gbIYNza/Ud0
TI1IjTdR9BrL1m++B4irMt+E+UvhS7KwslZrMlhQeqsEdvbZ8QVJDMFJ64iXBwyx
aoX6N8Cv+jKk4XINzv0lV6oxs5pQn3atoAjvDuYAtCa1N/HscIqwEkOS2/ZD/Fcm
DWSEA1O60UQK9wOYkZIN9T74Chhf7nZRawADNqAsrgHdrXeZ2QmxkBwkuGKfs91Z
piW/ISc5X3ErW8VF804wbQLiSuSm7VQqfmEKvg9meDAlR/xGrA1nX+Ajb0RW94EZ
995puDJ5aGyO1Nsvds8OAW/pv3sEI8/Bs6whnEbG+L3sy8hXqMmoqTHjwR3PHlAL
XrUDVI4+wNiMqvipfS9TrDCaWxoQV1Zo1HsQjTJnuS5/szqBlpBQ52HaOrkKy5Fu
MGdPvzMkipms1NHnmgWju0qSQYYJ7ctnILA/CSC5g4B/wu6QXV4i2jcF/PwnsXUl
x426JLR20xk2XVxs+N5Da4/I/kazsjDbDb+umOE1lurcgb+E9KNO5iP6OFZ56+kR
a1CQ3C7Tw8T7LvDfxOAeC3c8QBacXdaEAb7iwJahbK7nqjfH+1+6MJzPRstIcltW
C6ZdxG9xLVmTnXyPy9aqrBixR2jQjHst5dasp1B1elwd7UtlkKOYQiqj0KwZeN7K
4bAI7oDqBzpMgstZTN3btXe+s7VsHSPU0DXPsDjrBxCDV11ffxLUBt2EqT1kvZXN
jKgbJ1USpfSuQmlVnzqSxmdqwDEVP0G+zzaCDeFXEFKJ/05HORrilvCrM3ZUz184
QtysDRFsHXo4CYpqZIy3G6qDGimXQykp5Nre1WZts8BClon2a7bNF8LJIvZZuBX1
fuiUNDc7wZmsAFWE1VowitWDaesxbFsrPcfpTcfbS+Ctm5bbKPXdXPMp50qQSDeS
QsmgW5sNJf9Zf8u1tRlf/V6C7eBElUIp4K0XLatxJe0IVcQJ9e3GGwezige7rCDu
EFrOt0+fS2b+yGUwMifZrl1LOJ6QW5Vpik9iXj43zhbaasH4TuVYjf4Otc+qWpYq
AGirm44D/dY5QhSpRfggq+zTPTCp9Vx+R317TtO23p9MyGPB7tAE93iEV8GOgqed
nwg0WKcBJ/CEwmnKE1CN9Wgj7/U/TUcpCbSsYgcj19waTm3MC0KnvYZmLVsuWZIh
jdycGQgLVKwXmWdYVDUU6yqMfVmuJEQusRYJys/RWBSeuovUURj+DEIS+ieASdAF
S/1VOqqkMMF+a1e+2rhHGXQHf8gSiKx7kVfw7cKhxC0DOmzX99Bdo1zuIeybFb80
h1DJHM3M6WJpw4bflsjhdLS/myZrcCOaBinoiUzAyBWVkgYFkDL0TKcVFGUVrgVQ
fFcp1MX9I5FOLJldIab/XYaKdj44rFsABosAshMxR3jvS6A/A/0hhCvGR0E/2XcD
G96Nu06N+dgnx4VcZ8UOYo1aJZd2lpJQzZOVBaH0ns05Weky+AKnV1JpbxSdR1T+
PEVBwH4/tR9JNR0hlEfndbnHuRdKNzkyHARhravx5MnwfBli2FvDFg3Yp94xqTQH
9kz9Roa3SDDgK5H1sk0NHFop/kbXJMDcUHDOscS52PQhN5R799GDyS2W+YXKoUZS
T6Cr2N7Y/Xj03rKio6+rsY9M52EnMe3qzCJaaS+PgYaAPjrbdnaMBK/GR3Y0DW5X
QqFDB7XcyzCgs/Cgjatjj8uT/cikyfWpZePKgus0GRLnlZgcyXSTCzL5/bRpy2sY
VLRE0yd2sPi48fw9x+wv9z3CvxbFNtu5wuMCMAI8vuN9m6jPy30dZdZkywq2mI/6
pSGd66DF8Zfw1DJoCVZsqbC9v/RVXnCCVXBhpO1IF82/9hhAEkOTUcvumFeC4hRw
NlRVL9oa9i6BrWjw7q1KJc9s2OTV8Usx6jroRyI/IZkUUbIOy2TOym8h8USXdErZ
Nde84DnhAOHcdQlvjjeVWFu0cDVB+1WelUml6CP0b97RwkuQcj9msMk+JdiK0NW0
E0PqH1cboaUFbf3JkZ7+6sJKAaOnGsQGFIzfoZoJaDhDHTMrhxTK23MPgdJHJM9m
JdbULw7jwjvknYNw/giF6jO9s3id/et9xKLl3oNrS4HdVU+Wgi+K0dvTrAV6iOSV
EjAn5qmPTrG/pxhrlyWAeBfcjjssuHbeRmKIyDaGsey4k/lqhq0q+e3oluqgX/16
RKzeVvjMMsnGMFMPc1/Sh8Rwz7Y8v8nzItkFqCGqr0buetLUkeRTMX0OpVkhBHWm
seHgQjym1fNelRDyfVeCT7gRpBONkKMCLCQyc4qXJLDkJrY8/R2o1N1hsapDNTPu
pEABhDqt4b7Jy5ymW2pCarKr+wndvsL5qv7sksC8rGLKX5kBU++7xk/41EfgVFGC
q4pZ9Brh4WCJrNG99z2fPzRxjiqVXn1uvou9RYPke4KSZyf75aGe3lxpcL8fB7P+
4Lvlrpr0hssNUh0V6gzF/Fle1MQ2bys/ASZ30x9ITDQJllny20jm0HcXzwUy5mp8
ABBm/PhO2vDtfY4v9+niJ3hJiM8Z/ls77oYnDYsc8kIgr4m77XUPoxazAO6gdUkZ
iQ+YrmSpMnUMxqhjBMdrc+xj4eVU1HwctvgjaJ2EMRR1p+hT/uL2rBuncVX1s4wV
I862r5ugOGtMTeBkij28h2vRar+lSc/mx6HfiRaRU7wt30lGVOo14MMEPARQKVRy
UeJUdHvIzJxqK+vXtbWJ7o4K3e/9c/7INoYgCdzUkHTWBU5E+L7jqqTvakOcgwHV
87nkst8TXY3AZ8KhJDlE9d2534H6aZmlMx060aSAOxqnPGWCTAgQ/AJvuOqFuLbK
1wi1KDdmKb3smiCgn1OpuwYypA2SukyGRk5VdSOGfhuzYZ/drJKaqTkgEJOCoaI0
nVGPi8ehiwH/uMVtF9PNg7m7gqa3BwKhgE1a9BuSAian5PLotFqR9gjsUakVUQNB
2HRe25UREUeL6cE/uH4H0bGLFw72pe02IMNGjAz5hqUU0QYrC2K/LFeQjUXWwqsq
TA1XM7cUQ+UOGHtaIGBqV4fJOZC04tI4wOLP2RdCJnJr3ycIEuVUBzngd7cPaxbW
otJRSeL2BlKCCOZGfB590EUbQxrWSPc4WxSfhQZNKokx6zWZEmicqjSjUnZwOeY9
jqnz0SiD4Iq8vL2DUMlqGNu/4v/5nh1oVqXWX+myxBUXJVOoE368OZu6hcxOHXTN
EtPiaXC+axez0qGpgP7CvI6yQuvp1cu01nPV/2BfTQO4Hgz9fA4B+N5fdA6a+8l5
gHUXxXzwTf1JCVdcV0rE2RPWSjxYkTHJ/ADqfs5VE+ioIFPemXs54Eu8ViJT/ruL
4bd3XGUwfZXeQ2WEGej+whqwjD9+oJYjXHLIn5bu18iVo8rM+9TFoXorQHLXQqjC
njSFGe0kYjmB3LqnuR5qZz68WaDlByOYdbrfBIfl4kjyv6O2OBO5+oPvak4S31KI
YDohAixJrvRADT6bUj2iH3lb6I/WZutH6kkfPau4J+b/TGK+VVkoe51qKfzadQxg
E7kV2gs1hRcNvVuLZcOmuqxczJjv7KASs2GZn6WVSJpys/09X6yEE6SPUIZW5k15
VIcRghOJgHtzopMAoUT0rVVauw/uM1fnyUK7xwCYKy+aERAOmnRdU+POz+JxRerc
nf/qtdGO7g4ZyhO10087VefZZ4ZM/dZnlBKhB26cIeo34ihhn35RQGe9myRk0Hi+
6cJhKcaSQNpFR/1NKEf10OZntsk+qx6QS0pcxKm9D2SDhexOSvxsyphyeThZ5Ywc
IiKxkYohXuR6CiN9u5ro1ChlsSd3/kYvpQFPjYEz8oydxZbtbewhQET68G/oJdor
qasSRTFUV7N7t4rjSE1s6tmmsfuO0l2vq95WBHtEEF7UbDa3OYHxFpGPn7978LhM
uExyKM6jk+EV/yHhNCIpsPFXaIRw2uoBF5TA0Wqtmo1E0cbh3NXrS14GviwtEdwI
btf91+spWdG86LGaQAlqn/sdZzxVZMsXJ6+gNvN/5gOdW0VOPMTD28iQs/ZjBfHI
r5Jv7npwYt88ewR8LetyuF+nou6SGOtjRb3HDNXfREBOmL10phMrHvQQQqbWnWcq
sR9vHOD6JXbSb2XfpYw5Hh+ndNdW4IYhh74HQBznaeZhvJJ9qgxdK4x2BtnzPeRu
5MPfXYawd70KNHwzzmsBKvTEzD7b5c9mNR5WfXTTfRktMDlBWwfUf/b9f2yOIPKa
NF3ung2d5Yvtmo1/2iWLATVYIQgzIobrjvaVA1oAKbhlSQ5fO8o5Xgy672lSu0ML
PzBmRw5djJTMi5eIrJKiCTDsjm31pP8n+6SkFBbGRUNivMUQg8WhXdoqKO1Tgaw/
MNvsWGnbLo3KwnTuqNa4Ue4UfI2+LYvK5w19iUg5uv7p/ixHWETQQ817pp++eo3L
tre2OBQ/Y+7YsLuJNAMxWklI75lZB2pvwsoySxqwwurAOK1F9iO7BOb5MM/euTEw
F5+mRyGoBDCNtq5VkbnRoesKlIXBRtUBN6jDcZYqLkdsNaT1wgU4WMKSs+snKuCA
irfqCvaPwmzEG2Xz8SceExFYmyPbboS/YPq17tj2GKZMtKQxxc2FlhLpPt7ccu19
AWIAdNTJGb+EmWOheHaCVYOV0ByasYnG4kMSELhZJyc42Zw7Pr+trChgxGPBZ7q6
CQkf8+XOmdeLOLum/upimfg9JTtjDO9lm6DRhHrB/l+0JlnMPnlqUJox7YRpGvUj
t2Pm2QO6ys3GzUrHowYYXfW2LKT7qnJ292lgHfWaIvRWgDV/dfuX77sfIjjSdwEt
YHkrymCT232+wjDYNdfPfFRQv86Gj2YAK/JYVAdH5kHdxfNoNS6B6uEH3mhEOYPg
QVXjEFIux5CYKPt2khomwRYHkV/LSzsUY3rV56WJMvwZ14BQdwb8qpjYlFCohVRb
0qPFFHJPtUmQxR8mVbBSm5EOK4LkfNxNGNiAkb8+ZjgPjVIInm+FYHlhpnAqhuWB
gj3fAB/BnMgQO783P6EwqF1y50N8G0yS6mOfbhmV6xDjT3un1c3VQyvOE3ZUmUGO
ywVb9pY5//gFHNQKl0EJCUw2PFD/Zw4/Qzt9ysM0D/j5vjEC/vrfN80iXpdUlpzr
6c6eir0yvlbgBO3k0k5NQ8fxhCLgHisr4OiAoRKCfWau7DyOR855ETB8Q66MoY9P
v9FjEpyrthZm0H6V4wYvqimDeoSDbTXcJID6ngNrRwnHM0KUZ/wpbrV475c1QTUs
szBitqxCPADrb1vs+7nXgnZXGJJOBn2LKB3GPNHTrBEX0lKuB1bOPsyvznsdIn9H
RrwJfBlDPit2Re8jS9t6WyWsQ4Y//DuMbvBDXj5RNfrHcjhOq9VZQIJbNmzsbGBJ
CX169t+2URUvHOAQMkpdFCEqc0FHYCoMWGbt9AFhOWnJrazBkudk2Ql8ZYO72ns2
lwiq8RKKNJeJgZQmldUmg5BuY+WI15X6xyWOxSW093LfKAbKzw/x4o7Jqvh72MeM
hY7edlZwk+jGbIJRSGraSL8r9Z+qlq2VpLkvyvGj4lkyj7YLY4ZGnYtQY9cUEmbc
eg1qlzyPfJtO0HkqgLGHvAkw7rk0DuTCiqVlQPJhApsXKqzLxh2ZrWF6ArqsvnGG
lRvOWkhNhaAylVRi7/6YuzLK9AGHTghQ0+VmXqjZUrsnoRqLyaAQkIYpqNHkpfxC
V4RiqTlQs25zR+Uy4kGG5fWh9ubsyS38qtr/kS/HZoyrKWoRhm9vMZtHgV+pV1vv
3zab4mZO1EleukM6mxa2ErfA8WfjokiVyB+o2BnMVFFFRSrlIc+AQn7TvBx9yXag
I9RBaRIY086vN/cRYKWRTeQ6FDzTEUdLMXDd7AwXH4yaTfebpBp/RpFk6JqWn8fd
LeQm3UhQ3IfFk0WQtD23EcQ8w26UQU7onB6gBNANByS00t/wrCpDXSRXu6rO9kmD
dGgmq1mVKvrwq5XEiRcTS9ueq4t4pQWRUgu85penztQUtC6xPLph1l6nXuwfetGC
G7ZRtymi0bKljiNBs+JuKU27CZhjg8GqzQRD6NJx2cUmQW97COkRocepBqJQCGNH
Qy1zB98y6rKJVqmZzL9Qia42Z5SvRhTCSQMlsAISBj4UAzGpDPx4b3nZAmjtjyI2
z8OoiBpRJR+tddiceD40Fc8LS9BbPS8GYkhVcDCtp4dHoJOIG39LNo7FNf9V/Tb+
FEq2LkJTtT32v7HLvjA+vjkUSkAR7epONBuGBL8EUVkGJRmWIGyNcJtZpHrjWM/Y
cjqg6ZOGOEIM22vDADq4Smhmiz4CxxJMUVQ+cqu4cv/WBNQRqZqCfTmVvvpyFTPy
fZnD4wPzam5B+VQDWIfhXEcTrfp2C8kbVnY7Ngp6T80Rp5FCXB2PJPYDgwwh+sux
VhCT2mL/aDDUiABG9Gmyd8pdFMXRunHQxaq6UMxd0ORwHSRN132a8CVC5vm5nqap
/FdXDQStdojkSIOpCS+XsdG7J2KM1V1tiCO3Jk7uTcPYWrv61T9McK08p45jHemv
xM0wwHBBi+ZpMfi65NqTFXQCTsUT/JVM0COXvT2ow28wrzVKe6Gy7ldaZSzq4KvN
ZUl/JKPzr7z4ewzrsox07Jr9cm6FN4zMcRWeDE/Jnf3Fala5BViuwqOmosKC4QMZ
MVNMTkwEkX6hF4JACx76XRvC/XXnTFGRL2ADFDXrLTZpdt7SDeQakdqFqh2LhmWj
L20anB0NoCmN3valm0nSl6CM7a+At+F/Aq+QpzSSQZ72JHETLWO4pTeM+fneiRU9
P/zdajCiI3K+xdm2wrtntyKhAHxzUN0E5gn4wIqSoxpDxLqSxJn6GSn0epHlYdiZ
fc5ODAJWOF0zfSecUzA8zuU6u9cpdoR30ad/3Sj7Mlshg7L9xCSuME1T0jxg+2/F
Z7id+Okbtu5fhEesQQMjeXqCH8kvgiweah7tJrlCL/ei2jErcqsAjOm58G+KNwHP
jfbmB/1LVFilUfLSOKkX7kXB17CMj2fZsvdnzPw1dCjFQQ7Y7O4dpOZPrdoevN4J
8hadpxu1zlp3C9ZPua9py4yp/00SDSA2b86lQjhjEA5nYlshtMj9V7YO5baTo7OT
BiUNIOMiOc9+jMzqOZsUtyYEWQGnhsz128SXT0CYXLvdN0l3DB5CiR/f9AH16uCk
9Oq0Kx01n7SZ7+ai0EwnyjdUrkb4h7Tu4tu5E75OP46gLoouJdYlWZi8tOjr7/rr
ddTbrjZ/NiuchXVE5pedZDFrzY3OVasrx4MFYMGhEC0pIks3yj/SilJRuPaNPjH8
RUmces1ZJjLt10ovPxWikO/FCUP80PKbdv0Qwmug5OUHucSF97tE88Jc9MygNfjq
f0aM1JJe4xQCb1EstJRrFNe/ZPyWBP9/fxnmxSUPO1m/pmcfa+4/dKHuGrOY+KWO
4MmwsDeCPw9Ml1GuXSkzp/8FxCQrdxRuxzbAzA3oSdYz5SP6OJPEiRErtmPvNfpa
lKjReLn39Ls0bOQUqqbilem8nwCzhumE5aYm4D7YP7H/US9QNCP921MbvgxnKJ7j
Zi2FExCcTamaaqeoI4tYVBNiVp5O5YDIjqIAqT1VzPTTYKPgQGN5+0MRTnEgSZqz
aP2KMn4PcwhxPDM5sYFlh1998rg1sQqc8YSIICMj3fPC1YyavqeC5eQLVAcFp5is
d6X9pTzziTKiZeGH2aSHlvfGwGb+E5cv+zfDc2wkKent9OD4l7FhwjgKuy4qTmyG
M+2A8GT56pUnQC0vhs/QzwLsjCX3PlsOTfVf9ccaGsz8RmSv8nRNFhyJK2C4JpAN
M/EJ5WXI1RfHtiwIgWAABZJNUurDxZ+TkBDVKEnb+JglLkIpfkMS7OjkF619+Q66
I7xr8Uqz5Y+vBpuscZgg+FUs087HSWYbUPsmE7sUMNgmugJu2kkGmb4SIGJm06Sa
KMRF2dCLNIH7NnKNwfJ5+QLs9Ie6Nd6UI+iuYhjI+yltL+Qz2xQeJe0V/X4QYK3F
2+GkFd38eTYSot5dgJ2HyTC+iYGARSvuKLe3FnEL12zjIdFat4mxt2nfDuNfLUDs
FY6LtAKkFcUzjKyAbEOGG8AycPGx8rWBFz/Liw2Xme+S8JfhSbjpazVkLLSO+Kw+
dNqs2KkS9CvEDWY3DfNxcsErTep/bB7SR4TLEUjVaja5syNSg2XMDwOxotQy5n5U
W0DM6wuhGDPpcscuz8fyIswOVDtqbWas5yGPWMpUumpHGXW1sw0/2GqhK6jKAZfY
`protect end_protected