`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinrC15oaCUZRxOKQkociLGV
YDFYhotxbwA/khnbfb8aQMy0Nic0oPYTT1PeBRgvHfEZpas4wo+ZaYe0bKTdCuJb
zSUrP6/QnbQlO3RodCtL6jX9ueYmxfePX5f37FaIS2MAh1LDH3DFetgkZtGlOQyc
Y/S8xuWre/KtkfqgT4nI0QfmviekxzBGxliXTiN2Nr4BmUyvl1yKWN4o/8K3tAcn
jDSV+cMaf8FTDZslqwb+782mco8RcctvGwS0wo20IFbWaWDfzupP1YZBZtDDxxZf
RzyUI0+atvWrzVKB+OrNt3tTbqNM5udpGlGfJV9VHI127Lw2YUmVQI5cBMo8zUos
qnPl6GDkVmXr+6UfuWlaXgynk+++3bl6nptx9HTLAEZXraBeoQ3cwtLvoBRKypf3
Jo7pwHusm9SLgJN1AIxd2I57hxJ4X2q+VETQ/8CoKKL+eS8j9iccs9NU3qKcqFsG
qr2p8ChKQKwqasMWlAJggfmjxL2fH32Cz11Oia0mQkpZ3sOffcjik+mydaz3+ZF6
c/jCKS2409APpoiBsWHJHbAtY4eWnD6QQbnRbAScR3zqCs2w2695PV6IeL6BzDu4
AN5fsQW9ZcUq7U8sqcEF5xcSPHVBWOZImJ7TQVJqzlUyJmeJbBSchdZtvvJS5FLC
oOhPgxHSxtiTEG4aPaTlRBB89c9ro1WRrrwi9VFmd4Cm6ti/xA1+0YKrwjict6B1
VztSrqvSWxumRiCDzxwacKx7z3rT4pqUYcIU3LqhPfg7jx7/QVcloS7MvNHyPfMK
OM5k2pqUh1XAYwW9IXqfX0hgKivTn8eo3slVH47xrY5s4fe0IFFlu+38enQ9zIeT
smzC6sGfRUF015/QD5zkKEvJ3qHKiO0kfe+dFzcGm4khr128HQfKxhW1132WG9w3
F/hs5DbepErGwwgHjwWipZ5lXqLz1yY4k7jh4zmHlyKo33UlOH2I3vUzC1Ono6Lg
84FruCenu/i25oTNRVeQ60tGw5VINtgAAvDgGroyhcxA02XpkmjB2sjZ0TvvNSJW
ogA81aXawJ38EPNi09bICretLrzYoEdcJa/ItQCF+m3HJO/konFA5Dqw1MYujrRm
G84/yRwMzM/VbYqHreALsgz8qpemUoGqamqRdc49voTch7Byq3Hbpr5BQkJRtR73
v1pX3XLrHdka3CzZg3o9CBT7Vmr1zw6ekixPl8vib0HCwUKphZ5mBGAC6pOj2GeK
fkY7hnzZlXeqvvbQFzkDepv5SejTzB9W5mmm4ZsLHKsNyDmudK/9nBmQjGuhB+3I
VsdF4r8TIW2PsvFeOG8SBWFa/nB0EQ0EGtOogxm3rQSEkTyfA98U4Se59BPBCs2K
FFb/p+Y+oew4h2yqyMQBs6i7B8V87qLxv+64y1a2MEiuAoEW9rLobkq2dotoQ9X9
SkitROQu4gJnE5MLvhyUZZVpEuyIFbhtS0cnHs8XWWSnitEQvxKf9aULzZblH3uq
25qcwtZ88xLafCC5RdfFT3FmgwTIPjN3SkqffVesUWvsAlz7Thb9QZj3nPXChDkK
nY28aL6oipubKFE42yWS5p9gJYmNX2V7GGMZ0F3Ujs1+7OCb4TySj2izq0synw7F
JvOJ8RByINANb7WotpCB0QLnA2TafqBkj5dUwuHU5HuURKbruK2Ck79wTdsY5Te6
Iy+SAWMGVNjN7SZ+DeeqM2lPL6NYmK4L04zHsChqGGiVOao/Vk0zHQ3gXRAoT5kW
cwXJdZhpAFGaGMLJUshJO5/5eqxlHlTmW7R34dVYa/tSejsBJgNwYAHgzoKRq5eh
fyGxpm9Lkyxv9OEkInCNh8tFWBiKQ48OFlGPjkQv5sD3GafK7zXAXizRLNtWvRHv
wQSFJA/2hfFKTm/QW4IGNsan8M1BOuuUfAQQoATrsuYRVACegIBhRT7aAdTstGJO
zWT6GW44AR3OXjtwABVmpPwzkpfLj+HonrfsPh4CdP39krQn8Y5IwI2XuAY8rh7c
Q0E3LnYFO//Q6FhUBlQMV5owBCV/8YmDrAnD9AsX7v2L4mOdeLv8u8nBYIVg6H0U
bcParwxyfYtfK3dcQnd1glj61xERDmMwzEhHzi0nN4wn/x8T92AfmMHBU2yGrh19
7GMI6u1gDIuPKLDe+HUck5TfdYzj76Wm5QqaX9+c9kJ5ruc/kFu1/JfxZXcYYvwr
AvYoUW6ZuesISMaf9MJD13TpJRNhIoBGLG9rVGU/Yx1OuXj3/zeFBNvhM7b3WNPy
icDlIsOuOl6kmRiaaRkpY7vW1MgvhisyD4i21HdiOmsjfou12rwXxgqjTxoK22Yn
J0h1lLf1ABQKp1reyuI85TleCj5R2DdioeeDPr6XblDO05YN55tEEban+CeAoIPQ
VMipm5V2LFHKAWOoSaf9OlEuwxmg6+j3XOU458M2EufAqay7oOelz+he3Id8I45O
PICxH2QoDT4xyVimNfpoAN4AscBNR14Agq0L2IMKfOJpu1tUztNHLpwwW0dG/9YY
sZlUFsz2r81Nv7cgdp95R1m/6qbosEWSiZt6bVjRCdbPr1jo5Vk/KTVdRhXmw+Dr
k+A07pLaRckHZ7nS17w4/CQNdCCE8HQkR10E7NZ7W2akNOmvPtrbWwRy/7oIGL13
Ck4qWeqZq5VVY2b85cc0LD2UJ/yyiaPBCpqvMZ0UvgS1jtuhMryfMV94mja19Yck
PzFyiUCNIlmiLHZZt5vFE3oczOYisun1VuYDnbyH0hDQOZQvm7oOZ32QS5cx8aoB
IKcZhHwwDbrLNrv5+7u6H2vXysR0thjrcWGb9zPQEcFbe26Lj6HDVMGcHvu6TLfK
YiwyJtQlGN8pEtloLtN7a8tfPxybL9HBfCAJdD1/IawW2DjmvhRIUufL/Mg0K4GA
sqNLs1jNOnUBjiDR2eHNgDWE4JXdhArLn1YACSRZWku9KN1NG16dyHsFu2WcHTum
Y3yAB6pBeJItTzQKhdmz8a8rLfKplaMk+jpQMAu3jKG9Jk4QGw5xk4AtMRDV1pXu
SDmrfmicqzSOxkb/pBlo6kj4riN09fDZmBtlILbCAYF0J5rOoXUgvX5Qp/780nk2
Dc41SnE9bESM9HPlGmyqM5yYYpi85d19dUOku4oke4307Z6QjXHqxqcVPtezb2NU
u0sWyXa7KbHhawqOgvYysJSXTGLRHacVFquMlfpa4NEaVWxux8i/lzQl5uPZizRz
lwvGZ5mqwZpQGN0GriSkqRsJmaxgyfYp5EjW7RFoHfxOI/yYjb1TKEG0p8QR5G76
nM2fk8QdY/4JZ5PKsVLqd+q/Kl/dc6uF+B00JB6mG878VonLyu/Iop5uluUa/SfH
Tw/WFvi4bvPzt6/sfPsSVF86mgdf4+qfq03WOeiIVcXBF+iC0UKkefFwYKmDq1IZ
FL8IGSpd8SXlzk7iapy9QUoErNVFnU8KzYHNOu7aRAU7NMGwJeu1ROEXFy7u4zC1
gEWxyTa9e6ZhNxXeLSwDzf0LgLYSDdk8dcbyJ/2u8ck12wqo2STZQGVBonnsb6B4
n5RKeZbB2Augg9eOd7EQlPk04zgrEJ3HHxoaYQZtaN4AIWPrTl7Wk1b/AKdxqLDG
CGVuz34BPjn3CgCS7JDQEWhi1N/mi2cgYthOKC1fDr+R3OWp2PHOjg5RqpSbxfRb
tCijInaNUjgTLEHvpu9jB3sZptmVEfyl95iJZOGikXNa1UAl4zvIs2+jQqnW4QLd
Bkn8KdTtdyj+E2LPMFEbZ+awVsktEmURCN+/WxkvSDbbHOure5XyLz1vuCbb3A9U
FMEXuDGcniBZfzpXzdAZ79Z3si0I54ecQ9dpYvO4OHJrQ9gdXNVxTlD6+L3/VHAl
GibZ0RsdTcmQSgMe/4e7YiK7Ioe6eSSsuei1jzp0LOwKk2DMoo1pWYz8hpt4ePIN
6DVnC+QS/sLJl/Kwj9LLFLdgVmva+zOs3swhkm3uxx8hJ7IB4nOw1eF2Nj9sKOiv
YXU1wJ1LwGq1zeTA5unK2Q0Gwbpz/+0U6K8Db2eXjOcEZDYuh0nPPv3MfdpJrUXb
IRSHgCL/IL2E9BmR9Jh0byDyvqy3lmmnG+RLfa4UaXJFaVnqRzu3yAP/cBBFUbIO
YmncaymgHXpJ0MpPiN5YNiYeUWNfVEvjrE3DpfkB7xQQkqX/XNGlRNZMEFNjjQbS
x7+uj/s6cjfP7niUwKlUvdGxLfrUn9Xc/B0QINZ5CP4PMl39ubOgTyqnEERP5NvL
oqmFxt1YMRwpcWbGCoBh+I1EkAL4XRcQwetP/dPgZHLQzwexJrkNPvC/msmB+VeG
bCScO2SExz0n8qhLQoOWjD7/BxqYtRrIm5DjdpgEjs+Fu01mQht4/2YEuhoL89cQ
i9OaJtcf9DASJ63mqFS51XPgxS/O8zqrOvxQMsuXFcHJr88YvXJXMwOWO8EHOiX0
XH9gyyoc/AZ8svn/Gsaq0KZ6lztrFSDZhke0soAdmse+ZvYBqhJc8K6nC80Fi+HY
iwEvd1tZCFuWx4yIOxUZ+OHV59Biuze1VSQIfnpJjaue8p9YEm0uibZda6Pt/SlX
sw1UwIAx73cf9zqyaqA/Qn+/PJuLJAIMsagVHVvxadZxfEGK8CXxNBbfKP9BqK2o
iP+iBVbA8FCkkdIsIEJUWwOCy63Ap9oIHQJfdYWBuTSnbvvylaTPp5xNWTroex+F
hJxIiblSXPf2GhmWr9KogTJGPvjkFWXmpxua7av7Ah+ItjrYx1KNERHZoyCTFKkH
dJ8vqsUwh7CkjGy2Rau1WdstSKW9gCv/odktqv2WkgH1Arr2GHoArSXxzCPJ60wN
FhT/XzQZNS6nkp+3guE85RnTZYok+KiARGLh2KbmrXpG/0xKzU29DV9wccDOd5kp
ylxdQWt4fZPkggJPiAgR9gqtK3Ob8xF1fBC0pW5nMKmVoQkW2thpCLxDneMWdSO1
NtpsJcSHS1pTHnk24avemFdWXFX3zxAAKUMbadDIZMVJ5WuyzVEGfl1g78eM3gXN
VXeoiqtZQh28stXTJxwBoBjZU/gWeMk+MbEGGXLbpLFdEnNUiHTPVmY54UIx7Ewp
KVQFmNGVTwEiavBDw1g/6EFEpZ4zmhn29XedSN7awehtz16CkCWXBttCSzWbvdDs
sfpTphftoPRg8VIBr27Ar5Z+JYbHyU7yNYJk0s2TPsIwRZq/8KWOdF11w7Jy5hhh
eH/4PObyNr0bS9kW1tCo6EmQnnE0nNKEDtFY2CAGYkTvPWoPK676YpW0zDJWp4+O
yhzmHJVi6wudms43IndrOklRR8copINqbSurIeXONoiilo+F6K175DwAYHZDVnyW
wjkKdgbIjFZkaNVdAbwoGH3tFmAASR/0rnlzSasrhbPvLpuZCwA6ipb9V0WaaO+D
hFyD5WACVeriOsxIFGE7fcreK5eH0wz0JOohhX8BQLbHnp84+YtlE7xx02aitlAX
XcFQ3YiXJKEaK6hnWuxNp7PgoZ4BGH2SVgqbGyr1WiVTwhaJoT/KTKO+zC/kZZsC
B3kKRcIcD8ogmok4gB3LiAIeiI8i/PHVw1fXOoGi71VybQAlpGW8o4+KxmxbIUIY
4tACI+PCOURCk5pdFfV0rHBA9OSUDegmLa9V7qT3uPgJQ61NGK3rAY5k/7d6t7Xr
3v3SZnbpL8p9nJviMjgTKFDjpi9bKBuX8DcZ7Z8KzuBHA9Ob+uNx7R/hfOwEDTvz
1Te2ZTzLux41B/BKIvUBfafzy4uuD/nBmQijKo7oTGyPtpPKqjBtkMkSgEEOOi4I
WT81GRRCEO3p5icsU9F+g9vezg60+3369ia6HFy+wbs3r3OmTCEBbaSY44SF/ZQy
fN5bJCZswQPOTF0WTk/bHVjPvoncfzzF2dFLKWO3KkwddYNCWhrUAXnomfSPJCeU
nyolBVj2oJJUNIkEzG0easQ3raRvV1jg96M1+A2E+9rN3TSe5lpmc8uQFdbUmLpC
HwD/3DxqKlfnxw9qIbG0oyH5DkhVuum9DwPYLTZAJmQalJtvL23/X43VR63t7kkF
V5Ey1APDc9AHhslracKE/XV4z3zIN2V4a9tkP8iMwUAqvMYLgJcqNDitwyHcU6xL
0QWQY4jiInEXtVq0sN6dX6Cj5iADmR5LjLkiRzKDFDFBtg3P+W4DZuNrQO58lzor
K8PADQgCdr75nK+tIjL5W/xM0+MpUIMDF0/vbdGEgmnvL0iRM9mtlgLgdOaMfLIT
I8ULMjxDKD+Qn3+SblTyw9xE8hYNUlUcV8NXEe3E38Tt7Q81Nkq44RukF1o47GN3
3IvF3de+q62RU20mV2/ZfcYgTTeUAw0mDbKMWadlURTTsYX6X3As81GVXOPRNyiS
+SwmuNoPrqaviycNzwup7Dc1x0Ep6XFuf55cuMgJfRY5Wg99snzWGTqrN31078My
ORxMDP4bYoe/Nh7iErF+vFfZKzo7LWAxraudUGhP+pAwxLCpCjOeQxJ4zXVXslDb
fXpzKAlhaOm2f8UtBaC457OI5/MsTwOureCFloPBaAY5vHKQV7fKAmj5xl8dIXyF
3NkLnnNbUQ7Rm+pGtM0BjULiaOAgR5csqynY/iRNhGxMsaGQLfO7k1XrcQQ8bhRk
3HMPFcn1UpCP4jbR3KZuInUZQdCdsMd3D8oQITHFiMUTqA0ynlFOE5MT1Xek71+r
v7yDkSQkC/DCSFEvQxoG9c//eplpxH6It+du1aha2Z6tnJy0OiVpsqSbmyYLn3xi
YojyUoHwhqWL2h5mDs8CFjvS6VY2BV0zHvzHuP1MzIdam2gHCWLZ4U57jXlGfD69
V0BAEjFZR6uFzF0mDJK0dyKrMaO1mkO5UxdQ74mLS6XlmTsZzat3MIBmM02g+VeL
5zYzdK3NSt3Y5ne1e6/63Hr4ENrju04kW/60YdwZd7vbHtJ4o0v4GMyagX4P4Vuq
2+aWYV8/iqQrFxJ2kMdRWzPvBj5O992A5Luukv+9LRobQvJDijUWG6XuIINoU8Q5
7XiNvBs70irF4AgnKJEsue0A86vuMbTUT5QD+veQirGwVpZxHDbS3a3lL1TJT3Wt
Ddy4jKJ4KdWj3JGM69/HEbElStIFXQ7EhTqc6pDo2k/6kr7n2ixlgsSBEGrbUdr/
LDz/4pkMA4sI4D9QoRxyZSJ4BLJLeVl7H8/4uOZPQBzH+WNI6RympIuiAHQES5+z
FNmETet7TTN5b5WOMUjuYPRR0vSI++zO8pkVSdw2J9/zEAUTi01MMOEVnpp3mwBw
PgBQ2YFpSglqPhGh08XdKnWAfHoNpWTI5yDiF9L4NKia8VVkfHFv3KIs6fXr8u/F
oCDg4t24Wb+Y0qxHn/2Z1gNX8l3ARELM/aZ0AV+sdrlC/GJSdDYf21Sa4buNiHuX
7yys39cNFM/idhx2g9/pHY9zD/8RaJpbImY2r9UATGnktsdihZ0w5kZg2Oh342OB
G7O+OKgKnFMPK7pawKudA3Z5WMZyDR9BvDosOmFwPjQrwx7KJqp4KK5QnwQn9pLC
0fhYyyI862A3okyTJWxpeLmEgPuuKq+h8W1+GaPRSRlvNuC6RnYmwFCJm/sUEjL8
dae6a/eBC1+lnc8oP24lEVZ4jZA2GIiuEyqCwgQ98xNE4b1xUqbIV6X3ljvbi0va
btfETHqZhjgt5f9yBsPxh12k02YFR4XhezzxO1tEhLf6I044Iq7e++yDSXId0wTa
QEujV7iab0fSRg5CPHa3KkcvZqwT5clzVTKi8kvxqCQAEcCbxZWmSAJ35A/sbVBq
92hmcsCx7SN8PX6XbjGYgmZvOdwAxyibQUGL1irVIb5H+Or7t+aeE49ZPU5On2U9
4nEGlc6ixKL9IKSW7e+yNvHHL9Ypz8i0Q8QX2UPlnUtQHB51IubcBqhnyTXSQtNW
/Lq55jIzZgalCL7yFsE0ryM/chfqEGetOQ1GWq4jt8bH382uxXtMhFo+sFoCyHQ2
IunN1FjvIuEPgajCFKa/PipQ1Dg+RwDv1aHDshn7GvvX5bbgg5RUTcfkgkaKA08F
eSMAtjwGJ1/LQYltW5/QC6vsXt1FtyvpffHLvF5FPShYpWDbj8AgAPPLaxgXI0KZ
Seo0HnZmhMjfm7I4riHM5K3ceA3SoGlP5Bvy6gWpWJfRWzbLpPOi7J+8c/WzhXOd
hw3vaSt+w+QIYdq3rsQXgIjQC3AlFwJctVupXwx4wRPWBZUs7E4XKoT3pfrJf0Kq
BDAdYucDCeUY2c7YlbligLEtdpiq/IFOREZJDOC/7091K5TKu0ump4/E9PHqAuIK
YEA1uhykQ4p75PAtwoCNFirLpFL54W2enbxZ+dSa2TOe9WMSgWZlcOc5fR0Z6Wq3
QP3mIeH9vCiZokh71K3sk788X6/USlb+wiUj2Dtdg9y8ssz/9OSYdklcKEtGKGJK
brvusn7hmWYXzPixYDYGkgSF+yzpuwa7r/KJBoUDdmyrK5kEiqvT3aSsRdSeb9LK
Hyw1UArUGm/MFmEcU0Jf6cgdbP8KbZnrisVfjS6WPpr/iP7R7XjtFBNn8ItpYjnZ
ECEtQdezTe0hg7PyLnCLCwm0PXQbOEdMg7MHRZMttRf3vpqfG0EA5rBY2aqcAJO/
I9ZKSJ/3wqfabD5SU9xLn9nqIKbK8OLjpQ5yOh6Pml7FNytW2BKx8cDah4p7l6Jj
CbtDnJa9KMXLzcDzvatyk2wdHhAFr30ammXJ19fJz+F3dRX8PkUQ4K1bxM1IwErT
fDsnRwkWGbUZVW5GJJKnd4tll3EHPg43q+XZ4mZATt2CxUmtIQKxx1AdAvXvtNO1
YiOfpUr2xb3eFFyS0dtbpvYYsupP8wWgzHQDwmTn450SlZDXt/vIH1kQX67Ls+J3
GW/XV5THrjTK9EftPCFXrzKJ9DKapI4iSDZEsDvmJZe14PxLabjL2PJu9euxUXyt
ZJO0ry1leA3//P5fImWPFgSaNsIE9BTgdXOEDKqgCoI9h0XZGDCUZ0gVZ1bQj3Fz
YjW0pB3PlGogN9qLBUKn4Ag+QxoUDlQOtW9CQR/5ceuTJbyeMibYVmL37Ew+DEnm
E0a6xpzUAkxxXnuppVP4QfnvjjfGAHFD1HdukUwBq8/cj3h3dg8gUkTcltR3prlS
tu4NPsOA7fP3XYNEqYxjXUjzu78K92ztSiDVENwoAu0MyRvf9VlDN0dAJj/yCIYU
hcYgVf3M7wqvg5KNi0jjaVvAk9R0rwGUymRyQ4hsqu2+rBT76ikJTJAk7Gv9kP9U
02xdDDAXVeiWw9TZF6/P5AmbNKABF0yZOYu/M3hiLIDLwn+fuPVqHM9Bigj6o2sK
E7N878VRewQpnnbvnmxaf9IhlhYHi3H4N7VfcqBXt8x29w+V68FQONaVCD0V7/gN
ykTy0tG7ohyqw/lFuZapSg4hn25l36d0XSxZPr67102sRSiINP94nCkTIyQTF/r2
im15LP7kWgihyW9Uv7E5Z1XSZj2zd4+vaVssckiM6zqZubOp+R1vB/NO9nNwRvYQ
qUl19ygNAJDaQYfAr1Pg+k9ZtdF3oUWdr6kfcKvlHyu8juhEZKFZ06uUfi75Dmhs
mVrchM23Xb6kNZwG2mlJn3F0ZOUkj7pMbyByW+UrD8MjzYO1QJ8e2DmG1hHal8dm
7Du2BNbUZgCeq6NtzWaNoZGbVySwP0jfRDFN24CMBGVkEgXEyybP/o5SauYD+P3u
S/l/9HlanukRFr11/L466amITqwnhPirOkWe4fOdt9TYu/C7AmGVM3tXdgUyURiA
H4e7Jsj9wltMWdPPKH3XKaZ3OqRpN8jIUOEqkPokLPYdkeebDKPqMltyi0rfkX5Z
eSOUn+Ib0uCmL905llP9PqTBzix298of3rf7J2qBnRoOe8PYkSWXSCX4/qjjlGOK
PYnO8n/MDHc43Xr28ow68QEinI3P3h0DHkQGHT+rkYTs59ZhjvESeI/ZJG0KyLpG
yIyyjzH40Jkg350GQqPIxMepwNYjruFdl+vd207MpE+etNTgGoFSnPEmS0VtQUv3
x9/+QwtvTNgis43fBB85Opb98MuZW6aPQ86jBGSJtpOTvPKkFjvOwpCYhUjCp3LY
RLiMe78incGuLKm7YBQUTxR6sKjxCOtkhtRc+IJckZJ7AFW7bhH2jzYEZJEbo4qk
FOeaTyJdtkkf0WioVnQvBw25ImqXL25JMrY8OLy2HW93HBCgw1aamlAGlGHHAFEN
S8G5ZbtOCq7IrPoPxCzIDKb40PTGxpmZXhjY8Z+EBSM7s9IlH0tmpl7BMpOTSLHx
TefC0HZCQRghz6JdrfUcKrjOVBaIqp03XceJQJ37XlHG5Vy9xExkLVHhPgoGTJNN
jtcvhPmDUE8GVHguvJlFIBKUH6FspBL5Yte9kF0uw66hP+1NDzNFzO8zL9ODbFOA
c+IBDAvNvQJ+YeCv8/I85md1VUeiulRJti4TuCOLAqe4cbgXvuqoxqmXLHaAjWNe
AV6HpHUgLR6T8mYGdOOSsdjJIwnOGKqEadihamNGv7GqchSmtjOs7Iyao+Ku5+SM
P1MDqJp3d6zL8o0Kh8cr2zyQn2aWZ58BlLYWo1gSd2ysliQ3BFWXnfn48esmvdiq
k4wAMO3ryHY3rwwgfHAHn7AovxuJRfrz1qUVjUbaHzDo0D0fwlYKsrzk+dyX4xlS
L4f1uEhUiSfITssr0baZwYEGokedj3e6xPfFMk0NwTW/2U/W5qKQVCPylPWyNPIc
GfsRS8/fUUNcfpm/IosKP2jDEjCUMQ+NE+mrFlgkurD7BTbf8a2Gemrh0uv1TOor
rwKGAeJ1xOYrrsr6pWkxoen5pGmVpxcp0PInnqEIpoflvgh8jsy0uv95Uq6VvrQB
FzyvFxU+oN+swZ5Hvrqv9RPfxYlgxCq5VgnNB6vcj3foOOHe3GLSYu7UWfaMNWOr
HouF3Z6qqh3mM0Xxgsg25BXen9GKbbFdRsKNl2ahzIynq34gSoKQhPf2CLEfYp4O
aGMB7MwQKJyCpOVm07dEfjJIjDQjhU7syHeCwIq5xIJ7j83VZu6gVmv8Iw9q3bJn
0jb+dHwm0hyMjmYa8m2oH04NI6yTVSkyiPEkqGtMItR2q6j0YKvnHpLnnfXlbLRg
L7VyerIDbbeD3PwY0M9B9O/A0ByeZHcR+gxTv58Dqzr5Omp4mm1rD66W+gcjLF/a
o5DF0DxOJIU5AP1jE3Bo1vHvhbuKxD3KLYw32YM5Pc6TjLugHv4WX4Yv2LUGR9pI
Nnqdi5ku/gCYsGeEy78Dfbsf1XF8Im+7GPec7a/RvE2tbeLMrymkQ2K7JLEhA4kT
EUMhJtVZdqr4EZRNV7kLEr6IQG7EhzOpypypNqe+/Or0F96fKt8vnsdB4nOIwDwI
7QkwwqudUuwkpYgCVwX9p20a+5uYwwkN3n7t2W9YhaQB15Il5MmUSTidpTFlST2H
X5P0JeofFUjOODejH5nGdEKscFe5qJRsJjzUjAujz6ROyKENo6xES8dPxjTuHmn5
TqlqT2KnNzJEc6MrydCpDbpKmIlWhK+oAZaN6Qf1553WpTo/TfhPZOxd6ReRVwY4
ou0DWS/qqITBEU7vOLoz1VAb9HbdJzd71z2K/PTTfIWloIN7mFACcay5ptj4WBo2
ceYDn4alrWVlvIptgZnO5dt4XHM5ZxbUOCR12m0zAnp1U+UDARcUrY5Yl6/FDBVZ
7Q1SXoFU+CRz+RDqOyjL/6ulPQPDwSc41Z56AU5isjSo2D4c8LZOQkIeA1anaGJP
VqCce5aEz71D+sgqhdwVLHKU6lBDukScenrEg3XRk2T7X5JVNkHGXGzmlPNHnQgS
n7gorZ0IpkCuL/1oXQEkqQO2VHyE0vDzaB8RSCwj+/T4cDX1VEbZYkhwutztCmXp
yPOINj/zfeYEFrf3ZrTxhYCUOhD1CD3C7YpjKtJ0L0bFS5AO0TDtprkaeJxbgB5m
FtWkSdbTHZ8LCDdH/aNcJnmUcrRAbMK0HdzL0tvZhSJ+ZXPiXrE70NhtdCw/gU3u
B1A7gQLHMEi0V+DvPBXGRS/tPmGisCWZxUE2T87Pqk/BBY2CKPB4bBZch25LdCoy
fRGvt3btLwfv6pPmxXKY4EP2eH/Mft6asGHOueDBAh3X2k6OXJBuKQLazhBrgGFF
yRuTr+VRrPKawXP+Wf5SD2CgXgut83zRmKeFm52kNGyw34gLV9sI3Ko/db3iEplU
XGPpQyWf9G8umxv65dkASFyIrUQ/+AeQZQzJ/nP4ECeTaUkUwhNeN8E+Dxio/dAG
pbqtsCu/zOgWGiPhas9fGzXutZqarpj1YXUc5loTLUPosxOuUj4OcoBE4+tXccLS
CElje27aveOYZEJMoh43xXoYJvIoohOQkoZPkcUf1Fbr7qTt+DKdtwOGbY3eUFL6
797wQcCpmIXIjvBXCm8R2I5/sgRvdu+k92eCy/KuTQtAI0Jolse4dCREG12n0t1q
ptTGgGbC5SFK5nYilBIz42hxHVbWeK4lHKj/1QF+vbm5So00HadwV3nw7lWGezlJ
/tbFfdaU3UfjiHBD1o3asq1Z1k2SUVXsd5u2jugFgKfh3b16uaDozwcX0ShgKSxi
kDuO+wptWwF6khvRfikghbQvDhB0sd3IUO/mh2ul+Q1Idv8odCr9LiKEv4bl+ohE
KgcFO570LINYJseYvWwUIn8AsdyZ/oPFcMb6rW3UfgjJFDqHcH5k8OI4oX7nPyxj
tld5Tjquvnf8J6xgVhxI5bPEY68oiuKv1OTYQ2uusn5rlflc2lIM4eM5L5JfVYej
kpwHzkhLFwFyPGf6qXWK/vy9DQKh77tzsun+gGFeU5iJbE77cWKXl1EcNps5e3M4
kRhLWxpp/yKtQZbqJnTIPX2eFymXvVnhLVVIfq6Qug55IanFqsi5tv3gaSiQobXa
Vw7nzOvLJx7JJqDNBj+1wfpH32nNB84ny2oxvj+uotiXblXKq8In+jXCVxLslxRF
nfswBge+N7EoJ6e+uNqOj6/cwDmV9EybStuN26wms7RmWavmCrKY5pDiyMGioTai
0J4rIv2uwHBs0/m57Xre1r5sPfNICDXRBPTn+yspK7BXZr06sNkLSEU1+T3um1yx
vsQxbnDtJ8SqIi7w1zwy6+/2NmGduwx9xDgcQ+RoKTbQtwo08Fy59Nj/BCx3R4z8
3oQ15CjgcHrrqlFrHXTd/Z0qQ5Lqlt3+oshUD74dsmwm4JcKqWpgWBix/7HNVYbp
T1IH506NFrBtIW0Vrl1p8V7HsUHCYveXA38PTjieu+etuk2uTgm0vzyEMx/5HkmD
0pJ3oMd1eOF/6QwiuV3MTYaam7kJY85tc0pVVzhCt5p7APFpi27Dq6xFmiRzsT1V
qauBTKc3YVqYhY7xCawQHzUbH2IFLZe72bP1tjbd+gskybkFPZlNkXpOgBugN8yt
9CsbbtPOtvMMew7RO7W0VRnKNoocgYZ5cmRE+dIiBIUi9Km3/OdCDme85nkp46TA
Ksdi3dxEEfp48Y7hQx2og4BBm58rjbNVIsWjz3IdOA/K20h/b6tpfwvq2c/8LQ0O
KQ3+RiBM4hcTQA+O4FyHkAhBep+BGIDzm9+rZYxW2HJ6iavV04oB+z3X8pHPIAPA
aabA8V8b5i7FTrzyFriP3PCA/APt++1j5Q1TyEzs+uVn/phwgZBY1KrzjQjGpO5a
QOKKdsGvpYYMRMvTCkWCUNNoOn3f44MNvDhvwY0E5wlgGK4/elW1APtZfAuzIbNp
P5ZVf83NkQLNlPGAXTUdzD18GF7axPz8LaJ9/3DC3QukjCCXjO730QyXrJ4cEcev
MoeaweC5avR4faHFjWdBr5rTCzjIA4ZnkWnSJx3JkEAzhJB9BhhROxHQAEQtKOqJ
sQ94jjGmYyIELsp1nEc20D5IiDKP+A7TFTUt+Rpph/4iyM4w6DDMg+7753/QEaZu
6zwzxa5kje6XjCYb/VWM0Wef3+EvSxKGJZrjcEZp6CovBvwgQxnHZxXYJOf/JO0Q
Cen6E7rcl28InclX9ZlwAAP7nBlYh8u9vTaPvyZ4X80ikNUMTBljXhRVmzvSjBUU
Q5JS3X2g7V362xUViMSCB7Tt/GNBPXv5VlXSRCdP9P0Tv0TGWLe0p3PnEniCyXoF
qPU01OWC155LNQUoMn8YyTdILPSEV4HXxel7BCwfXHW4R34649kxS17CirKlH7We
68twbsKdv1a/D+3Rh1iepG0H6b8AJjJkkZJEMGFeTYmZ/lP5I8PNRpbOXiHCa3EK
DAPVNyc6fmFBsnDWtwg8mqcDyF1RQJNT6O1AdyDrnLxcps6YyNQz/EBmt8FTtVMQ
P207YCw5hDG3IBRDkU6QxNsIa4n8zO4C7ah5PLU4kM3q2KcfRO5Ly3v0r9OLMAG0
Zo9fgm1aVxtNkuQVrQZgbhQn0jQpeiuMIskQadi+hFxxYB43w9abPHiQ47cCJAUw
RzGRuJGBGWv03GmhZqX9hdpZ2ilXzDXOn7gIlJ9i6kPVKoinFCVBrP71BVRBFnNw
Mjgw1MirrtYJ+PK8FTdVDDsp6ac85w0WJM8UF/3Sm5sPq4B5uAPf8mqeN3uA0l4Z
72DAM5ADm9jfQ8T3n+y1RWMsVsvzYGN4GzzFGkPM23ipENWVXg3scoJI/YRnuBsH
LS3qKdci3WaAcxGLuxLZkiU3cvZhgC6rFKZY1sqCBmt7utP707s1NcPULdNqC2Cf
WbdKsnYoOzPAtFwzGR9D+m1OJWeQoplo237htAE60eqTYwRRXe7vXXo8zTVVSZ8d
pQmsG2r8iRZ/U5yHY8rSTW4nE0cvgn+cXD8YCweVY7JgJVdjKmJ4nLoEvbMY0KZV
MRkQ7GFSBnsaTIv4hIAK3gWKt21/Rtry7HRsmsyTgLftrwA2bjvHguLmKF8zppIZ
QJIRshb1Q+gOXTEAo0AxDNGV0ZLD9m0Qten1lE0A/wHN4J1Fi/8IUexXWilxkvwC
Y47G6bJFgyxyn2LFb+U3x2joEWOYDiw78yfo5g1Lbf+aHiJc4fTZi/8ERt8/pxAl
oMIOKsEZwDPIHeANCUI2AFrnxCmKxXYIMbXNbFPfnA4mtUmV+3SR3TFFmQSg+g7s
iy1a+yCEox6CzXX3ZgM9ZzElY3FeplDFEm/XXzjdlaLyO+p2My1TwEh4nunw+6bl
Db0TY8xkfO4bIKrAEmkx4v3Fv5Vv5ostBoi8H5b5cRXI029QzovK/CVCZUq4WmUd
J6MYLBlEf6mNTXtbmEZFiBU9iW6v3ylV7rh5EaN689ZFIJcaPFYkYqQMHjo+BLxs
qDyMDf6c3e5S4FtjT8bx2xbo1iZXcfH1qz5sip2HgqJZLBWXrBksQBNVhM+LqSxb
DF3zs/A4WUBXkSSjfHdjaODY63OwiqaLEsV0lykO4hYN0VpNY6Mlm+B+ozyex4Ld
Abu80hLQ/GlnqT5K+e1shHrRU2+Xd2nocRSZWCyNEdX0c2UdOYmzZ9xVLZmJOnOM
FJjb2cqUKntZsZZ0gJzFci8DGV+oEJJtVkB5du/xdfgd4VLPYvd5n8lNp6Ed/8G/
QCvj7lsBYxPueM227jv+qmvTfOijbcaKe2JZF1ufz1nQ6j1XNiabVuZXKoQfKFz1
ZoLBrnlFPnDOBjbFLVITx6xvuEJLccjWq/ac0zyYpWCWp8abtazl4u40Q51bjCS4
L6FlNGi/K12TSwkm6crZeIRUGs5i38xGyD3ucRjlVJyYIFd/9wsanMeQE3JMz/Oz
4Sp2MRArIGMz6uSk1/QNCTs7WgIVe5TwUF3YC6rVNkALz3PnKPJD0oE0yCVa+/DK
V4JLWuSFLCOBtvUZMyMNRRd+CBLPr29zGTIAACUw9bZAbIms6cpCUU8gpK08wuN8
OvT/bvbcwS+nTSHmsbVXJ58pQRb5f3KT7tJkLJuYJsUVVNfCU5OdEhpDblE8tV39
s7xevmMVDHlMqU8B5WdYDM9EvHb998zwybHkbyQGWQvMdptZ5e/fvF/4/Cd8yOk+
EItwRT9Z6dh9Wfy+Ti9vOTX424sG/+JOeSGoAItcPbc3zt9FAtqPj7LXH78/l6Fv
wY3jLZenfKLKXDRAz94CZpBBQ1Ifj8dos2oOw+arUf4PYdTX0hm2Xmhv7fomacty
Yom0xbaUsYMQUrfKeoYPygsG+SI0ystamPwt5VXsWZWAra9JUITNY5QjFSmPzgZI
6Ktw6iIpUSx/mvegSxcxoqKsaNjleYzL42kqxurvwD46QfaCppT8vkjJhV5kAwJF
n6aai2n1OqahtpzrMhAkloZaZ+XuMK7WL/1puiejqJPencBfX7Yc7MpLchpaj/eL
VRPHPdyNr3n918GifhHcbIwK/IbZx9GhKdblx4r1Q5RYYmbko8sGIjw4H2mv6gn4
tasn9LozfPCfDxrdZGSKUQPEdBc9GsK4X7iPtI47qblK9rRHTykXAqTPZDF8R/F7
MdBCC/XCNIrf3VRF+uarblhOfnuZYGhTZFxGaDsRAEjcIjDEdsuLPQ6ptPK1paWM
a/ZredU2JE5RVXEOKn5J9S+Sl4KlKxHF+7rGLSRnkfYWJu0ihXAPF4FArFR2PivR
wyDnkQ2efljdquikEkQyySI+rgUqMAYlKpCQnm8rQW0V9iuBpOj5mCUYJeg0m6i2
qfqLoLpoA+cfu8GbYbKmD0QBwKOx6Wl+I95EoLvyoytH3RgpUeuXqWo5Xsz1y0s+
2oqwJAEPbKTUbAI4cO5y5jWu9694gYzTXu9u6Qev6ccbwdRuHGIkNNzmYGbnvf8O
LBA/Ius3ehCCrnqgRXLVvRcd1smW5Q60rEUbo6Qzdv7IuAIN+2DmZGGN+K4oSEUz
VEz6yTsRBvbCsglu3P97N6uCfadbPXVslraqoxSUk2TRFoaTwqiZ2d/caBiybZQ7
irk5+UoR1bLIIgp1ZoxJjf4ziS9TF6EFb7ShX4UDxGWm3upaQkZFxZ+TtoMXsSn0
IdHw1/JHBeuXr6fszEudRmoaKCxAM2KAnFs4DPfgJZq2rk5gcITZFeNjzV6QVe6B
lveAc3b1IZKCYrk0Ri10Lv0nIq2TFivNsftyaUEMt522D4eELOsUL5LLRSii/ZOi
a9TEk1PuPuE+4Wsl4QkYCb2y95IYnUQQf0rVxEL36WyzhiFkF8FSB/Gnw8c9zAuF
/hJ5g8AP9Q29Z3XqDnBwsel7agb2RQdkoA459vFVWGASXdtzd67YQXkTBi4J2D4e
u89vKnMyQqWR6KNdw3f6kVQBpolJpScJVAp5nFF/E2yTLKbqNcLnVPUpTyabZJlE
+f7Qrmx3xtO/SLKj3xdFdyDrT7tLIwvvarl3AW9Pmxm3cw2k5bTka2imWIamtME3
zlhZTHulT3bUCgk9yHCHRdWplJnXuTEBN5UXanFaxFxONa+/Yp7wf1m+LkT6LG8s
rNZR6KYBjpjIWNSvgPPVCgsPFIxgIkzKcn0kC99jP8F804ScPsr+26JeFEUKZ7fV
ajUKBryd1v4+4BxeHd3AxXKjWzZyId77lvT3MSq3hzCPqFuefe8DTWb2ez2oZFpu
M46IjnE12ak7hDBiWR1rLNEGM+YHms+ib0TX2UCt00N/DDdSXTrJ/E8pYvdrLoBK
8VD87EtbLWV7nuNZDjHG9MfLquteo1KEqS2k80gkMKYQBuXx7q0GsmXgPilpy1Xn
SAej0zOjgWAkJEJqbxG/PmClBqgvi+ROEjCi/FgidBdJgKN5L/eLC52EfLhLQH2c
3syqGcOOSIZqbkztM5++WFgmCb1TuXY7qNbd20fqA90mdRFAmDyHrtdxQZzPVy8E
Czfsiokn0bHZIMalnQ2WHABCj1wyyd5yh6lMQHbytKtP4BRu+byO266rGYZjq8ml
PKWNWlQuGSv90RRhOLrgx2ZVcEkNPxtWd5sssA3pzSwE1S1haYuU8blXgJem+Jnw
yOG7GFH9yzilfFd4323LgixkEX7XaE8yKAyewCTrE+gqStGt0uIur8XEEAYSO2U9
vbxbbdwMCbFreUgDjBltnUutMad3KiIc9/CgWomaB3LMr9hAborXS9+aP/qPvCx2
Jn2qae9v2MOK7eDSsz8EHMEpsPy/x7jlAo6umu0JF4jO5dv/K9NixoGrx4b+mjSM
GJIILiz92RXEz04PsnqpAF/AwWejpfuwG9GUpwlvUzBUnubNUXRkIhC22020F3ss
VjWpAMXUn2bP24x2Uo85r8fikAOqctluGVu1w7Ra7GcojUluXaDD3TCzADhEUWho
57Ji3rq4xJc/TeIirR5044HK4P6sDEsdjetUyQVisSEgFzSRtOLwRvKkPtzf+Mpd
wETJTK0uD5KgadBz/N8c3dELClF6zPFQR7xvGo7FJ1RTh2B2dR45EwD+BFIUqLo+
nScxW4dncjVgSSeAbNtJCSHnIgwH8Y8cBsADsoXxPj0O40++mOw5mElr+V+/AV+L
oAGdXnTgRhUe4Pghl6Ka0I304dEnPheXstd81zDmwkKeDgVVfJIbK3HQADjghj52
7Ymz0WB5R3HrAhjguNaMe0jHWS2ysjdGWsYVzTt0RDiOayJiuNZVA7n9AHMpZKgS
h9vLTyff7QA+aFnOh8asLptg0o4ZSlQP+nvzdbJr/mci3rCvSm2hL6UMsQeHeMoB
nMU2/CpW1w6435Q6wunj89DelnfL+JbPyTVvqCcuhhvtbZGiCX++ZcpZHt7N7sBm
fcaWmhYi/RCEsSn10CuAr826kT1VUs9SKhw2MRSfF2orRlhg4sBr9k35VAu80TNN
ry4bkdIU5bnRz/ySdXMcfK7hRgcfcVTGHQCTMUQHB8GOq2DALnXesiKHeh7flAjy
jBvk217G5ej5wFHCjdc2J8MNruOWhTfX0i0tUCFSg5NTJcPzhHsRTQdxXQ4/XySp
IsGnTe78ztsth6I3eBF2Df3pAP/hHahWPy+dZJIVdB/qAPblNylRBvYy/g1lDIqs
S9nBNWoxxj4qyLgEDz2PsA8WowvIzzgRaZhpTv+U9rDsOaq61101cenWnBM1jRgo
pk2oXSGjyVjhp8KXUQj+TQFQFV6TwuYJQagE5GJnfWv+QDHDdSPoct94QwWMhC6z
/Nj3X+N0dO9yzJgszorgXGWX05W6nvoIqMAwHN1mB5OzmjoAzEjH6b40m+8LYLFl
T7J6XRZn8cZzTjzKovvLa0aL58GDbg3xsqorHZzO0ouXhp/B94Pd2V+IP7Z2ybQh
nKERHA+OdVgXwv/GgEmPrXRowYbO2CosgUKUeiuXvNNsk70B6rlDvN6D0EGkfdtO
JT8EKLXD9srkWY+Ezv/Mt8OIvrSME7WPFJY/dThxNaFtXierlvAGW4Y1Im2CkRXL
4mNeppApzfPkJyj8hDACrJK/TkFMoKPSLD59xHuUWX08ScAhh2aATVn0DzO6EZ/W
9YrylX4AtTtLtZgkNooGL+ECl1HRGqNV9yLyhSGf2sq/rto9k9l2k64/ORFKweyC
TbiAXWKdgFXjK13/o+sXms6Ah0Ypo2JtrhEqRbxJmi7w5DHQrmEEPhIStFOTrOEU
w7ryhfFNU2qAFGi8dSix624N1mEQoLfv6Y+5nZiQ2Vs4jxVAXO5e/ggf3zlGGnpp
w1moqkZr3o9dHOLe/I4ywbNnk3ZVQoH3qc4YrHMVirwL1iYQOO8ZuomBNzpa74jt
vajzQClcgYhGOCbfeSA1PqQdzk1jGYpATFKK8VvDgwUEJwnZi08UIqkmpu41sCZf
EZJU3WGt3LAwjgcn7KFCOqSsg2gQsftOaBUCLg6gz4D+hdDOg4Y/XMOx5b41qGok
zM/wTturxchCnRsRGnAJZMS2YdsRLDpe+L2JL6QUQKeGlc0UiN1Qw7av6si0ftqa
gMPwViRQRguijiyuazbYnJ9rA6lK2/GvBpWbI50qYyHuFl5aFa4+M/3SYFzt9zex
UY9AJ8ewcMwCNbihoU7LMJbSFBCwLbnHZkMrKiOGHJug5g3D3AT8lfBAovLGEup4
MNiyDpbJMmobG0+NLXBgtEhztFwzXp8dMAvpYQYbI7vZr2RIv9GYJb+4M2aFudFq
bBTLMfNYMVtneVWQFTVtjcTKOIW9e4ZqsQnMGbva+YKc4DDm39FYhvRCD+qHyYud
qi3T0HZWQCetTlHGMn+yvDunqxBe5BIcD5WEklkQuDBzPV8CYCywYOwcAgunYOSk
jNdYdlBXSat41uIPTgmgJSUNXS8JsUte99Bi94YuyrtUpG+lF8D1xnPwtVSzunfi
pxtKoy5/vhsDhaS6I20R5UJYBJUuCfLGZuuThZfKqgTZpCXYZonyP8WV1A3Qrp9m
JP9/BakvSMQUdpMC5QrQuMwFxPBvlPMzfML+xE0Orf67j1w0WwazbfPbPCQIj4+v
bS3/BOUvCuAv94Ueo2kiVbeyEeyd+hsu+MSxeEgIXqXrsqdtTu26iYs1/F71RQcW
jN6LCxMI5Zvz+v1QOxNV9hkctbpxcgs9tE+RbXNQKHrrScNTC3gxzY14Hm8wL2DA
dy6nRqRYZWLbvPZlw8fFegWRBuWyXYQo0mJkD7GgdQ7kBhyuAh59pnCcdvLfqZjA
RCKGTRnUV+thHcRr1BeU3jE6ZkyMUrfWV0Zr7LkfLUTjF1xAqVdI/DOWRmfPT5iy
xHqlEO8I47I7FdUMP6djCoN5aXaZEbXX92eY6I2UrTWidjD1chD294hxkEl8JY0C
LTYpxylhzjb617sPiSdhZ/mtLGcdOhPhyCHpK3qkal5O6g88F06bZJK2f08Hj+T4
pkgm+lw36cvtqq1fJmnsZRxQMY3s7V0iuwvvYrQkbrla/oHhKG2fhmSzCtuBVaU9
0EoHH+ukI2dQnDEz65NBfuGC7gM2Pb9UFpcnmIv7jdPlTO2mA+i3U5QM7FxxSbO6
MsjQBOyqEe5jI6MlbaKg5ZwR8PdRPvgaXE/OhHfYP0TORzS1OWvXonxNkzWNCW2/
A151sB95wptzkCyTKV3Et/O0RKz2k9FkOVbhReqXaUUxppb8E05RnB9+hNDoeW+1
1IOAVhTdljHYby3Es8Wnx6WS2Lx6SeuL6XbbI+aQnNdWrLIogbiRjbald10r7t6+
BvvF7xbHdoFQMMARbL9xhop6+zqGzcfTjT4/M56LW36Dt8CIdp19m1p0Tr5/V09g
3CqY8/pe0RUoQS3tsJxAdlgbeVI0L/LW78f2bXdpWRSf056qFvHYDaUjUVaMzPAl
OaulwQtCF3O0DEtjSkqlvGQzkxWQafCfAFRBebMgJ7stOCBbDDjaOfwWA68Pdb+s
MPYfERej/r9P/NQU6KnynWBUBiTxL29n23Ts2MkflxRICMFSxVKvqSepX1vYiha6
mE+L5rHIWv93fZR/SF4RCvxptpMYpMQKDjdIWtmR9GUeDQD3Z7g8d4mF5RMV6QP9
204Qcx1usO2i+hmD0wAJsYreUcoItnM5eW6bLffAgzlh3QjWjB1bQQ3tqe7/UnnS
SjgWxBShWN168hRJWh/ifL214+a45+RULu6z1qJkH97AzLj27qMekGa++9177yW/
bcpSTtV6ZH58KrmBBLnKcNSd6IGqqMZ0dyZyh/OnJqSNn7LkZfZT+0s2lA2/ZxvE
MyHvZAhdFuypb+Hm2tn5P3drzoqr/DwB5oVDSUtvSMdT4bz8zMHpO1za1g4eR74D
42sKuQ7nFBOLev+4JPVplrPkHoetZ9cF6cvI6urETatuY93CuTjHVntav21Y+Ep4
2rrNHS3Cw4Foz8Jc9Jmklr1bwwI/QXd08nNijFKEoBl3gUo3qZTBkI+BgasKiZKL
4I9cE6m5SHUqv8wm5UwcmM+q5OI7WkGUKkUBYiNLmL3YNx5i0J+otCcAEhwYxhum
BRoVCGGsdiLVrP0CpQ62zZl1lKLCPlYHdaw43YrXiztjIik6mU84DpL3478/aPiU
0jvzhD1LYb7kb+4nGCiJMUmWeqyQjSO8RSaZcMp/DDFKedhf4hZRyyMLvvfEAOUI
INQHlu/HfQzRdmq4K3AuFAHWwvzj/9ZRvbxcbi/PG8RQLmS5eISlQSeBtqK2j2HY
6YoX7HeAcgOVRGlkjSyCLnZV6naSpCcPSVryhI6kCK7FqQeQA0lfB2te3tX1bGYN
BEj305mRtKs+q2qzlwZRZ/NewgpzX5tig2PN6a8WfPolum0JGcYNXCRVnUlzHTEP
LLZYSI9VmQatggcpdbM0+uM+e1XMxPrCfMpANoPPsofdn+fhGLiNX2sMwP+XBfBI
u6QhOeyHt4d4tEU1cN6qmiOUut5pUxCRvpOWpe6uIiAT+Zwum40TFcbqM9tBavcX
rxGlqAC/BmhH1Uc1+WRPPz4az9cqitIPt3Y9K7MifzV7Dm+V6RTcmBn/mqABeoLI
kThBAz8KQZi+e5rGA9WJiZT4pSuKij0DczEEiT4rc7uETUvbNQ8YQtCZHk6sVnNM
gXwHYu/qDJOqGlD//M0K0/tzd1X62XO35IumlYfcz1lGVl1/bk+MyLHpgb0FBL27
V8HnIfNiBpwkWi3xGLiuM5TbmBKlQtIQDcUvGSF2wFoEjF2DQnPKfyh+bSN8lox8
6bRLNkST+pl6Z/8399OR79vaHjhCLqpfi2bMrE0Rrv2hPwjcw9X/WARH+zBzUYYf
9H0HghzILl90/6XOAkdseFWXJFZFIo6ZKS/NVLJRNMEaqd+IzKERzbACuCd/V2Bg
OQwD9XZ7SXx4lq8U475Mva6XSRqT1p3NZIYg+NWzhC3UzrEhM5Vb0JeZRJ9BDdgU
WnRQ2Fu48qf1tlTi0USMWi7OaGFS0cDJLh0fot+zZOpU7J0Q3/VJv4QGR4ZJkH+P
/IbfCNmrH8el3aUBDPdWwRa6eAYH57HqJ2rr+kqz18jM7pvBJpnGiGD2/bb27r14
97LjClIcusfqUNWsRz1kiOaatmt1F5yJnlkJUIAws8DQ8FS/MrGXVxi3zd2DcH/f
zFXk4RWHecBfPR7u0tZNZiSw/1Iri1JVYtdFc8m67wbm8rIKyiIEPOJaYldpnhoV
z9sK3ZHVlRhVU21KgJthqGzGbqHAL7HI8LL77qbXVaphpRnowHb6pIb/uKOv3roS
yUfU5H3JAPkHNuYqtztu9td6H8wcDxgreXUePQ7MqbZLubCQwzol6EqQIc6QGy0x
1Hi0PFHa3rtqF9q5ckl4PhQNcqvXpWgKn3XCk4Wldr5MmwOCsmF9TVr44DkO+bHE
mvSKkYv58Nflp4QdkMuiWYzaRVUY6f7frISRcCrM/lr68kC0tEkAfKJLbGvNCDq9
miY1LANVNPRZNzUKcIBVxpyvlLuaTxurq2kYaDDMtYOK0hWwuR/aZ7YVONCSYBvE
EMAysZqaEmP8YlgCNosEW7UJJUW91l8wOQjTatW5O6+UabwihrXQjHcWUaRMnfmS
C2XNaWLQSWAhMnNzlJYILmxWSrfVWHSG1VC83gNamX+aY1jTDT2AiHvVwKKBY0WS
u8Zz2uoRz3MzGFRVtGujH8p/ksti0Q5nJvT2UU363HJAiOASGTwvnXr5zihmVrZh
y9+xiWZ6S4gvF4wO/FN4SJRuvFatw5hVkMgOGFlI1p7Eo3/zXNTDdFK/BMzuj7f2
5pHcc8CBFftByfSGtaoPFIA+FFckAHQFOcMw60B55xEwtGahVB3E2UirJjgqT7Fp
05qG8/wwiuUE7o2qouJht8UTtFnOZL4A1oxnLJAPOmORTtp/QbjR3Fw4deoAlbSv
IjtMq0Wbx0PPpu5bLTEwrrHwCmlFVFeLRHHPJWAPYffgRLMWsOGQEAwBBw2NfFuT
03p811fZGLmnNzD5CRKJS9lBDIzNBCsoE8kGNMUPWM3PXKbeboqrlbjMvY7lk9g+
A/qHq8AXqKWOnIe1O4BHkATBTKUiNsPC/y7pf4lP2wPvL9ljHP1Hdj19onQgt+Cb
3HAnPg+qFG2NYecFJpOpSjEq1O6KAPr5191/4FlTwuQFcjIAgIovB3GXPduCANeO
qmZoRKHmnWlkkNzcmO8ds3IqqBFoY7ywDGRsvsOc+HeJsSeE6ybnJDBzxo3lNgZ6
osEk2VK6s2Nup0FgIANiog2Tb2pdwmc3i76HruglB/nnzjgpDq6bhNxf/etPwdNr
aygoYezb9FvjLoNiHiIPolctqnbmzRux+gii+XapQ9PYDs2lPe1wT2+JkvJN4nIC
pG2uOyF4HN0yeEklJyxOWOxdf7D4MMJ5Qgj2Wq2thMtMVoPaMRMITh934MwdJAnW
hYpelT2pMJrtAuN80VxHd6O8IIeiCBqky2en84Ri82fmgGYrdm5xrYwDkK5pT3ny
O2dAK+dZeIyD+kILguylOPTOpjy6uFl0knIXIrIy0q40mVfWn6ws2JAySnF5oAK6
ul0F6mGgGvb1/cHvhZiI7W4HC0zJUn6KLKtHgYe/cT2glxrPswWlxQFNpsp0ZgaZ
bayf7xgPqniB1hgffq8ldzjIX07YvY5eC6QStg2pqtp4DIZdJ0wTF/a2qYvkh4Oh
GsDO0w1j8Zxv07Leub/fUG+5VEvUtKeX1iV6cbjxJiDBee5yV620IOs5da51wsxF
YYhCno4c7hRURlyvQwjH7rHiFVF4advsms/7Yca/RRoInJ0FTKvvNQFtrjYb6qsc
gyJAX+WRZiSwr58SSj3XH7ER3pw2tU3LGIXRP75t/8lfODxeynpSRkk5/01N26MB
+ypsFxXf09OcBA/qVP1mH2n+uRj0yfHTdQ1nZ+pQpQUDTJkuGFdXQfoasNeunmsR
JnN4pmDz02beSQ+jmd77846UWWtva74CIq7fYbxnlyb7H8HqX4HH0C5opCQLkJyT
Cjhdicw2+OEuRG9CmrtMn54ENMoaAZt5StTJPQwbbbeHWP8Am/oT6qj48YIRRkW0
Tj0jxXQzGr2UawseIleZwaFqmGomUmgYUmsjzwcm1SVlJoBLNLXIO4Z2kB0dhwSd
oEmblmeIe3rDcp22V0c6dGR9eNFrMgHVK9aQ+CuPYjn9GfXN64NVykN60mkUpfFb
8J4CObsvg13Hw6teq/10Ctj70u0YLA39GJn3XFtwKLxirun6VBOBLYgaraTO+FTK
5YLVUyAk2kM9uY45d0XfTLxN+r2a4KzBH1zDe7DgeQ+fw0WrUVLZfB/iZ5bFkNxB
VNTLDBdJirxiugRVhtbIEaxn/GEf6OzKOua0TRA/+NbEqb+0JbIEggeyCA51lGL9
53UWOMnEbkYrJ4UUn7zCuGhf1ozqKOc9Oq/mcW2d9WX8AgKPnSkKge9CoKaWf4M9
mtxGz+vFSbixSH3ZQMoixlRylZO+rNHP+fG9U8UuvDY3nO/U2OjEJBo5n6sPC6o+
8xkh8aRGYUN3Zm5+hId+eF0E69tEV1vRMA39H+xMzMn89GMH4zuAkXarJcYq/NdH
tZInvqLbUoUDp/b6LqYhwE5PIUmmCpUUXH/irkmVtqcL+jsCW3Q1qGjKjV53O/lX
ZxWWOS4rbmOZLCgA9H9/rfIZypeWTfuneL+LwvsuAT085TQHlKsBw/i971k2M1Rg
CLMlH55wR/P3efjiZeyHudMfZ4KKZAAATKMhDIV8iazE582qG3FCo8BLTnPLUrsm
eCduLcdFu4rNbdEuJE6YolT/yiabPOmxWGFbQxwY50OrCMCzlYoGeg46u5Ml/Q90
NNMfe+VGxwsKxByuAnEMpz6umJ2wfLqenvTVHZ5+p1fZtxxO47sGYwIpl8FAnBt8
eHlJPD30VW7trGFNRrimCzTutfqyhUyBl1h9aD9qPzVnNbOo6DbUrxDfae1MROMH
Qc3+83MPPToX3BoEATULgHJeXg0kq86WhijwziYEo0fyEx+QZjmRO46XFkBW9nHa
RgtQ5mumKCRqgYlRyZhPQVegFkIoLJXAqXEO6UKTRQS0oUnuINl85bPkYKlFN4aD
V/hv2g0uWZDmdrU7Czqtsb/lQbFy3UYLZxvnyne8wQp9abjr4yUgESz8OprwiuFg
9HEEAc4TpY7WA7ZAlfKSGE5tr7bfWKj2mTI4ZC8p5iWE9u6vI/DDGsv9Avb8RDxm
chpZ6/Tk9o0H574LXfP8khlFBtdEo4rFjreR9wAKgT1uQ7ZukiLJnEUMHTUfWa7O
CTu6W6DpI/7Rfcou6m/IuQZtgVN4x5SsQkKB5nrDH3NTrsNtZBIeMt+I5mnFh0/F
4vcupTMibH5TeCAV7sxDqEocmypNAVlJ9SC7F7ubKWUtThoMXkEWYaiZ1QX1ma4K
HGRFh2Nc4P4T90T+/cC3y3A3dYfSroXRdFAu9CCMoGap3pZY+bpmXL0OaeNhu+Jy
VeXBwjVoxrXnnoUJMU9o2qPhk76kFMvFQK/Ievf791xGutoMrHXiGYWT1ZtNZjW0
j+Z8W+5RMJc+ZB9fV/6GAsnN04aqSNeHJbXikGPGXV9h+9VT87m0C0kmp7kYlH9+
dmqbHKIcCravTV+LK4MkYka3yAImbWfJPKk1PL1R60XkOL5yZJX05rt5LAVbths1
87fouP/UkYVZYN1+ea/aERJAajKyCxNMTnpguVHkpQ/9pKRVUgIdqc41ptrS2aK7
20RK0/7U1fD7tIDEcZ3SnhsbakzNz8s6oaw5L1DkwHn/E0BZU8mPY3qXnru9y7RU
ugue4EyI+Eh+dbL/Pd8BZYb0V+wh1H9qhPNGszds1f3fuKSY4++wLvBU4EQ+8sT+
fMWOuAFgiPaw+w74WzoiBTwzED51C7VGIVSFRWptWrAPuuup5L20tuiOEsEaCN6I
OiPhTrSl4v649Sny36kQ0vprnjrQ4PUfHiR5LOkxt++Zr+1LeT2rMT4g7mecAE3u
gEzOxbkF5fI4wDHxMduQAqh2V/1djYFBENnwEM/2ETYUfpqr1eGiw9TX1X4oGY0s
ao3EFUFOWGaXb66sDladMK/ISb9TE3YOMe7x/SkvrB7fZAgcySq2ewRO4QQwWnLQ
D5Evyvpse0luLNlpot2n7eqRsdIuwG54nfPB+DOI8/aJUJwde3UqYxQXN2NoRZTv
MPsss1fKi1mhfJVF7913MTm9z+Wi1Xuw9LkT5J4g8B49hhiH4bfAcLodknj3MboS
AVSo1HFZcu1yI3Tq5MnRCRoO7/8sZgUpnRq40RWxW8jOxPLUyDo74t25+zTRp6Z2
mFFRINwEMPXHSPx3pEQWjxKFGYXAz2VXWrbH8J5rXF8CzFMli+H6IuLbq+TEuJ7h
sZgde/cW8VkWWpm47bQAWUh/zObDpfET+U+8nDgWQU2+FSurbRU5JERcp2o97YSj
7X2mXeMRlA308EClS2KwNTYxCsFuRl72SEHsmDjhYkzrJX02XCdjLqTsCPzwDxv3
gIiYzIKpryYmAtHbOlLtMEUh6K0Ic9HwAG/rDPMBCTlKWBJT2Pd4a0lff6samdQt
9xqPgsM5SASHr8S2ZlS74teS5NVuh7TGkQfb1Dr0uXlNnvZ1Z9yTfbpTmx9WpRix
ED3qZ+JzO177aZW80pvGC+NkeSIKgAfNvNJt/u4bTZsiisE9ikwFOPw+VJ+Rzhau
pleWAYf1VWM+AapeSsRMqvzW+UmNrEQcEMwVxfS2KJSOukbipA+iuTlnEV3W4KeK
4hfYKEmyS8wczB0jRpkg5LkMhPsWT6U0S+6LiuJRHwT7GLe+OKeT7FwGQhG0nxBN
UxcfFFt5T9dqZgAZV+Wx82TXW7nbJuA/kzrHRQ012AaTjphXZtIDR7EtzaDmsJ+K
qNDVHY6SJbujtZ8xpccc63l6dIdkgOj+Uz2qLiUrmPq0rfh/jE/kqEvVF4Ml4ika
iqrFtV6hF3aGHVmjpR8X81S27DeW7IytcsLdRRnznWuaYs57qQTiai0JqmV6k8ZS
As+utjW4HPR7u2ORp9UKLAQ5TpDauS2EXsMEkFH6cimmkZ8CTZunZjrdPplANlro
UKPZ9LTNmMFPyQb7Mp7DMdD2aOM8AHbVAWOUlkf5VlJfWCEd4SQzrEH+BCzDt3ge
aMmABh6laqvHiULbqVQaZ/qzx/Ve3T1PD+3fvxHAalw7T53jS/pgvnxWiGY72ZCJ
NbuWuFnCm0pBn3mWEUsBXjMtgVsNApdhLMKcjYEjUYc6mU4CCCE/xlORy0npgkS6
TisTo4iJaQEiACdMWlBNcpbhYjFNrEbgUuz0rWJ9l+DuOKbFiA0lOhmSi7rMVYuS
G/X/bPZH69ZcEzWGCrMwd9pKAdUckTht3easGaJsDB74YL/sfVDpwy8OEGnhX2OO
llwlTLt9aNePVz4CCqkCyf6DIGySp2CIx1fPgFG+uPGo0rrGW4cH69ilkhde/s9M
2ZG0bD6bjNItgEibMOStCwwxWfDR5ZT21jZA7cP8krji3446/8sH4V5YCwVvTO74
pfnnqPEGcOyLTzJuaxOFBwezfzSRhYwxrk8B9Fgx77H+9/Rd1U899qBGrGZeKghD
FsxfUYtB9vC86G0fNUTwhigwa6o51IrrLQCSp8uik7Y0XmiAtDLaaD8wrxF+i4ba
4bYu8Sr8u6u0CAAA3MBjBg==
`protect end_protected