`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
IFaXCgmPXCdp6RyUymjEidpk3pC8jHhCrHKpk4TdzTOLhQKjdEV/jAje5pOHmWOy
tUOJdRqOfSEsdqYZd9yhcBl07bwgXm26c1+7JBaK9gXE/9DGuAESGpB9VEkeuLoo
5kdOToqBsk5FvQ943jzzBw0WbbP7yJWFK5/Oc8ZP59PiVOH4CiTITArsS7mzVEt0
ibaMUpULpzo3KEhqQH8ue+nG9+djNPrYIx3qJfYb41bJYcKO13LPyaIUjsRQxJ7p
eqYmS+qqoi6EKvJl7AmqLtBRC/yHGp1O1/pcu3LT64Sjafm5oO/mafGym2OvaFa0
Qu2gsPCsA0kHkVBmEzVTqA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="IuaDaeh4TBnccuSYYfnpqCcDjQ8OyMCoYBKLT4Bu5qY="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
GSO/8r2MdLu21a89JEKDDxNjXxQH2i6Inm609RP7LYEdEdtivfYa4w42pj6P3qQm
UNgthclLZ7fKxzvL//JHcizKNBMSsxBJwO257qH911tcR43lglSTzDFtYrgPFtf9
tCRvn6CnQq4+0cKJGmEPwJlmM1Ijeph846UteEGbP38=
`protect rights_digest_method = "sha256"
`protect end_toolblock="1bjaGR+Wh+5fVOrqHT2gS8wpttTkGADmfRGgWcbSzdk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
xRXUX0iPNhYTJISIPGoZ9Ao49teyFgEDM/Nk5BvAjQNxi24K6q30PDEayKE9GrzE
oG65OqFnNOyGhqKExnvzm2q2smlsICjph9cqNKJcrinUQYveJZ9MaprJNBS4wVqg
OjaCXv/RjOWdtIACqCWOH2Tua36+HbgziedDEafKaMciObKwJp8ZsSheQg/YUuwA
VdzEUe2OilT320oGNLO54Fwgq95gpj5xM8MklKOmkQJVMdvN8Uv0cXFnjnEE17ru
C8owotPalOr/F862cIhz0NiOvvINseAegL+FppYQO0piuH/HRATDHVC2vJq30Fh+
hufO4qOqPepq2RLCgeHenJ2lG0APFZHNylM6BVJTTrLA+LyEq5JdDEy0GuGkQDi4
KC6Qbh+YkFz+C5PQ0CK6FQ3e7CsawKbkyS40dwa8h3yslmNr5kIHrDwLdQo1sIda
n9xHUUrQFDIZmKR0ZqfCx+LEc6BtBe/DNxA/D14m7QXbxaGRUPyab0zwW3LAorOg
toSroLZ7KW/WnGGTOd1tKPuXUmtYx7PCVTcfhe3S4SQaWk4tIWG49NjIfBJ4xOQe
Up5ShNy2yhX1RM1bmUcLLaatGvFPyy3nQv8OeW9xxMCeXzB/IuhZ2llnKWb9SkkZ
zrhj49IUXrMhc+lMq9K3yWXrcpxyMrsHUnyFBDwpBg2X8+neQ3ij0QWoFPjNhgf1
F22eVAwQulqRLoa2osun+JxVlF3M8Qp/Pe5VLlsHvsAwghUSQ5wEXDJjjE9m6GKu
NEeklxD3oRl/6Yv3OBBdVj9szdbAWb5bqpa5mjoWiIgMDFFYegcWteNlW6BqLDSM
7tFdNLs89rLi5Gd0RD7z2C+TUzIAB5MfWSxGjuESVB+cXxIs6cNOO7e9cxvRrUOg
pX0FMnsPiz1kEfRzUbnxxGeFpRI4sg6lvHu0SKDIwzY7R6gFAAOeaOVVljd/nGtX
tkHNvSRA2qmlNef+8/agynNVzM467Mzbdys/7PYrK4aNhMPkcCuMAvm0fjRLkWTx
mgEZ+HMj7hVnPOqb8+JrTCCEB/0eD0JcSIFA7T6PzUj/NtvHrNkX+N6nqp8P857F
fHrW1jY7BJc/X3Jby1dlf2KpZOfFrkx8GeU9N10RLMUKGAoUh9ncQgfrc1l5uPgI
fa80RRzS5jIQyQN3tmXkE6cDvHRbyrluQbvLftDibZEjUWZBqbxKdLeaakqdfIRa
FSUhBZ5Mnj10g4vXZWm3+hnXCbEvpzAlWZGmgevtOMliy1qYhAKBVhpnyHR568iv
L146x9wTQYIdDUMikgOMJMhBpeZuMn74hYHN9dvs6EDPN3kh6xvxD5QVM43Bx25z
bE0drKUfyTIEZ/euYPA/+Ibgwnfelu3TOpv9D5kiqjwYgMP7jQA6a4KK2LmJfPl2
Ejvv0Kut3VFice3QyGvNbe7ZZC4grRUDDPBogYr7JHl2PfeYZp9Yqtk6Lcgql0TD
0piUn9zvb8Llw60OEZi6RyCPHZ75rKEqw1CSztiragJFUFWe0eTVZ3jyKV6rLF8L
TnZXQS0/zHdWkozW0sbJZyn6hrIcbFuxNpI3vS2ctOX/sK5PB5zYsZQT56unQ55W
5e+5SsrDFInjET/RV8o0rPJq8xuQUsQr0e9enwMvHCKM6zxMhoniuDmwhwUom/ME
6kHIcHhZd3rnL7uYQCLKYZwFJ7b88q/PR9OFy6h/WAYLsxeb+WNdokLLTyKCfpe3
mwLrrX/JPiouXOVo9jYX0cdmlPJz8WRYML73m7FIbIQMlB7cxqv1NtK80JPArnTE
lKDIYG94aTmUKgD/RVhJekR/7XiVxLk12m4k4uT3vUYT2OMU7rUbj7OmEOn17Gik
/72vUfad9JbUL1NWJOYixXhh4EZp5JJsNz6KclfmYicODvFZvX+qXpETcAPQC7t4
J0tHZCSflmZPZxTNhGwh1wiIh2dv9F31agkAcpAL6mO6QxTnCYZj65zGXfuy6qMH
KNwN/US3dDV1wGU1rTgeiPoETt8MVWem19IUB12/wbHbtHcHACiPqTMCemk09pB1
BV1pB3FxwSLZB69sEUCoN0jRIL1sJ/yTevOkCoqo7goQbjLm8EdT7jblCVuuTFsf
eJskNi/RNXS0gO0dnfc9aWs6yTE3pkoEIEE3kfUa0o5Xzd4+9v9JFwSdE3kDpkMY
vzYZl9l2CbxT+rquEJfC+o3SjzK5BL8Cp9VxzLpbNihGklk9M0miaued/i+LpRS8
7JFzk9zB7JR4gCdxGgCOgmb648E7GqbxHJrU+jzZXXy8zxWDCNUcPdzEZmEGLWrp
5CfvE1TPtqL5ipRakjKXuo7Jf7Z1vYz1OPhaY89A+a4Nv6yf2gzI6MrVsgfc8mdQ
Vcgs/YJRFw1YBzGZTQJWPF6fn+Gp5IWZWKQMQ/fjE8FS8qtQTW8PdglDtjVFJnZV
gOI1iq/DhOS7WTZUpXlOltn9KMqRU7+EHa0YwRaH15OG5678r9TJCfv/gOvY3Z+o
JLnLy7VA6+C1K36Gfxis4B3T0c7Mxl2qOHv+VC5TwFmDsIBtvtJgsqwpS+hNnbjW
IO3SIg+n8JSVpL/EF8nYvkd/Hg7gKYe2NqpBh592IzwgxwzWK8t5wTAOpssLOUth
jmCXGjDUYtG5TOsbeGWEKkGedjVhDMtpfxTjJchJe9ftiYghULq8QE3aCAf5b0eV
3Vje2wgwRrNVCTOvjfxZ+N2PDGLxn4e6fHpFvCATTpfOKXEvWqDY5sM98JZNoEGM
JqvLqzau6b5EP9s9ki/Hcw6S8YWJWxpkmSwDCA35atVoigotQwl8HQTLZF4Pk06E
KNKRQdMPKH6XNdJQVs97AWt3N6goiuifXHdb+4vMdagT8KdNvjWXLyOsJ8502i84
jCEFqGh8HS5DPdoeQmMr3f4T+2jyrTcwSUwWmq4RMW3SmbCnLSgxFY86XmORvL30
MRbr3oDXqgsXQgRxe2oIXsTmBWt9hvDhhYHlHH/85r+xdr6IsNQIPshck3uB5n5E
1R4/9tKkq94yyJgvPdWCP/uiIesEPRkHpZYRNHk+c719UhgYbDU/FY3FrmoiLegt
b5DtjKPPEjhLhXpnUssvSRvsEMxtvmOQbtKWiIo2O0oLeyBJNC3F7uxyXqzUHnBm
me8W8ca54zou5Mfg/F5GtF3t9Qp+fu1hNsUPS5hONf2DLFNAnGFPPMjnzivNMfZB
yrHF1Bx2AJ3IXtqWIhhIsxWXMhaxaGQlKeCOHKKJxHF9judxhkeCIRrXedIczkOx
eizf/abVl5qhfQGwoXg9Ap+IX7tsNEcanyMOvFzYVD+Y91GBlt2pfLmqfdAtvgjc
VJPbuvDqV1qOqA9R7Tw+f9SXpLPWAVuF0tKCcBnphizjspP6IWz5fLDaAIkocGZ6
JrsWugRmk//odysJU6r2+rAmeFv1Sv5HmrwHiHu+5hLAIv0PH7VjmL4IFuX0fbdB
r2vorH0vE/q9TbVdWVrXwW3RAzIJfi30E9OnyZpw9Ekg0a48lPw7liwbIoOclK8y
DwLsHpRvJCZsbETzPbUs1wpfxWXu/ntTwSTJKTFCbBXJaeDx7eCZTNdRMl2XNi5J
Rn7QzdO+MipjZYaYfTY7EvsshoIKLHmnYtZsv/eysQBhIkNnRCp+3/kcbgtrYaDq
u+EmADPXD36YnAJdNwwQwUi/RA1aavpnbWoDBBpCplyrDby1liXmLHfXw3SV7bze
S3DmZ25xYxSw4Zbucfs0z+ZwbkS+zmrKh/ftCwX4QojXYZm+j3u4xLJrtAUPqgKh
q1KToyncyW1+gw25KmyvfepuT8GO2HkcAmtcfSEc0P5l6NysRUHb6MOmP0Xagl4u
YBZ1RWBBalIxlHFuUjoxv/vRqyGHLxmeORJOB4UYH5VnIJ6NLPpMIyey6fYDlNTw
jxUxZiTdquT6q+dGpMHyrUjhs7prQrgQRHfjgNVXPNToak7w2KSHwP8xic46lsj4
dpS2vM3+pGmSEv31HIDHLfkiXnydxLoJeyPX3d7cR2qDlO1REFnaNt9xjMfsFLOD
7YxZt+DOQtrxvKli1UeXDY/6VEtNbpByjkXNVer8vWRGxKtq88VfUQzHbshmS3Tq
NN5G78Fu2V7o9kNl9LLX9nvVOVJG2YE9+NGtm6VR2CIGp7s3HrA8jfcXrsGLS/9e
hGtWANnICJX7L1MxNfRCNekU8QNmQPN/1piFhHf1Miq1YT3n339Dg2AxJk2TF1j9
gUS47dxg94umg0Gl1va2ZKhJ/jnZ/iO15N0kjr7emN2INQK9UepZRYrrpD/n7FVo
uVfNeEMFlABdKXyoJRjs2VF910Jd7UQkd8mjrD6/DbxdZ2wSA7A1vZNEGCMBG1hf
5bD64FRaOEJs61c5d2KVbFVd8HphAdaGeYnRVjJJ2FjweASjzMdF9TS6zKKSaPh6
GCIIsoqp+HIt3gptuM3TsbV2IvHxEoDUbYuTJi7yEHENN+rtll5fdVqJXo2p6NZ8
ZTf1dA+7Ic/1YUJ7EvqGVxzb1r82SAIVXXEZHxOT4EDMJK6cM8el79QVRwLTZyOB
sKh48T+KSD4UhAxYi86bh0nuQ1FixC+RWgZnPmoTvPN/MscrND8xe9KhaxUIJz5M
2T044M8pGTc8FkZah72aIG1/FaAl8VPgGZSbjRb88dc/8C5+77T90q47sSN8qa0V
vIcmKwgaIAEEDQrWudatcOcfxzkM3XXYqE5tiLAJGfhSoDOL8dJpUppnx9lwhEIm
BEEbaR7r5L4FikpAlldR5tVU26s6zNFA6YDAbZZoOuzONjHlLf7GprQl9WNjFt+4
VSUpAMPcPwcb3u6jjrDVgB7fXxCUeGaYYwWIwMJA9sLE60/JftftWv4E1W0kOfeZ
5OnXHwmNc5NU1M19Y0KNi2m76yakhe1r+YAkx69vOta4sa69NtSR9IPJrnRh95S6
BxksX86saTtTK0tkBZ9kKPcnsNzJGrTDId40njc9F7iFVIwNXnBdZm7O20sO+T9S
xqYf9x5YyF4l5OED8WbgLrxIMDpwjpDd5ezR0uCMD7EZjjqB6SX1EGUmJ4yhNPXL
yz/bY2Lp2UuemYePZx20I1sz3ynDRJhmRD52vuoG/IxJcbadQCuCOyHaaahQxI3o
c7+9RtOVy5GQtOqGEp6K5ap2p+ANu8HkBh8z/RnIQUcPyUMw6+nvv1yt9QHg2NTB
arBXW59Ijv4oTafkd5qf7LX7/NAL4naxL6ZH9Qs3gqfaOPJs8+DezVuuOXQTgW3P
84GorU5sUdXUBTHMHrlB3a4FzqulNISANY8rkg9vCjXqfNksh0QVBnXFTzcgsnN9
16diBvMMoYhHNLUErkY5o8eXmNLTzIyJwsFMwaIJgLX2vkiUmqzBb3DLFdPDSOUs
PusfbayCjeX+jtoWrVU4aXHXn0ih4kUKBnUvWVOdcnZfXd4FELE/rUPa1ph8kSaU
dPxnZILnRqY4VtvohCaU6pNX2v3r/K8XEPrXb9WidKwxJ1wtHG/Kj4m5Ie98eoxD
bCKKJj7sHnqzvsVGsp8b74IIZB8QV6LYykXElvqI0DfYxVHIpO6fmXQN3wQy/qq6
en2vZivhbUEABrmHrMJ6DmV+h/WjuEQeLPLQJ+5bYh4PzcuGvdb+v7DXzCg/ifVC
0doTcTp6pK8K2MEIUIs7q9vbsbckoJjcMX4zKn6hcrlBk4cWTKq8Nsb5ccE5Gd2z
J5NFm7pKah/S2HPeD7u05YVlby6VAGGybjz33Iv1OJKV+GMeEuOqbfxvtBWtrRfd
sEWNafllzBepdNEpQb1JTSgLzpuzaFvvH3/ZTRQ2GIGtkVGBRdlok+vK+iUqF7c3
hZOpNXZy53arZS3wLw0DY76YHzRHY+ImHCtH0mNZ3tmmuNMyhq/DIZOoQrf6jKhb
UtZlLLlG/nDCutHQwZBMqUKBJk/i5f1owg4/Lksn2gcvOWSwzVxtNm+QMa12oA/5
Jf7fmeNejrLKu8v/4P8RNbqFAJCX9PM7cRGbsHduScEx942DWYgfX2jqQAfWnSY7
vF7q1nlTeli1sUqYe1+CtkgIHWQIGQnGOSbhLbmTGJlGksXNxuv9XFl9WgsyntIO
q9YBRd0gSfwoO0EXJNGavB+F2ZqVf2Wz9m8liNVD7KGnT26IEdBwRqyUbWL4BPzr
aKL5o3/LNbZLAcb5L+BXFoAItFtz2gQI9dF5lY19byDsh+Rt02dbB3vZCcfkkP63
LdLgMMawglVf+yWnInMmRX+23ixHLeXJbCHQ7uSFRqcWeg/IoTKWeorqWQGb+vqj
l73CuwKTKgpIXDRa+2/ObEr85/viwHm6X/UaT3hIjDCdEqIf+0ixXiK7ytPq/XKk
kOEDwjfMT/Rw+gRDGdsMA2M6000/1+TdeQ6FacvXOdLhVzWQh9oyflFU36jSGt5S
YolghvckRQ8/uaekaW1G1fZI9NKtKy0349Ay5PTrusQZUN7XOzkA24dHD9IsRP3U
Ly2B8oWPnYEql/AuAvodiBdBR9wBtLT7kDyuaZmIbvVMZZ6+JKM+oO2iSQNnHeeS
DU97ilNX3evrr3jEbA4zpBiJZTfi+hoKiKfFHLPJokxDBSwG8uUt0MPEgyMiBEl1
6t2+QFSI4vC4fCBmB+KIO4yx0eayZ+L+IIZUR6NE4GOpUhCPpO6bhSHDQMgSfpEx
5hRsU5MubRzfz2z7VBTgT3h4XP/QIIL0TAJy8urOkZiPyqoNTCgLrmT7l9hztqh0
dyo+hIv9U65TGVQiofDsWYbdLWcUs5t1hVitIn+lIoVRDzhE/YonE+ypbFl34A8k
ZucAwAk4F6Ou5BIShtQ+Vk2vpCRksu+eIQCGLMvEfW+sowVjFpmJ2uAzDz3Y3SeH
RdQ/D4I5maQsq144C8ShWWohMQfS+OPILzYJBdK2vX4z1BbvASPenQ/1yKFE9aJh
uZlEFF1GcXlyNmMn4CVtQUjFv+w/wIhym4Z2q+54B0IWSwyE3k8DuwWKhsfJZDbE
OAEUW2F5fhRoEZi+Poe7H40XTMVKaL/LiyImFapbMxp5qChR/fMYTml75oQ6gW2f
Wo8YCzvLurRQAjRVQC+Cg57K6Dow6N9cLk8fMro5aeSC3aHG9CVrH0C36E6F5M/2
WElzdsT3f9A7p8qGsNiF9GtylAa+DYY34VcRt4jJKXJ8IVgHiKIOk4YpboG2iKnN
T7n2o4xwrERunizlOal+VLXGMjd97z5zhEb1lzGEBnxEvsjYW68FCfBH8BLXuS9Q
SaAJQPwwOD2qFJ4/LTA3yjLKR7MvsFJr/Eq+Oj1qmlgrkWali6VkLq5QCkbdQ0gi
c9nfp1UPORaxuFkTqek6SrjTxeryVxwakAM2Lpqpunxm/DjsgMJerrz6tdEni9hl
iGYESWjqTLD6NOK0m2CmIyOCwuR+qE9/F10KLp7rs8ooEOrczZeE5lJYCdQ6BtPn
8nYqGQcSm0IOU+jQb2uZhUwOBL8r9WC6GO3bBCbCDPwjgXUqATvhJnpNysJr3Ier
XPf7vuNs0V8GvbPX3SZXAbqzKTYRHsNosujxjnOUKhUwTCQaThPOS1obORgNDXmi
v4ixJmbzmkACG0Ex49A8IJo2cNdTIqAwJnVlcW6r8+OYdAQVZFfCMmVPyMyWzvOQ
Rz6OexbA2ymP+ni5UYqQ/NTvCLvSdth8Z6rFbKwI9/ptOohC0ncuomiobHEpN8Hw
kvU2ORoYZuAk6wOiyeB+4E9bOUht1MPPv4s5j/fOJOOYQdzgljcmtbmySHan7c8R
62Vfs1VWO5+0wCLRdzpoWfUI0tWe/XzWZ7SOgJT+TdX6BcTBIKEy3vJ1K5zjt5cg
t1xJXZf22DIOe+e7Kslp9zgKKwvKL9BTZ6HL58oTCwUq2i7HNT5nug0VFmq1yVw3
i2zJ4zdTKR1Cs6wreuQ9dP5hGERAmjQvOLlMWHejor5NzdXgnH5U89hd99a7pnnJ
M8b/FfPUMluF2VKCg4yTYfqqcLQN9L7rO+kvTStg/AvxZ9RdL1AGITYaFg/Kha1y
RNX5E3LaZtyvtroGKk4KUSS+hkyTcklZLNRqrsIMT8MPMmrjsb9fBmHXYwvFZOOh
bGw8z6RJqvcxns7gSZY8Feu9Oj7eQ5KRJNjlhw1E/wDJ+eNgGbXr1FGBqXycSOtS
9OPqhF7oBLXgDW6l1i0pISVamS4WAWxlaz08/ZwNE2mTpSP2EE+E2amHy3NdvkY5
9cY3PADi3F5YasShji8CIG/ymFUTkLsXIlJwonv401DPHH3aO3QqYlxOHTQvLtrG
WVr1pBOWLXqXYQairgfhi46SsC0pfI95kufM8OsZE6nPeaFQgpSuaIgiijjvh1aD
p9+L8IGhkm2acwTlleZPt4iOpsxTXNkXU/YCkt6+lUZFrj33ycwxE5y2U7YhWQ6u
J1Htm1yQhe8VF5UulJzNYKJQWCXBO6yfeGdZT31W0NGosC195Z+7Y33ga/yIXmWo
yDFmqp8uqM0dwd5Wxd5rc9MTWZDLpDnZwZeWq7l2OShTvFWMJT7s2tRgvR3qqy1Q
5eVkthCApvvv1RMWJL26CrprTIXmOehTcU30YTsoltRvimX8gVB7+u2L8ZscBYGa
lyX/1sXbd0MtZfnVQEIapvB+yto0pMF0V13XqGd0/13uG2On6DTRFWn36OXDOSqm
z1NE+DcIeJQ10/a6kLYW7ukNKrQ2l4HjYdQhRywWEgo/S9gW+7u7RQOg54mj5+Jy
pIgWBE6lCeQ72yky8dqXGCDE+tFg/nrFAGiLJeib0KJ+5irJMKJ7DaDEalIIpxk/
LiOgtykx7ne8Ij8ligPUrIfmU4oVDm+50Ft2gCYeuYbiDjafTGjXDnUNLtHwO+nf
+RGoHRjah70PoM/m95Xiu3THYv7bUy/F6NHwzPy8LOYAIvnaoTrDmc9HVDJtRcD7
IZBOjpeejibBOTMb7BvPY4g05uziNy0Ht9TqLARx32vxW8mmc+H0mtcZ7wAzJdYW
cQdmPlrUTWQgtT1g+U9Awd0MTRpASwVnjSEUxO3404HCYOJKg8eZfT1uR5vc4Bjs
YrWccXY+v/h+erz288UPmvk73+mkSk5ndCjJtDkwYYnVZY4/NpM4995uyVc7pt0v
u6BIp61kGz0UjMLVHLcpS6eomMbLWphxFYVcAVC/2Fx8+NbJY8lXVg8Wh9wWfcE5
noaqvXjWVaaa0m2JIkc0Eh8c7hHqok83rgxb4GzZr4iYs8n7KfvatQI7x/0UuAa4
JHOp+igsUWv2nSWWVe65vWuBu9CAfrzvnyrOktFGJgv8V9sxylh0a9MiCQ6XpCio
lOtV1+X4Xoki0LeBbS9Bp2n9j/xuO32YvKWOIS1tyL7ntLHSB317Ta8mq81/kPGr
O/g7J8ZyfsyfFK6XaDgoecqbyZ0gcE/uMP+6h9sen8yt2IXWaX9SMMNxLcmxjct9
N+19nLHIRpFC611XHUdVQrG98SmOk0oBElbRiC1mHn1Ap8tlVcvJZ4BUyWCph2O1
cy5+mlBEdiCRj5nv0NgMt7mfA0oaiXrD6KmCJ0Lm4x3+YR3fYsLjN+JABN56x+LO
ECse0YbW9i8Gftzcq2KbJr+8VGe9/NT2s6FU2nzCPdjru4v2Vb0WasnYggfj44kD
rRhFwEC9TKR95WLNh6QpvHiFLNfcTZ05FNYFkrIpr2H4Q33mw4dsXk63i+XCJdg+
BY4dD5BK8vWZ8TWepTbotanzUC+CpTA0wma4L3455dExB3Ojg0NsuyPHatevLoy5
tQcyiM8XlCCbWP6uEOrNrtVZF1Nip/DpMYjWZLIegEAm5gEMgUTmboZYXtkD6a7Y
2w0OmXcPSpSpvcIgyy7TQNPxVdiLwdacAF6I0GoHKr9bgcGEVRWYMRj+6L+F9rIe
ohyHQ7vlhpp2BQ/TBh+2sZTY6R5YzGmYR0FJ+3xQOt9EWig/Lp5dR5EOO1wB7+Cb
5jvNwoTcbK/4BUZ7+mKOwIVWR+PTgFhaCL4B0GWKpIe3rXC0DMM+iLVU1O5RfW2o
rxDH8L1PWdbJxD4hL4BhM6gBBT4BYjtrNYIrz2Yb6rUIM43QWhah2XRhZhJsWEqZ
yZQaFUFy2eAfe6YnFid1HrBIuUfwzjHtsBF5jbAgH5vYmpOI3SqDZfdHz5ZxWSIi
iRwUvEjCwUsMcA9C5k0FuHOXkHDaytodVt+gR1dJWSu3oMdnrpRPqTQa0y07m5XY
YWAE6S8B+IjS8f3GhDObJv+jM5tsttyPrqa3YbzGTGjOi3/S9wenFLmo5H2izHIC
gEXgoNT78Jzg7y5v3nM3DyLa3fPrKWW7MryCzZuS/vCYHDz209cpTeuAMR3P27pR
hVwa7lt7g++gqn4HJTjApmI494QA8sa3CvHMDa4CW9Rs07A5n3w0PqOfrgYf7urb
f9O5NoxT52rU23Sg+yK8a5yZy4dkIOJUsWK48/n+vy93tgFkPEn+HWb1NilwtD6j
+NEvOGF54DOtXazvAepCciE8fboyeZiax2KVwj11t9X1ljdnB74V72o3n7/xnzE0
ldvOxdQ/qAcdRHoQTeDs5fLIcqYttgGRunJj9W5Tz94YZIzxwedZ1RUO+ZXISt/2
N+uriuoR3hwFegqTAyQ/gwGRrixahZL4UVqx3SDPnLgn518SMSBEwpRu0pqbA3zN
mTYRDIkv5S+P4kdd9HYOYAtN6VGDzMQWEucctWPRtzxNBbyS7BNCTmRvnlFbPzNi
OH360qvtxjYBKNcm3OyV3olIigLifqBXdFbaPpN8L0+2TPRKroA8r4hzGzUKYVTz
DCgXfz94Z4LpIy8fWJbtfB+SBKzxiR5JmeSP0Epg2UW0NvSPA2K92DescpngYNnL
bzztnslMPV6rQIIFG4MfSGciGn7HkIBmist12t+ULmt6FrgJ0JZgoqL3BDhFDlrW
QU36c0jgIrJKS/FtTRH4xZ3N4fzVwIt+0ZjBAr1Vp2LQ7InW3KYjT8Nes9aVYM37
0OSoiWg0VvVTCQJSCknU8u5N6N+8v8s/PFkNjbm0M8rtVoYvOVkgAt5h7KuX65BK
CX8MwnbfTVVwJB8hG1iiA4as6mSUagBOCF0MHJiicSN4lDMVUXbXJy5nT8cw0Axk
f7/zdnIwksDteXxpInOcLxafSNEnmIDeaKGxkQwvinDSZf6qOXM8T9HkYtycBTDd
3yGjVZ7qWP3iRt0QSmRLZB7zdgkllE3uuWVsBHRRpt/Kn5kSABByT+F8paAJR9AH
5WCmi7mTFKoc48cgagn0Rjf7sCBBHbiOTPVlWUjgR0SAGHsXDFgIrul/ZnR4v36W
y8cORDNNmwMnGflK+q/aIpDxtNAFwJadRCsEocvWImwWum/Gg4bxg3wVReyZfoKM
Sa959EfxMocdM0o7Kot006h8Z8PsZraa5hQsP5j6TLw3GlTYWEguK03AicfI/d8O
U0Wl7PsgzHf0pz+g0QSIKBpfEnqmlYkZvxVNSySMvh5G+dB+Juk4mk6yqYf0qcVr
8SIVCTthy99l/oT7j6TP0faqXYQaM+qZ/Qi6ikpmWhocohSg727JzJA9wU4FijJy
0X+x3XpGJssP55eeqVjPJA5Nf70EGs20tTnanEAjfak/5K8BpdD4eqN6m9Sm63GA
kUjNronPTTNgTRUr+lgBOLp/MCYCLuGpozuu3dvXkC91Hg3eUwzY2oPnp3e+KObB
AA4w5sW1FeMkFUgIUKrd+CLj0HGMo8yeK96VoiJ4kC3duBN7nu0YaNzupv4MX5y7
ntNVoPaunTQRAmPzZcxp7uTrrgk0ueRXEXyLjcg1HLMyo2z0irBBwPYZ5bOD1ya9
5+RFHRFASjznSPiRbUqTAQUI/oJCvv//tcPqFP1m6bybpPwnABquJBYi9TQ1kVQV
vrMeuzrAshneFCA+o1BVd4fROoF/fjOl/spNILX8bDqBp8NxbQz0tcnM++QyN+G/
8oSv0yovmLuj0tBih+ItespoKb0+7ib2uLARRaEr36CH+Z5qxap6wFr/ECB5uzqT
aXfXyCVyVDqv/8BXUj/g+bJtofcFO90bot6c4F4lbHFesKtCImWgjU0NYKDBOPXC
65M01GyfijjJLEr34HOf0+f7RScdp+wbyHkaU+AaifvfR4y/jzmJ4zKV4PQSiaVY
igHOEmpM1eG49o3zoXDhm5U2XpBE+DXvILt2wBOXJi9wsFwyHtyjC07B3vwqIxtm
26f2pN3Nj+oX8IkH6WoXf7+Aqj/Rl+C4thZ0Y7aaMwcaAWhaMl7U5HvdUh81q4MV
5K+zWpHHz1aaHSbgAsdHXbny+18aGUWHJakqoWt6A7QbQoVeWzwwA7tCTts9nOon
AOgmopuq+1lPscjMc+ZKfE2nArIHRmWxUX75HdPW8njqqDzpyHSUna7BPW32eNJm
8bszd4K0pi0BYgqW1ebiceqXHMFrHHcwv1ImxpZdN0+9toLA2hwVuG/MXL1fZLt/
1Sk/bi2/WHk5XjuvYzIAa4V2viiIigIwEbhjXyVc6LhSdRHG1JUEhjMH51EwNjxX
d9Bt1UB4vrH7/V4y75UnLQh6c0Xjy7+oOCIsNWKo0l9iE/S3ve6UjLiX0PpmvIlu
6szi/xICsj3iLt3X2OCN4lyFwJpKXA/6R2KaugwAtgkbrLWZD2/7zh5GbWq0ZQ1b
Q6UBxwHiHDe6PkVYg5K5S+tqXHEQIlZaZuRuBlysg61CvvKRGCuZaCyKkqn9H/sb
xBQ9UikybdfUumkBJ2PgGBGrlGB2OekqzsNqOJMDpXQ61fLyoGncr9D4ja09o0jt
SlwDZcydfOYNYtuyOSX9tTtiHjNyOdtksWmZkF4osfZDU4X7347JjN2kup8SSDU5
fHBvcnPGhG0cN2fBz6XZdt7p4u12E5e3RmNqnFs8Vh3jKnt9vW6NvkR+lSc5pvk7
Y4LIqODdCQvmQ3iH3UbTnM3qxSsoLsQP8CDCLWX1ejDm1RZWa+Oy0GvqC0OYod/F
ps/wsNQGhNOwHl2RKejohxjFCixjNlj7tgyUkwH4rkq6dEkNHM/IoD+c9s/B4pTj
/KIdG9D2QpPAoWIZKzPyHmyxvNTEKZ6pUnW+ASwFrtjvouf/BXVPWBL1DFcnA9tw
R/5pLDSKllsyBFiYJmFcKbpLkw8pVEPqEstYUdZweDFcOHMleCL3wgmqtanzSY1/
CA68cAnKeYgDrIB5h6RoeKNjqSQp+1w44QI9FF03LY2LkLQLoVxq/xUSjZ2JBnmm
GYCN1AySjpnJD1c9JyRtwYOqMiPkng6XJ/MLMSHfbh+5WCNrABMYqL+aZXi8LUWi
KsaJQgI9ajkY6FQlxWH/bDjsiJht6pIUvxWnaxqA+ffrlPioGDcpLt6zvNt0M/TQ
2O18TnH5aMn24FQ7s/x5gjDs4Rb+6+ENLCtZpzu6qI/But9EPouOba/JUGXxV7yT
b/B2iGebpqeklzjEsHxk1oy8lNS75+ByEIz74tC7NLZJ/c8IKQ0x8cfMQ3uilJCT
ZMYEag7wd7klKwYHdY15r9MIM4uaP/QscGari4iL0ZV9udJ6KNeyHkzgSfN+ThA9
7Yx4btiVq3AJumYeeCiUgNpmcoa0RvmSuxqCeVarblZzuyQ9sYEwlymJ2KhBtyoA
D9PmKQ4fCfFUSZA3o3e3FF30JunF8OxYm+3zCJeeDox4dD//l0cZgOQY+Qk5ZRN1
LtXu/rcmvbVb0fTkN13TRjdFSS6hT8ux4rwPDCGTvIbJdKwipAC7grWutC6FZLXY
kfa2ONbSW8t+N78w+r9x2PDUudvNJmxiN2VK/l1b79Q9sR3SeqH1soX11GT64TRt
zUorrJruPmTB47XxAQL/Um+nk2cE9xCz5rzv+Iyt92CCeqf+7apbN14ukFuQfRY3
SdJ7aaNwb8BFGEUxPcCoEU8wZxD9eivOcGhSZhAkh2WTps8PsC7C30R4fJpF7IxO
67zSg+oYqHuoclgu96NGHULCQmm6ugh8WzrPoHre7+gE69/42LnfFGM1j3t7W22E
fgLtXsLzrm6GPegqiBByugaadsrakw1+I0vEWNX111m1iiKGJYFVUOsiOwwktJ1T
NaNGtIQdP284mctcu3HLvneqyw2P7euL1yIL90DJrOdBBUr48rJnPEbzeQLOC3Tn
ShimIXayMmi8zevRYT62B1q9J9akf6BGFQpUX+KiLHlV1lJyfUn24Pfww9fY+ED6
I9nMuC4l8f8nu7phmhwrjOjo2k8B7IjIvecwzAMBeZ2e59IrjrX8LeybMcHGWD4r
/zPXH1mIVDeqfcXpyhJFgM7M7L/koS7Yuow1/l8/UUuVsQC8kpMLsiS31YeRDzDq
rISOyjGPFFNfbSQLBdT+JW8INFDdHSJMMpYNRRouuz6cZZFvbRR8ItlkgtSOPBrX
8BdTfZ3tE9z6XeK/J0GAjen/HWZyqtrrjKa6rr+7awJxwY9+lM+6ZJTtItXOs8/j
tRBhkBLYJYV8xPE+GpZ7jBnMZL0AQFsxoEojqZ2gHxHMhDOpGaB+VhGPV8s7WNJF
BgAQGS+oKTIDBHCwOjEoH5Twmmi8fIOCalhp2lzIaf/dmAh0CIy5E2nGS6Vco915
35cRYOJ9FO5PEMfCSlfrEuarfYFH+BK70wQAEaTOAX+4Z6dyJmV+w1Ev2oGnkfIr
qshVhPOScZH9FqQPP46wKBplp28zFR3v3xP9SzXWdOURltbPxKMFp9YXDWmdfJyn
WEMzmooZJov8AfMizLAS4jtDvW1lQlN8R5MtiDfLVcOChkg/IasdUGHaMMX6h8tp
mmbhynSaODvqYqOJRbrOOteNlr4RyZSt2ZuFDoYVH3RGvHhMpF9DBXAZTPpgtI8L
X1GlUs32ch2fZCHvPD2utkpvi77d5EK/BHrugNYY0Jt419FcKgRYt5swgq9gwJXP
ChuTExkvn6Wk3D0taOHHYbMdOOuuRfrz+QrejT+YcN/ZEW+WQNe+BTx9W1ckpIf4
s3JfxFHdf5NliXyaTgm3pf0B7TL3x6ur9wZD+bkM2X01y85AnMl/8sgAPfurxoze
WMvYAnBL6ADtPFotpuUBhZRjv/pU0FvClvt4ReCfQpXIQVIltcmIxBZt3Hhfo47Y
Rd7yGpxVlUQo0TEZ1nyZoXEM3X9ub7PG1tGKOaMYn8NalqvkRz28F2kOmVzeZvXF
TxOlJtdXLU7XmFbfMAsvteMvyt6UWZOe7bOx20tWWvputLynB08pcr6vO/C6SmM1
lluQjGkpGdTt8L83W79VPZw0lrzHefomEoVnHSgX5k37meBIgPf8qJy0wktKM9pE
VwvQuhBjropLeR72Fpdm4Toyvkg0u0sX4st1P7ZIYWPhOJkRCPjX8YUY+R9R2+gb
N46RB2DY3ddMzzfSnWu/aipf509Kvkukg5UZaAdg9DK9mwl8a2YEcc2WbKqSgRvC
6nmqysnauVfxwIfMcxooyra4p57Vs6fcQM2cfSfzOlKEMANP9OLqCf3XIY5azxl5
OeLvgVmmxsPQmnq2XQ1KAEyuqICe/YbXsbz7xb8ytnW5sRt8gS4eQgDTwUinzx9J
mbpA1ggPBroh3M1a/70ytpdAFABekeUdKUfhltW0w/vS+f9ocbn2TRTS9konyJYi
lq4HZZDB4U2OBPvmPUduaYz8UGKIhC+iF2QkYe/BTt5QvWUT930FSWlRC9W4/C1s
6kKWOtGNq3YwnaG5EW6SQ3DAvm8/E1vD/R24cFfXPpTYCrFwL6Y4OHN+NaDZVEdK
Bi5LlYljbKhqkirRVDT/0NG/BLThHhaqq5xPjnNnWGT91eygKzwqqQGODBAxIOVA
HRmg2/NSZ5qQJKFrve8226O+Bme5oqm8l9a61IpuNgou5K1A8GicLULsANe0fCX8
tHEnYsAjUZrcqwInJJadFeEDuUoylzf8JLyVzVqS1tDya9hrCI+BkKueetxvRFcG
t2qPhf2ml/EVKW7ic8pFWhscgkRSW1p+EEaU+LfcAiz0yG9eYuPelYbkv+Vpk+xv
AEX4o0i3OHu9yFUDaLi+249lQbNi/XFTlPOspC7fTRkICExh87nOJEY7AMP3I8K4
cJ2RniC3mOXnoev89GceaZ88jN+obpWwbi86zu6GRQ46Qx4aEXOqpj2YHPhuRjH3
cYF6EnflnlhPFqlT1KXUp6WjYb4Txpc58RA+at3oMIOXM+t89OAatWyetOgxtB/T
ULuIH/WEBMb1AH/aKuxAVarQaHFMBKmiiaIx7oeFoewFEs4hn6p3qU72i5BT5NmL
tGEyw4v+ahmnSf+Ida0e0fgegeAkBn9QwylWBHcwYDmci53Duf4s01OajDDdkVTH
oM0bPI7cWGKZDIwj7mrgjEmiuBdeyyA5Eyvn+18Bw9eeJKlq9wBwDJvgKR65dmfl
RkHl1GWN66NL1FCGCKuqhVSUl5mGD3yXiGRW5pOQ9tkcr4G6U1nPYyChC8kN8lqj
WTxeC4I8P453SbQOkGNMEgGprl3nm5uLUiCWIn6hPc4umFA8YjwuuqZovDrJFfw/
9XYfqgPUCIHMdGEUctBUSPrls6XFnfFP4lgIiHWqBMRfdMkB9IEq3VEC6XH0nsQv
A6TeuvAEr8R1zw8kHjsvIUoclAxiK85nprk45XtK3DJh6aSvq37M1CULcCbngq6e
NESEI2tjytHD7UQ4Kim0Z+EaOWC+huqAZ5Dpqu4H4IwPPTdVQFmKku28AJsJCxj3
LCv6GmAvq9OayxB7oAzPKYjlLmXavWqNBGVcyggzeSwKaSBurd84Ev6xyadUAQu1
+Q72dZ1g8R3alImL38jSE+PWDyAWFQhU32AJA1suSZg/rYeAPPdzuolxPnkpkjzW
XZvdeqPgTBersUdhzwaPglTf67US6qWHUgvvlRXse84YEEmgioB1C+efnACmlQeN
+m+BeIXrE4FUqsnf5iNY0EqX4Svg0yNSYtOQ+Wz9AG3alB0wX/JL77TCI/fBoD6v
3IxIR0iJT+EaCVSF4sFQT8lwjBmYQkNDhWiucazPyKo5/SkAusTa8wPDibIkOx+k
xtQs5JAcM7VdVjXpL2FiB2a+QRt8g+ACCDVN0BuJ0raYxsE7YwGgpbh/OGSVST7D
Tzq3sPKG35sh5Gq20m0MQHwGADlojP9N/ZE5hjXOI69E43suWBHHW9KoE6T1z2x4
tM+VnktmK5iXLQEWbNquJ/IY1PuSwr9QSx7iOxYIoGF7BLxMMFT9Y4OjPBltqUDw
LdqDtQ/Me4PppjsA7TrsEFGzfpuJqZHDQHSAkrv/+gNR2/LAR/AE0P9SDOk0sebs
wBtXEebuGImCbcsMbA7uETbEH8J/yU2aHKI5B5iQzeYEwhKy2nJJN9PAyazNAhB8
Uvq8fQzHaRgxh1X51JXCGRSXBO6oMDLBmroYc5lJvRxlTx5nn57AL+aD5AwznSdW
kEu2HtwOYBnfb137AqM8sFI+YPrOKylKo+RWHN3B+hedP73znGyQMWFheOv6cjUG
j/Wk8Ime+RonRVK/zJMwCN9lJYx/32H7DWOT2kH4ojupAhwGsUUJhfu8bqNaa6Qg
lYmi1U6hL7Cfw5vTiaxgV4UyI6n/lQTkqaM+/lUOMd64kMIThsuw4W/9egEVH3ZX
qqe8dqa5rkn+TlzjQWLgNM8fsB9yYwFaQxRsiNVV/hlGo2Tv1oCfHyUGoXL1O2zj
yy/wAWZ4jou3HvvWmlBKB1rJpZo+8+Ve1TtO8MCOZvwxiwcYNmNZ2plM6fFDdm2b
5XeKryDUQ2MmAFKtdlig+7J6ORyUr4d7Z6uVAiZfVzl7XcM+sLu/jAu3/cUkiVS1
gGkuX4af9m1Fcu959Mh8aXO91Rt3Mzn/EKyNz3lOHP/7mEc1cwOo0jljVm69M42D
E0jGpM4ZthXS6uGGAbBvziZ5aVvaAJPaKcLms8aU2tPYosYMRmJdRDaEzKcmaZif
zaBC75pSYGgv9nB7ar/70gOlZsG3BoDNhaGjOEA9uOU9Ku5DjT6/MdkgMiSpsk2E
r71EDV2jQLhLc0da8CqYSsNnCFXUemHQ1FSlS9nEaznqL0gDxA8heD358JM/ePuz
0LG2Y5i21ghFjrOumGF/E0EbVAzxdJ6VvMcKmohMuLWL1H43IssX7H6XsMQAfYTF
dgv5g0IDS2PhXQR0ttuA9Dm/InAEKGiJfHoMwgz44o/EaaG7q5ytYvWSmU2B+nZA
05pkyyfy1KXS+YWjw+woAPRX3ygjIpaH8YhM9X6ZibigajdPFVb5PPcRCC59W2OG
lChGE7ZjmtNZagn0P8swTyH5fxWbvcvB5CVSUwY5TOntorg04w8sYNAxFs9zclan
HdsUYNBp+vY9Q38kqBkRy3impCjg8BDMDu8coyAcB6l3jUGGkIVM1hYjidUt9CqR
5a9lApEJpx6eFUeMYFFxd3KdrJzl/MADku5FYOL58lrFztEQd62uom0bzf7bKwML
20H41IK4YFEJOIuXthp5g30w/2W71+FMIdiASZRpkno/9c5T0H+0Xd7ASUHa2UV0
Gwkd8q4Pc0l4GZPGK1PxirL9owpCQFMvTbmBwtMqhQbr0jQ3zbyRz6vUQbfezxTf
m5khQ7X8ANNRO4M9AsrCUPGec0/NAcDqbgFPJ20r+7xi8d1OhxxVz0tNE8Rhu4Xu
LatTnsPrrL2G1Gs88Ud06Rj86PDut9bOQXXc1wDa15+U2fsPSuI4Lqz/VJLcJCd4
E9FkQKws4d0qMYOw/cH5u+Qo4ZlhN/6pFy5F8RLBAvsVt7onjvLgEVOjDy50+aUf
h0b2yHu5cFV+nTdWVIekHfgsDNCBNHlLjWzLwm+4Ey5ObBFWm3Si2AmYNPkUCl8S
7G4iSyHOtvPAJh006H23RQ60Xz5xNaAU/LgD7R2f3Euva0Jmu4VSPqc+N+j+AOX5
mlDDH+yd9o9YEzKJUFArdRs7YyQixJPtove5M43RbwRz50BfTchQXn/DBz28Fuh/
Pni+OAk/fK/rCzhI+OW8qjNxPNheVp0N+552fK3zQ3DtNpVbblJnhGG5kp0gHKmk
oef/AYPMbOx5G3GriVejVRr5qq7lBCxCYg9Fv5pcDHqXi8c/U+0+sQTffHR28x7s
5BABjVJnqyjmz+AUdjbSKVMprtZNDwBy8YN/Dl0D9MMwsxALlhZVO1LE4ZcXXIUk
B2d/21iu/ve6X9LgDt8GvZkWmg5USBB+pn45GLRdVWRr+L50/fw2PiWPC4874t+u
MoUzW104k/pyP9HFtjmO1+qvbgH6+rIo8klR6YGcmF/c9e+IDcgG1G7DN2UnYYtm
OXHMfmP6Spn00B7fMR8d2+0JtTWRMUzDPkONCQyflBYblx3OldP/dIrFAxR2x7mE
zO6ZO2frw1h1sqInooM6LmiDZfGzsY0gkqEtU1Xjd7FPq9kIaLHS2imaHM+tugaR
yCkul/4jq5rBDOCjM8za7GLkPamDTVihvZeYXSxOWdM3rrKyArjSKQQFmJ5vOPoy
scmRimQqsn4dCQW57IRqDHBWVTIe0dveN2pXOdss+FI0OciBILVOjMUN5RstpVE6
NLi4SvObOiupCWl/jXQJwM2X+hFlhUXVhMmgWvwhW65PTs+Rq/xwtOncDa8l5a3r
xV7RPTaCsBMNVf1C/P6iMT+GiNDBzbDh3MwxL5qFrCac+uav6t+TsokGSOmtsf1f
XR+Tw/KXgSX+6xJ1Mrrs7fl0K2NC3QQlpkKoB6sfg+Crc1Qr9h+GrNPWay+zUj2B
aeCSL16/EcjpyZsPKNXy9xNjoWwaHurvZzHX1aCerRzt2c+RyC0wHK9FWRJEInHx
J22KVAZA/RF16w2By8S9Y7d9VVbwqWqD4VQbzxYD7OvYtBeHCZOAJft8cOU2nrDj
XrZuIxRKR/6cVFTyfVklxwpHTx9uhqbS80qkrC/GR8+rzyX0QwwLme4UPkjRB2C3
T+Gy+8531Dd/YV6WijKUI5UPD1N5xQxLOM5phmaLYTbL7lds7s7DtAsOHcgsv9kq
eLcHnApLF9ddUM8UOw2u/Bq0vffAxcjO/AzpzyL38IvAExW9i6jM7ysLGd4AUBcS
NV3VsqeFgJKzSc8fYNfRsjQUsbSEZGWWSZCAf9EqRpSVK6jb5ns7iSjODYiuf7Kc
4n2AWf+CwserGxDzoZ5LEK4mP69Z5oClJtqRJ1Oeh4fS+cjyA95R9tf7dajC5B9v
VteR/euRxjyWhOZSxLDg8raGWuR0l4P2f00YYSEYWRa/ivnzcuyHCmSanGkYBHzZ
qCgUVEwBpbbUrm9igqrOw4tFbMWlMHr2oKTcL+anzlbPBTAciG8snwLkg8gfVBd0
qlC/y11yUapi7rw8pEdqHJLl7UP5Qy13Wx35UZE4lLzaltBrtfajZUk7RaPvGcxq
bomfypJlaFBmomxgvypW0B16kYGLWu+pZ363+y3+mIbSYhd6TrrXz18MIGoFUPsb
1s9sVKOq7P54bYjW62MctmIGKfQ2FOBGjjMQBxr8qlcVd8PZF0mE/zvu/uv0GBIR
TV8Edbq+GDgS4qjGIScgBJE9CUbwz+G4httHHkNlZg/OKLCjXmBeWg5u7c9ESS4G
lZRBEP6IE1q3vtsa5aMX7XVkzK49hIvFMfGiHIa75mpJTwEx5LNsD99RNiUShlYu
XhoefluNPhmVG/HUpnwYwSKa0CWPbwl4wGnpHBhsvkOTllMsRdlUJchsHfjTMPKY
iM0pUY2UBYcW+CDl+sPHG1UAQIQf6pirca0FxwJjvIatlfEMij4zRpTPmamqGw8A
1ElwQbrof5GrdEsEJYITJnn4GpC0Is7U0xZAX8JVDoIooSyJfVT6hluLruE4gsiB
vs8TiyS1KMQRBozl6AOJYOFgTakBEc6KSovbokHxiwXJ+tFYNqMRUHFvbc09agPq
gbRBIJ46+QUMEj9RAprakVRYcNhXVdKCPpoYk+dPQ8kARpzZMQWzUZ4am+hLDQXG
7BUEefoOF/IOOLXbC75BP4PlxQOHgcw1L0r9cEW8woH42520eD7wfDf3nGYYj080
2HRC9vg0E+bNUSiIovrnM+IIn4PWs4UKVAzfqxg3PTTdLxeAOn3zbvDGCelkHOMX
jTuh9Weu8PQAX+uyQk5/bH4Vj6fRvyLMF8LMuhGC0bSml1HOe/KXqZ6LtIrXZ6o9
R5rwEY2CgnpBSKZGUBWLgiirVSyBWGB4QLL9n4WPbN7ivLX7yqmbH5aSgUYntVVb
ojSBh0ub+wa+RfRgsg5EDcFsQDIu0Qer9OAL9eZ2M5vKwctEog673VKTbXwnfyPx
elRjQ6oIqAln5BTbZ4QtHwKDYNAruN+d1tdIm+GC/VtvyhtfDOD0x85pYlrZWti4
1vV825ygE+oSmZdm7OWVuPYdAec0HAh063AJw4eMG8PZPZUuZ2/zfEVa3Ki0lBWF
vR4Eu8WKuuS4oVCRnKY6gcRpj+FLl+cxZYpZdm2iuBh8PoTZDxfCMVGYVGkSCJf5
EwU0TpGScf4BzZ82UnL7gxoDchiRMyMzart+i1xumimyyHQiavHXWyTLRRbnUEdz
TgyKD+KycNqchGqHpz2owUTG03dbE0N3nvlpWsQ0KmuoQHlW7TeSNef/GolMYlz0
NDaOz/N0ISrKD+/EMq6kDO+J84t0D8o7tOnFuIM9WTELxdid4YlSdLl3ElsELTSn
z9sTM5pK3V+Smldu10mGmBcxc7/DNMIIiReQeLpSPuQo0Oy/WC447GhR87vJIT/n
53snX/xnTZxlaCbEfsSaSgyDZ4Aj0bmomOl+rQ3FbxT5guqDHrvxE7lZ7gDpQU8C
nUtVxEZjzPMMMi/QOmu9tBxYZ8JRMCSQmRejhwEsJBpxyKtjprzN9BgqjumEGQeE
GgzLqsSw028sseNyVvkt3z8XKgLVlJsbQ8ZvhZ+tifGs9ZjczwlLBHLYG+cw7flG
KW5j5Te90ptYOi3a3nmCWdqZTb9KUJn9cWIqK2DKHlyiv2YlwrL53uFG8P6OeMAC
EJcsnDywkOofxXkzqNuq0VXptLNaYQtLNV/mUQbj0X423MFYDeqxqfqTHP4xj4Dq
mPVEQBP/G7jL1+KfM1sL2hpeWORuCGCHBOFxYxBJKjv7byZuV2WC10RypkCoVu2f
9wLVPMyWnL/gGh1IStPuyFH2rih/wkworp1Yt6q1SuzJ4geo3Coxvh/bfWh10Vhe
XyKp9BXcb0Akx1ySwhFOeVpdlcgF3FE1xhTg6RKYr720zYAy8tb3XDBLW+vozi75
FsY0ysLgH+1MfU1e+7vcCHZoE4s9ykJsc41cZf9G14F55uK2dwagPeokj5MFVYjP
fHnJwEmKAvNiauv8AzO6Hf5Y2VoI10oZ0uRwcvJeKAiFlKotcOpT0G+9oKu8WomL
y4RgGLrtJIvtzhDAdhwUTh2LXECw0BBKSEVXfxpwvntvGC1XUTKXko+IZc+l3zUC
WJo4T5jgPskJMwx+lCysZYko5GtDk+Ki0on/U+obJfmnLNz9WMCZweIGs4dXgIlr
XvnmZa35zNb0+6b9KZvMs22jQW13MVe01RROiCELeZshSuj6Qs2bx+3TMQTVWZ0v
u8YTZx3fpROl+6Rcsy8YEg4QKzj18pSqe9Ky2ljutzdaWjAZ6yqMGiUfz2kdx/NI
NfN1frigTF6ZV532QqeYvXOhudMIXbKe/ptgKSLvaD7hEXaVaqGfetM7OZ48coDh
gyYebFaqgDo2DiFL2mEVxZOGyhNCoPGsGKXS7tD8PGAaSq9HqxQH1xBvRgVpPqFp
hRvZMDqeO1ygBZsGwIIsfCHtng1ihsa6K1fsml94xhKQOoiFrEyZ3IyGGnvPrRmM
R6B5oJy5KdQJlCkAZp0rbAny66LnFldoX/3vjLBR7fmss206E3Zv/8gzCIfIpBi6
ugeX3e/IqKcsVf3IVlVpJ1jg0tyU0Jh2hO0qw2qRFVUkABgvmc18hgvE8ey0exMV
cJrpQiE7/SLhETyYs0XcIv0fmiMnmX7HahtxX568FVuKfv6rfwt6qc7WNkg12iXO
+GLCsk3sLMXw1N9D+PEigECufEfSF0VQaCWrxLQv7bOB8UwpHQfQk5gEAF5JCyK8
jVX4MwjDdwfR00f3jaPoE4SeW0WI1jiCD8xY8XFXyQx2QCGAY/xREXMC1AmDbyaL
du/UzAbxC0FDxZrlO3D1GDSFXMT7zZP+bMBI8WeSXFZ9ZUN8ST6VAq7oXNI7jhvC
QztwnlpDFIJua9PvciHwkSzFTdo/0mFQossQ50OD8m7ODo7vrt/tMbPEJrHmJKxe
v3Sn2GqyImX5D2nJbEpwE6iO9U2Xex5Q5dD1gZwIa1JrZY9+fK4zyweJCoCcTk4k
j8XvbsBs5JW3o4a14O+VYPUBoBeBtDryHKB+9lyNQeUPMD5M60qAQxb3Xjz59zyG
Pud/oGMbt9mVeJxgD6zir71C2c1UdtjOJsuO8pABqYorvsfgSGlUFT7xjqbkOXm6
WkVg6MxsWXpccSlLYy/wIYSTIquQSceh7EcLVD03JAzyudEgYqyAYg/2mYQhSkv/
Z0F7Jm8pKHdncEVuM84t1TZ79wWNi/qglaa94BQEMmIufhQNijcGwv/PCTwwCjWj
ekRtiShTqsMDAqazII8C+PNEB6z5U18b6aBko2zIyneEt46BJyvk8qm2fd4eWTn9
WbcqcysGrs0DEXfbk6HMwg76GGbLCmRL0XndYyVO9kHfySTkkAFWW7m5khtMP9Ec
co/pJeerz18/Oe7GDEOXS2eYcpqYYB94eH0AJgTM6e9BuIVNz/jEXaBPPK6blqP8
QiYN2c9M57J255nwXJ5Und8zzFKHsOfASKKf/6pdk0CgHU6j4k9xRVZwLMMIGfpd
dVV68tvIzDPezjAwumqu46N8jIGQJDJZSthafhay7FTiHdVsLTFvZf/FuqHF/FPN
W0x+rm9JawZ4oMbHoyrsykyhy67vAE//GzBtxcOSRwUzAT7AO8tKpnacVEaXnkGW
OVeLcotn5NM5RHtZPbOQpRJ2YMGtZ9ZfM27UDAZTsc8zVfESaZiOC3InjrcXgytD
kWMJPkWtWcSX/jXDVFpUA6UcYGELLb09Q2sCmt+ZdIJgrCTlTtWE2L+ASiS7c/zD
mEOzkySRFB/ep/EY2lRohZsWKTM3BhxPM+b3oTpkLYYlanI5WPvrTFHSQRiBvKB0
QIJQrhzTWK7JEExcYZP1oMd/z7mzPcYOQk7Kc1VXG38TqN/XgfOOVJ4Q7X7BOeuR
Td+WsqVbCi+kLzqWKPHFURIPQc3KX5nFm6GZ7m/3xhtjxRcPARZYXROK622zI7X1
mgBx9FhaLJVHjtTn3vfyKDKjZLUny8kHwXHXnnPrVlb7AAO3TILkXpH0+Sy2Kpxw
Ovw3WhnLoG2EynKuGXq1usClcoAH+gQxt9tn3QamtRfIj9eJj6Z3LycTQjKZMqQq
9L5i7luF9l/03GATV1KAEt5kl5LiCiDsAPlYff/7ynVS6DNtsk6ojrlNIPDh0SwG
mF+H1dcQs977l0lwWu3lHDiosNadqjYG6IYPlvJb0WmLypKvgm9NFNYhAA0juJtL
mA6PNoYR+1rbzRSqE9pJqv6ph3m7ptcr1gkU7GNdAoPNiCcgppmpK4N3W2EZCyZi
B5prkEg/N82CpH81nOAXHPfKbY2yki12ZYsrTUl2Ruby1fTpSAN5DefIEtU2+9vR
yxDoY/lpjoO4ZYGOFyKlV23pA0BWDkxoxlYifZfu5Dyb5EsheUO2qfBs9LP/upYU
9JtAGohd09QScl4mSRFFMl88L7xPAzTRZ153i+Db1kr5gtk3hTAarOJTZxpFCI9T
4RimkeKOOp+GMapajAK3nQbTKMWjDdC2ccgwYXGDb37DLq/1paa24KgtAsWheeib
2cF4Hn8+/DzzQpI7ciBMyktpJJPR3JoZONKbfxRi7YfBEjl5KF4uOiSz43CYLRRP
J2G/ZKqIK+k3M3lrPCd4rIlA4m4TtB0tBB0EM6pXa6BIT9ZZ2JzfL3cG7rHGwnW4
vnIx2BNmle1Kqcn2LAak7yFJHBtbwZTCg/0K/atmTTzuZNYupZ4OTl78XYUR6jbl
3HcAlZzDOcWurDLkI37pMPsHcJiO2BzSj7bHkyZJ8iPw+6J4+C6zmgVWEnYEzA7D
yaXxwuvQLIKcVmjjykAnBKiXD6QVCXVivCGKnlBvhHhI3foLKVi0Itp1uo7T4ffs
C3WDMXcaIb4idroRYdjCaLQjNy8dcl96RPFffkeDaCgCfXK4A9fRpYSAvjL5T+TS
Fm4MDV4i8fDmdefShLHyyGl2cEv0BLLau2sAzqVrIA+N3QRLPjawWnGFdKPr2RKu
qblnkUdqbMvrIkN5LzzFDWp+F9m3eO7LnDFIVUuLyb1oOamMn592q27A6DqA7M9Y
liPO5Wd4GiiAZ4Wsq3+fMUMH2nHPz5U8C2tyLDHJxef1VSfH3kLBpaeZnxG+MyRV
auPa4Xo9YiPk7gs68QJpjuY+4eykv8EXz1iObvud659bS5o/idEMwHZ3lcVfc8qd
rUTue7vQ5i/VAFqTY6cfqq6DJc7pE+s0rQFRd6wCsfQpjAyLd8pUQXVj6aff6MI6
zQtLI/MwpfPmhqVNdtt494UXARf1KraHdiQs0521CaXnVkBB/s56GYII/+E3fjOT
YUbbs1NqMCpZBDkrtAakePYZstvdTn1wRR8Luo8doggEUIsXlofnZXfEGlqfJQtG
dUMJdaG2mt5NBlIS4S+9uDO50We5/hw6W15p+Qop9+/ad9XuaaZwt/6zqZ+O2abc
pGCuYMirA2kwya9+8HckkBH5wFdbprxe37JsmybD+t2JufBi0X47ofJ0NkrdINEJ
wPWzOMWMcykcSDVjW3kfEkKTZebmBNxpuYjTHLplU8xSKH70Ozolkd7hYIMViNd+
D+QdE7RgEI5FuHe3YgajvS7jxkrKNvK2i/Jnv00UUlXp+bEr3SmgBp5v52YD3WYi
V3U6ebkrBtyJ714BOXIV2J/UrclkVXoiZGRO7f8ob+6JWgOveW+IIoW8kSBYKeSV
tgnaedJIhVmnqeS1xXrzgeTdgbRnG3LiM4MumOiEPq+9e701ge70uLxzwQvbY7/S
2a5m/vwPywkT/GdZHFcVnCbqC9hh7exjREP92/doGtO7CD6BhroZ0TsV7ndx8VtN
vYJO6WtKlMwnwmXYSqMjKrARZAtNU6Zf3X9tsZ5XimnQvEU4+mrEcJjvWGXBQKXU
8OvnLXfY3s7sVPRhHICn880VIY26Y3xfnmB4cF0mTSDtnof9Vr2Jv1WdU/lJeHcl
Gd1c5+IJ6VULI/IMhgkXPt9jGSKaUODJDcW1CtaS74hj6DVjnVdFwI8VyPxn6QK/
VtGLINZNp/phdTcJPRGdyu1IcbYm1X5bGLnKte8XvDoO2pX4zWLWiEUbXCsK0NoK
RdrlbOm6Kehfp5k8ltuJte56cc9pl/IHMB++oC3IwPWUnV5bxHH+bzK3HRUzlyVh
QMvfK87AHFpn+PsRhcpZVlMNGd82ZMDkFFBHBuSV3NSF6bopdM40uqYIW7sAVQy+
J3hVfYVSpqKjXtqJujdChYCqk9LF8q4YvSJ0TD6H8npVOrZoLnRkZ3qwA+6QoKa1
whmImACkDjNs4BJF4dgDOM10rHo51pGBV7MH7gUgJ2Bmd12qHk9qTxVr92rxqRbg
PzzsduNdyOAuTJwmyWuvz+Ko3hQ3sG05Vx0CKGFIgdnnPwQz6qGD2QTq+EcFp2Xo
BEQAG26YTI0LMSQAQw97+XpCpml8EmzDWLUi26Z8vsbhAaXDyvwv0cOsPqqTjTXJ
f+LOL83Q6guWID3W3GAdxlmV2ASkpY9GANFSk5ZvA7uBCTmmHgYn3rbRKE4RXlQ3
flhKeSPsjOvfMOrIVbu4c9U9YPQ7LXbnsxr74m2S9aJ0b9v75NMhYrUOMsNzznBu
h2o0CK9C5FIMVVU705+3woCbHWm3ZIxgIzJduG0LLlC3xh2Se9IL/LocQiEB+hvF
hpu5nB/8WsGknWQoxPrGEYPfxsW9o7EjQ7gkAvjIfVUKj5BeOqvYOAcVrbJimeTf
SM2s7Z/zCynMAGSt2D0iwOjspAsELUGvcLkmClnLMdH/Z5dDwd8wcdaN1mThB8np
T8RxX9uIxOUJAxjcvwQ1jFWl9oo2rjdYF2HnwY/hP9cWIv7D/dg8N1yodQeSfyar
4HFvJ+4LnUDuJcCUoPMVSpb9JItnEYDIUmL8q6TzkjrGqMoeF0mQtSTyTw6r6Bnc
N3cTNt3HmJfDTflnWplbp1h+q1c69N5EAgV0wdBV+hdda76X+ngnZ+vCTU5Cq1kD
HTJRJMrIzITq2+NhfKRze4/C/FcTUiy7zZ6NP5guAEu3JpMs6o+EgS8qvTUacrff
Yu3E/rdmIEsgeKATskmIKCGRtnWy7H4d0ynzStQRqxIAguhxNBkDvpNrsagH9Jvj
K43DkcvXpanVfupOUggkwgSDCyNImYLCNpQuUXqE5vl8rD5emnHmYJBXVQipiKKz
k4axlxOAdTtX//vR5BbdmhK+qKQifiKJuGqaOEDjrItE/LBgTRfet6Cqe757UOfo
TK7oaJtTqFnMPQpyx+y8akhYXVKK5hEWo5n1wr6P3PyVrGo+i8+Wg+sxFpzm0h77
rj5+JWiEbx+4/UauIr2etUwyGQ6oc4ukixFi4UmgUvV37bwFulbV06XBKteTYMMk
lQIXaU9oEkqS4/DK4QaHTT8spBu0YfYLkdLLdLv4Yk13q7DeUUH+eYCjK9Ps2vln
/7Kp7XJjWDk/moyzLQzmltvelSYtQXba1L4D3C8MTlF8FYkYW52UNRAdB/6/33h1
zkvhLPft4Ifd11NZVsrlvpW8DEKAATLR9hmTRwVUpSvW3nL9oqN8/fcXDsyfWI3X
9d9xrH6bT0zjdUidlcvSMiZ2oRxsCpQ80Tzya7zofD5foeYn88otBvOfPTnIhM9o
sTSLULzTsDwnn7LqM/s4ylh5XDIegBAP+G6jBp3bQCGEFk/55CLNweaPsJZqDoVG
j6IOOWPIWoEKHTuu0R6IWq2cbGpQyPtbz2rGp5hH90S9Mrm1+I+Gn6QbZZLOWLUY
T6KTdljP86QdEMrjAjUbP/Q/NAqpisf9/Z2krXcLZiSLggm+eEWX7ZkR88ZY6vTE
1gWHGe0y8ZxNqBJXLjDJ9J+oTUvJ1zq3aGQzKx2ZvjgRBhi71jmOu/tCBaT4YIjm
SHKSac9zqm6PoeBBmYWgXn/zDyVx1XMR9mhYiLLWUMwrif8JW2sfTk1V8/GyZitx
Vi+eDo0dnh2Wi8c8aautMPfAuGC0NNYSJ4k0F6xJG0EWJHRioqfglJPsf+Glf46y
uRNbcAVB24MNLfOgdxjT5OIQO826g2zYpFD3Qf9LVNNL/Q+HCcUOyFXnQp+8UWST
/gpGlUv1Kjrmix2D9LDuxgyMLBuEMTkvL4hGEEGoRp3XIEwXEa9Fjgggyml+swXw
xJr5f/JItUeFdPgbn4WCZ9zibT2iq0NOdUh/8tvitOXkr0pTzjsE1xWSvVE2zdV+
z/QiQc7a5OcTfFmq/UR9pQdqR2yYq1H9956IhcMXcBrhIn79JcvkeQf2d3noICcZ
RVsZDaAhadmzl8b32yKCgS10Wkdadeg0ACPuitjRUDZppOuQtup8GSfhgL5HWp8M
P1EEYUL0wejXrhHoSkAtZIBL++1GEIQKfVrbZhTcdWlAfcFGVjxr8LYaWKf0DW/k
npY4MgARZYCtj0c+dXDyaabcbpYvU+Q/MKcTgclBd2hCPvDDDKi0Me6YXyFlApmI
mvb7j9x7eUTicZ+YvtcfTSM+Ipp1P1dp6+N4a1clDG7DuqfxWwfiP1l5222n0CHp
wFIOd4uu9qhpL/nWUY9HY+5P+uprgYwZe2kFCMR8374WBRzdmCmDMvQEQOU5DjAi
HibExPF+Wq2z8oWMhTx0I+a1RA4n6D3PXjgPefgn/W0oBQOXDlLNxCmtjKPpUkcn
dW6ODwtclQRyymu2HX2w9DwtOkjVUzgafEltXGuTs01dGZ8laxSKnvsN7gkqV/9t
r7WMzS8sr0f3u31bQk2T77TJnxB5zMAtt3/RhwbvcmHYA18P9hWlEMvUGaCTJN5A
GBM9unQ4lZC0khvDPKIgUzZ99O6Ej/nPo8pqgjS/efkdnJijqCJU0jt0VDigL1L3
+exLXKWKoaFd6gc9Ln46gkTv1XT68JkKcCrY3b6WIJhJthYQyzOfp0k3SmQbv4pA
sJpfcSQeklZt4QYBU3EhaiU3LHdPuSDDc9d6J3cSYVOOnpLtrhhM00tApaq28ihv
KgIlqGOogd9LqciBkEtUTnLe9zvSZLIViDzZyfKQ3kNPB99VETfNf7yKDf0EsLwW
q9ujhtOXtcdcnI2eknif9ymbdRcHBeIU0oBQOpOe+iw113CmlMWn4Ju3QS1nZhsH
r9Wtlx2XyfeIwjQ0pw0uZxm53puYEZROr5d+JNi1BrGYWOEj5JDcRMhrp7/DP6FL
/BYmrWXuwJ15TY+i7WUDhczF273x0kd+6XrYaWTYx5dfUdzSMpsEsxIdnZ6nWF9j
5fPOzAlW15hts0k/RHQlfZdSS1iV6Yxtm31K1UAUYll/4nku7zMTPEFtML73xB3T
9JduzcC9J/8COCicT2WiETWvnbMWulgP6QQiXJFxLFCfr37md2MIY1AFrS9nsfNw
GQIvfPBqetnmUMMOMkE49G0WEZ8ttLiv3w13oX2o5AUTyf6cgaDllemVAwy3KIWX
v/jWj1ZFmFzBo1jwRP+r8ags/xEQCWBMJniObdK5hr2aiLpxTNaekAJD6xUtQadR
l2qC0ugAjKqJY0Qqb5bccSvaYCQIbet6iCU31kE2e+TYZYr/JnLpF6wj8vbvpst6
DBeSOE/Lj6uz7B4VBLyqnRE4kAia0cH95LVawPm1mjyPJOnWRP2ZCck+Lnk6atrG
BdHhhoMqEXjVKdnAvbLdq8RA/Su5lVeSjZUNTdvwLpf9SF5C8S+HRNujZzBljNox
IKMU83ihA3s5RDX+lBzgeQ65SjYs5mSOashYze7inZOTGKRFirD8mD3ILtR9PYv5
a3O1E8Je9jP0iJWK2Y6sz1M7uR6aFN1odt/9V7mfl2mKZRJ5YIRj2jBK+O6JOIGd
xf7ZPwisWzI+8xrHa3g16415be+b8trkuF+9ywHau3mNBs6spGLGI42ceMNBvJOp
wxzzcCmxWa8dtWsn1g/I0E9Q4zkV2XmPIdmUgy3xEPI5R8Y3W40Ky+7OR1Evv1uQ
syqTbeAahCL2tzKXSs/jpA8+XzE3qDFqC8dN1vOHk65Wg3ZBQRrzS7cMAu/t2KXO
9vcqP+0kPu2JGfDxZGql6+eerkYHMJEghXfknUWMYA5cx7FL42F16LFdSsl/JRPi
mH+ToclM6hzIbbdH6JMhNMaPUstpUNldWAionDAT7kv9dFGAaMASxUaeEVVG3e1m
UFVeLm4oPG/lwpCefOvxEs2UA3bODVeUbqa/vUYuK68Cv83tIbjkt0h2tozuvzPL
Kx5NKtCCAdeDIWEkFKVY41WVYufYZZnoF2EwCr2ZqQsU60FbsxgmSGCw++ztQ8O9
7lshg7NDHJsaahxYmbP3IrFkvEpV0L/q4kFwikEQLjG7zdQ3MyPkXk1detxL8omu
S/nipTtCxUoUBotJf6QFMKE6bimN1S7lrECBN/jYARmzUEpQseixPBpsc40H38Zt
vS+HqAYkAgq/82Y36puaaUPRfjUIfquwRBKJLqktEMpLvBBs/HQHkCshvnJLfu59
L/Q7HPzGc/E+EFMTxFnnYxTH6UJynAlv+K/dKBVygEpbK0NPE2hTCPHJjnEVBym8
QStl+a7Fl3wYb9G7PLlzoJ1aVZ3gQqsIGrHb3UnN0ftNZP+cjy7k6AHDO7vCFmi7
Gm65bEBJKCusn1mFiaNJy7W1lO+UNx+XGfLCJypC2nZmRzYZoVXxQnsOg+pjzlAS
cSQXa5GGZCuyFADD1ilj8l+wknHWc6696u6VZ9vNYPkMciQHfZ10FroxhEuIUsqv
Vz3KkdAkri2wsYwudSsi3zCxhooP8QZewf7P686exi4YUtjhDyiI0ydU+/Mo+UGs
q5LcoscVp9gttKLZyjLqDUa04UKlSDYz50LG6hXJowGVll/rE+ioecsLt0mgY18G
QW7mgfa0A8oHGHzzf6JF4Wz8f42L+OYWQcReMWVglt7Iv+cnhe7agH8qAlQHypoK
K/5LXuB5Kn3QJe5OclL5k5U2EePyPyigcs/iD6Yv0XGU3abZs52OlET5Fhz5rRts
IsFj/ydapmXRbyx9DHjArugChQxLMVerowu2yAqprd71VY2jaiCIts3dq1Ve2iPy
9qeIv9aM9WN02Yd80Cu1PAqoysjRj5mNFiLvhn9wh5MKYvIOECWzOz8bAETMJLjX
8ymr5Eeeo3fXPUCSPHlMqwYHdFzGNVEqY8/d++rj6M/gjlLcMvIVyHCEm2UYjCNT
pTmpzgF4I2U+/XtMtl2+U/jsYXWhpRDNC8K4Xcge4YzShQdSxUWkD6FOLGBhEjb3
795x5mkNfhJQmu8zul6YRevZ1Pmx8a0eotUJvU3V4SfJa8tyShUzvlQ9XxKHs1Qc
mTWNnRBHVRqjw0SXtc8Az91In3WISQwolDoek1Yo6V2+iI7vFtSa1tBUSml4unEq
QfB4DtcNk7knsjx68G+bprvakeFtJroZ/O5YXomfK6/4QGAZbPb2QkwQMuCN0mJd
3StrJ9j7dNGeagtTs24vjhZLMyKSiCmNZlQa05rUm2GfcUw+KIMs/0Jd4sBgP/OH
Y4gUomTZ/JqTDHjkNE5tNhhW13jMrMiLjekM1PUubOnqsl+GG0t0tN9KrmR6kajW
SLbHYZEkWxnm3AwcVf1ag31AfqmfwWPA9Uj6zX3ca5tEfw0KuFlJU9kOe6/1k6nO
2Tc0rl8KS9RLldNziuh/XZvHqLfH7yrs59/UIvjntnU1bIrYv5ouf7coEwwBulNS
wDNbN+Ipn1y4lPBwMCmNFlBkEHbRiWtunHzxZc4YD5ZFj1y6jHCgeBDtqDJgBf7A
9TLfJU4TNwwmYJ+aYVWk3n9bsFFx2/4EYZZPNiydbPfc0Cjyn1nkpRn4XXQpm5Oq
6fyCT6Sm8fJHYs3hmf0OpukvJnql22f/uMQJZKsFfh6s/78L+kZQoKBABjlIGZJc
mP/WgIeiYsE2yYoPogfoC3ddBYkY3l5vSWuOmYF2VfSrhHWVxRS0es23ywpkplox
xSCKKBpnvaqLgOFYJqrADYP61kuev+BZkutkXEVdKRVK7fQ/qSf1Ius1bldDLoN2
tsIU+TCeCGAvgllriPNe5PmW4XAqQ1n/b3sfQvwmXuiT0FaHI7n8ANsRW7OV/7PS
VJKMT+lC0fwvCUly65GRudBjMq98BwjuiR6LNil6MersMRF8FEt/sayfEbliatWC
Zu4DVv0JWV0N/6eWdC/CWboFxonHkVD9uPrYtVphLsqvqxW8DUBQyJG41JfjMAr1
vaksJNlFs20erg9Iz3ybsz1JwNtyjtJhXkeJH+DACH5KZGM3Vu5S/kDfpp/60n5M
SwPrGIHjb0QO3K79ZRKPPj1CvC4n4/lLSzIPz/q5oROJExI66eesXWaMv88pVoks
qyVwvTl8ricOAx+Z6yCEKfAybHNxBUTbS3Kqyj8HarR0heG6ar7FWDeXpmED5DHT
GCE8ESmKhlZtUlPNDxD91pFOqz+UmF99+9qIycaP6v8ZdGj6mdx1Wup/l+MAxIez
XaqQmciHuCI6OHU8xEnTTjnF6+vlAW/6CrwVpLcyrJv4nT7NQUDR3yozjz4ujOrf
wKLeGOG4Cy4vP0KY4vJ6zMrtp51j5Igho/JCA3Dptg0/pLGBu54OHTx18CYfui9N
eb4fjmXAIKTjUbk0IWU6vzsLOIJEIaBso5ZtY6nHjfRRQZnRhUWmlCmNTSXCA3Cb
xTAgMlMq8O3CTdw4SQyaXvZB1myDg/YRRYAJV+/JZ6tdHlxm9YzW/5Ka/2Qv0avN
wMvfhzoQ0deakljJ5tMAF891Jr7x6WbYrfhoOA9ZrWIwyy8BJa4TXFVjA3U0LSZH
ywt0OGp+heLemUKMj8sA1Ah/QZcw/kuEbPjkr6CWozQTCj2KihbzB25pmk3s598W
lQzc6X36ACeGB+zptwS9fH5Ld1ByPMrt3UnU4LZWe/524w6WoIF7LwBuCcO2ek62
hBlhkdxKiOMpoDAbv5OGtkDVFWeXmoigQFek4CYEy90H1CvHeclkK6w1qZ3A9Xpd
HRMFZQUZcUKd+1TjnXnqRN8jLlUtpH98H/BxFtlSKCXdZae5oepvKftxE6LJwsip
JIcM2vqckA3re6pyJkaiKffE6xEacK6z0tzykmQU3pmZYYMCMFpPLeNKyPbpxkZZ
037AR2oSOKLz3JXnmQ4WWdN+YzdSC+y9bDF70P0/qwBJ094l1DsYt0IIj0WsKRzK
oLA7BfRroWP+5lCVFegsPy1McxWhmdeQ+RJd82a4I/WRa8cM/A+oWCbXHjof3pkS
zW19oDtTw0zW2Hh5J6px3r7mrQyzjhXLPVseUmsAQZQuF3M6QI6kMtM4JoU6ldJb
cIbmGuB0EgkiVG6h9yuOLwROtK2jaTKMNJBhMH1iTWs6EX4qd3ODkKDAkmrelVNx
sOcLkbgHE06WcWofuz/6/MsWkdp3mTfcmXJBGJ87XB1I5GQe8yeuZ1kKuumTigYL
0oy5zDV8R3r1dJV03ZxPboGx729MuckjR6g8OF0iLQtcF8VXpEUn7pZGdsI0fTZ5
EBkVLSHprr1Eakjq1FDV5qMPiBbdDl18K0JZqpJzGKubzMdzTw9TzwzVEx/ZF32p
eUqakffUU6pGzFJFSiW7esJVxtSfP3n6I6XDux6PX3Bfkvab7ZYi3JYKh2z81iGx
DmQyBquz9VbVQG5vqbws6il1ZsV8m1YPwH4lmCHzdkrph39Rb5mV3o3baEm2kk9J
DHs9KsY1dthSL5phVxSWTKl4HcND/HA7OikazKMnwdXswAMBeM2UdJzCWiQXxrUH
QAv5OHCkbT6vVjQV95UMzOoNxcDi/RMvj/uD1T51Zl3SazJytD8xT4x/H4ByHoaQ
p1qDaUXj5Lg1yl19vX8sBza4iF7OnmHdQ1klT6T1+y3VdJlEVm/UxD/JoZLgYb5B
qvWrUJhN1gtuLEyhef3i0i94BxVW+NYIicCm+nVdA1jWAM9IP7LYPjXff/g6P9Cz
YRftnqT/w35wgxZiFHzEbI/LakCZoFfnEa7fGqzGFnnscA6DGhJPakb23GAWNPBp
vAlUQ2Ce7YlzMCPMBA0wEADODCnayk5Zc2QH9OrKsoJCVfSO1bgIvwtKQJCb4fjc
ZStFXWS4YAw68GsTZCOEx4m1sXunzZubKQeL5NWI3ku9MjAC+n1Vse5hlzQ8HIUn
SdDURnomLX5zy0ARg6j6NkR2eIX8ygk4GCHe6EaTAoUStmszlLxS3rYnLMWbfbNv
TyBf7r3Ncpp7/1cpDcMhlZ9+hNkMfUhGb9Dbb1QrCKXupDegOo6KBwipuwnHPU0V
X6GKj+TGOsRV8RqoaYzd+r9EIyT7Voee//2jpC4r90tGiSYK8CKKW0PsB9q+yZS8
c7tVi+D+gPLYrTdD8wWe2Ui5HL8byTafIP/d/wZPYC1g0KJYIOy2AGNXWf7/FESi
FqSe8cs3XN4yJN6t3jkobMms/UY/kqN0+m4wqNtMcT8EoWqWKZ5bJEaampZxjdSP
olD5rVFV379YIaouhCURCwkXUm9q4ZvAfrXsxEbohCS3Xgy0TzV6sTywS81qikkb
ON2cUN0xZt7CmPpatWAvH/9kGK72k/i4A5DLN07f9UhV1yVLCrk59XW4kspkR65x
kgrJU5PpejlU8BG3NTt/S5zVT5kU/ZMOVxy2IBv46fwzmDMEjPt3fcDVzSkxPdMV
T/B+/UjjPJGS5rJR01mT+reO2Pe9Cui+rU6x5wp36rgMnmQXLKRtgh4cHV0apNuM
sJ64ii0V4RPYjiWAhmFmn1g4RkXn/r4JXMGBZArpYXrSJ7Dy7gWqFCSmXW4RVck3
9QyRcAK93YQL7HV0xy2hb7WOuOKN7uAxIOC1H21HPcrU6x02Ye2oLyRZwStU9CL6
4A1Xo/qs1lIBKmyoEH5EwE/7NV3Zn16RnbiVI6iKq8iCVz2NXlKheabEx+Dib1ba
shTrG1+kML3+foiU3PmYT8gePJu9GaYq5vNKMjvNHGTK1k2qKdAYFmeK3993Mq6k
tShXGTWp50ZO9rYMHul8aGnaT2ILY34jd9CpdUgZki/4DHd24zPSeY051wXzqR6n
jhJebfyKQSddP9otH4I3D6hhTBPxSUAKyJfw24pIsoI13dXf3w+ipbWd26wt2ZRr
jtIsHzHvZ19ikRHbLaSKRIcgE+AJT9NFMpaB99019rpp9/YHPhXsdM0yQwc7b8Po
FbnCVOdmTYkqvDXs4QvzfBLcLqGfEGIeuubdI7AWrikxDKOEcgLWGzwfAvkb1pK3
YF2qBd8Pivniexr7YrVKOiawV9ctqydik7tDr105rUVkm+HvNaX9EL/a0bASt+Hx
WEJQEy9xWso3EfQrcIlfbCp94dzzi3opmdr/Wz0hRMn2fBkwT5zGhImLpvspKe7D
L30KNL9SK3HwqMGqlXFiHGtpXot5CGlLMRCCmMLmi4O7pzBhf3wt8SNeB4DQm2ux
nwi9BtCQorZ3MRemDRtV1CA0Oft752QYaod/p01m94LS5TOvTBf1CXS4vkRoLijp
yUZknx7/nCEyeqH7IucCPOcQUpAbmtVDD3BwUj6WB14KLThH/tP5Txe6mGxG00vw
jLmDWCXFe+DVq8AkarS9NKZcw2xhi5Q3I8EIQ7Y2aVsSVm7SVGalTznmHRvbJNen
Auzs3wFALLrzH5H3ahd3Gr/P+YV30UT36LzNFkxDAFawuJ12rdF/jjLlitFooljQ
tO7NwvYj3ZsTC3a0aRucRksTOVEI1c5vsniDTcUzs0TUVyYPo+ORY15AVxE74pER
Kz8INOf5AWgaYAZ5AN05lCkSdpBfZ3ono9oGoztuFuL96odQEhQdmA8FXKzA82cB
jysyUYEV/CcmqN4PLOaBw46i2i8qYJdKI/lEJRLvDbcl45lt+n61SCas0+eDfoXh
R731xXyS4ivJ8D+JwI7L0Q9hhGfquk8/xL/SU2NoWcTS/g+7DdlLyAbXwMKO8IKF
rgj7Y0DMGz308oU+cNvlW/gQWidVLv6mQx7ncF5Gn5a+WgmvNZZy/uermw0D4Bx8
dnn/XGRCrZcPVIK7HJHSRDCnkOzG/LpPVGLJ1AENPZoZ694g5KFz2eG2CZt1HVGf
VWUrIcEn+503DbvEPQTMHVLw5UpyZJ6Q2z3UtERo+xS2Qk3qiHE2utipZ2C2CAI7
bT8PsFQRNMCiZ+7UcC1ppFRK9GPYe4BZWWvLJgBGWRCKvzXLXvPGXNzykqe5E0Tl
A4BtRc4CFVYgUWjRI1h3Uia0EH8f4Xq0+Hn8mmfbwYKUnyBeZYtpxZyfDwQ7P0XA
aR58z2c17zHXD5KkNvY6/Ek+ocDz9juTaNhx+nycK1bPFfAiLu0JVbHfSwTLyhwq
/Qsxe92qVIzKX0Pv/kfS5eciPf4hbp3Z0xNdJPBCkfXKNZBE7cVWqGuDn/5zFPOA
BoN5JlOz9AE7c6S09K0+33e1/7XSP1e9ZvwqceWsrotwV/V/B6VYjReCA0LKA/H9
vl+xY+udb6nH1NlSLFcPLeAcJ8sJJQ2TVO/8+nVlYmpK16RV23CMES0MS1L3ljbm
hqBkhPQBWFDgWj2Dbo6OtaX5/BWodICfPLd2JbjkoNMvDjDYvqXhzy7ch194H3yN
TNTXR5RrBlN0AP0zl8lBFjhoKRO0M0jVghqQFMDziv1M6Iu4IjLFu4xMSY4fC4QK
Ikf2GjPaCYLeZbDZ9pwPaTt7jHWPBpJGhPxHYt0LXA/JACgkh+rXJGtgrHDZ6Aso
7Zi8WAZmsBtnIcAB6YJdrP31Ot1eNbXcejxXyPeFtLVcinzXeSPTLJ75fEklxpFz
JUv0JFNyIiWqejzSfN60jxLZ8Y7Bogsbj57NtlvjVwd/d7ScZGERnY2gzu98QHjt
LMV9an2N8xiR3+jll7MHzXQ8O1HPAQYGrqUOkomZwN8kNdrObTNr+YUIMh5m2wr0
AnzCqwsShg3M/H71lqyIWePP+n/r7l0oPEb27LqYAz09EgwWNpHxEvVt2cM4zdna
nHMLf/DNp/iKvxrcgVGub4UUUOQ1MDwPToYsYsNpZJhWqDG57y2fF/3TFFwf6itW
iNsYO4E9ZpPGTelZvh5+PIHRLiw3+sN06/b76VZZ/uAh0Jz723/HX80R3+y67Lm2
dqG5G7pIuQwTmZfQOqt3oJRkifIfyoiaYVvvrzwvavSTiZTt8xdWsZ/uJQbG8CVW
JljSEz9HqrS9dk/awFAtxqu4TQMgXaBMsPyWb8DqgQ+dS834B+WBMTB4uTXSfpSW
NR7Z0vGRGK5M3MvrsTIxRrtsjR2fLoLhbLcbZNiW8A7DIJwRhN1fXJuLuMvMSZIH
lIVF2OTCy8VW+o+q6ulvSEjilbK4EPIaoC5adTmisvbKlJqvTQxgDoOWSJ2vd0h1
+d4DRe/DQEUhN6sKT3rL0i5/rxhfZjUHxR964LD4uJQBIDe/d+OJ3hztFabux+l/
q9wZLSk4p9gWLI0kOWxjNgWcUi8gUV7aS6wxXiT0cefWq/hkTthy42P9BVOXpK6c
nS9zjzEznqRonvFyG0qGfp8IvlFjKNfUPcFmj+d4az3VwZNEKmCc0j6O/wSvapAm
m3fPzARudODmL+OhG+UxqyJC0I5YlQKpljF+UxBnrs/bdCiSCqqCJMpNlTjdqcZm
6XSW4qzpsVNSEtiPhu/ES3EhQm4p1UvcvebdD/c+eYHuOc8xErrKwSQ4CcpUqu9a
lJGXXQx2nlg7ibfPTurd1uIAJfPRyxbxfYyu6Q3QddYcPHradd0YHtGm5sC69DSs
q4GZZgk40kUn4sdm6zG0NG+L99EPA7TOE4lesGJ1IW1ejLw0AP08st1oWgFKWiok
wmgr0BPGt9/H71Oz2yPVQFEX8w3bNbukxnaUwrBpAp3j30BkufAuA3ZqxYf41+1w
4oosCYjPRyHva2nknan2Qyi9dTy3Nr9UO1OsJlwIf8ByJyMNnugVj5LAd/QIAL0k
MiFxpNXy1m8zI/gk4YNdLBNRclZGs1JsG2rlblrB/le/ay2MUyNdQSc72OiElnIv
0bxzHLmWkQn47v0hCIC/USaxK5UBpKDLvQVQ/eaHUMi1kN1Ln2QklvpEjusBFKq5
YMr6tccvn8n9W/FDblUzDXxiApm0VnqlPXqE5RBVPMbHPsjuBxQZrInfV0pZQD6c
Bx/svflkv6UE6+cI8ojv291jBij6npd+U5prjnjQMRhwxExnGm9kwvaeHC+NJHI0
dXRVpezmwJ4bULvpNSa03ShhajIsG22rAcFQUlPB3xopl5ETEncVprWYaXbInyRl
/WWRHRE57W5WHrRWa/eHNB9EPquN1IzWiH778i4O+WeUrutgnDqGYjqyT2SR4O0N
EQAeEjNgYuUK0f2I4ryWG6ZPaCQkmKSjf0YKIvo6Wx9PqbDF259OrMoz45VxZ34C
HlDok0+TiH0/svnUWXvOcstTXLUIvmQZ2fxIqth2KvRfV9UFZ7hwU+GVR+PEk/JG
eFJXlsAojYA+WIJUJhNlQ1WXxOcpGZZ8ApkxXBL9PoOv8XmF6A9+gCwoo50dWY2V
HogxVDdK7X8lg1p+B63qEWjIkRJ8ROvrnfjMW2avTyPV+9falK5Xljx25yfJA6s6
p8yqpoDvh8KillbN95E6oDa8UIVSOqMCREAkvGMia9bVHgLKEZSRtqxBonTDiJqI
k/cLkI25wpp1F+mpXwlW722/PjiBtL2TybFEy3VkxW5xUqfaiyeUmUNmrhC1ZG7t
IIqWJ5r7myIY0BZSAURmUkbokG6YENI6swQiHo6Ub7jpuAhP450OyiCP+NcYcnZR
vkafGK9odHfneliI3K+RgrEnzY8dtS6dTX9ZLMfnfYWNOWD86gqhEZ30UF/wzfK4
4RTK+/D7l+gtMYTgKzQ9j9CNXLmSWoKrmWJr3wb6nwXaKO0WIewaYb3kkHWFAEcp
gFg1r8x8JcGa4WxDEGJ4bSNzgavo0QUn4iZc9B6azlrTDxHkyoIvFqqWKC35Nhea
CI6oEkMBlJyny14ChNajb3jI+l7Tl8XHC1FMk/Tyh40gtVQZ3U/wGbaC2lvEGWWc
fjpIl11Q6BbhifFxdMpBmPoFN3vqqll3b7uNRo1LXOagBEWwS3F43EcFoFRUwDop
pEM3ECoY4vsX+z5wjaiR4bDtRbGCcemTDtwaJeDFI3ioGOd0m8kLTW+R3MNYZcwp
jelc3YfV9xR+NxyiLgcJsx+mVtZ6eL58dUcBmsZSckyi72Osm81Uiec3BYv/ftxV
prBBRYCuGsadgrWMCX5PbvtOBYJ7bBy2CIAmftym/SZ5IcjaQFfWTF6gf50Y++Po
+RtLvZO2hN0nBoJUDtd0ZV/svfOxzFNDhxsK4QSvdE1Cx6hQKajUF8MU7M7RTf+O
Lr/U3f0S2ZNrTxJ3d+KKgQOy5T21G4wHboQgVToIlXlogOpoCCLcJqpUluVRJTJx
v96edXT/fJj8V56UTF+OBl4F7hqA2fBJ+U917vRejzqCsO2RKDej6S3Xb3j+gN8d
jxyCIy+xrEC0Gfiqpjbf58FkFNihYhXqb4psJLkxPlDk7/unGm6VSuHcqo6Fw3HY
NNn64nlJXzUWEtf6T5FgLxtbChpvuiuFmzrXGTJTYkFb35+arYlpJ50Kta5ih3RA
QURIxtYDQY9mDVV+hgcYMZyosfrRpsd2syuZzTAhkV2AekifmvuXVVPD++badosk
F6IVK3FCTcu/pLcrgatrx3F8MKPfbWMtcRYyodV1vfunNFnYuVzD+MjnEv+sQbD2
9fz3/Mrzfo8M5UYaD3xmZ1dEO0qElhEgpTQ5LxMPWydAHcnYXgCd45qgo/fXwhrl
kDlH9DJb8dDgKLoovP8oWZmnqXwxPD5jqv3kPE7eG2hSL+xAzxJE3qKFtabTGENN
VI/GFRsybrFDc1i0y+6yOXU0vGxzqnJrF5Ry7r1dF8+9CKOsg06Y6hI2qKgMoXJP
2mlMLTfsBVh7mjlqy2QmjAjoqXO6qTONmeNdZ2hV0/aDB6uplNERCGHZwlUMPvnI
BMMCRZRErnxzc7Vo2IxyL5JgwmKfObC3Mr0TQto3ZnlqJIPmtaziHaOM3YeLO9/z
MkGCj3+ccYHF8A4yL1hJb1Wh5pxPQn2AoYSjR85dl0ivrTEpirhPX0BBBAxSgDbt
YZ25Gpx4qriTmMgBx6kfaKr3ePMir4rHB1x8yMpQKIWeythzyAPPD08s7bj+OfrO
oTQuqrgtmqvi+/0ZI9Tj2dGNdjkjMrr/b9Mx6C9jxuI7pfjK/tGD3gSstGdUcA+X
4L09eTaBN9WH3Cl3SCjXparcMC0VqJSacBnual4EemFn8hhjCTYhSxfuQjw6a7LI
+ylpSlJ7+TpuKnzf788l/c7P89zNL6X0ImliGxpCIlXmQktsWw7zzNB0MyMVKgv+
rVZlZGZ+Dadgs9zPEERdaSF9QT3mMMf4r4cSFRxgHTFucBeuMt6qe+U11kJY3lso
tkXc2mNPO/+lf9sHuFn3lU68Jxk6Nqj/PTZdTExR8V0AAN4L+Mb9c8LABdNidAol
YT+0tYBdjSYymuD4yU2Ma5EAjST6G0398Kh1cjL6Q9ZWMfY2BvTz56CG0waC9QkY
vFEVHW9wqQEEQO91FyHMVcGHo+YcRqUQXSYHMg2t1AT75NKD17pFurVdrWC22148
x1k0djzz1XEXGmrLrnPQnatqBvNSysVC78jTrV2/bvIShz4eWsjkp6toHBkD6go4
s69LLNmoEnYiQoEa9xxUw7C1NkoG7JXqTbLwSSwRkP+Ha0vzXO8DXugcdVjWAiWo
p9eB82+IvLtlKl+jKg9smhs2aih6Q23/7gmO0qBw3TEpQLZxYkCtBP9Op2Y3c2EO
Nj+DwMuF+QLBpHJUQAKjONxHcQVKXCgWhmK0oXuAYt+xWLaY49s5BHbWHcfLJXqz
a5u468YGXXmrdfkKMIz4EeT5I2lTC+n3ySBXxKRB1SvlcKwsVvZCY/BYHHshxTeq
LkCCFS1as4hnfhK43PkxfPj3HEEpRRIgEiiabYxRd+zsTBxFFCPIo7cRLCVR2UiN
W0vpIZR7ubLqij9l5T45M/g/RIpXe1j8lwqiE9xYfWmZ2P+z/Qv2+ZpDeVtt5iNP
iIOoJBTF/lZ+rFVIOVsN0szSlFsT0YzSeCiRJKV+SJWTN1mbMEhdcRQ2hX2M7eSA
EaSPjXy3DO53aMpuegGvdzReYP6AQcxTmQsr53NeS6UYCrzkmE5y8BJLQQZCasg3
61PrXelRSDKJ6+GDvPrWSzos5MHO0BPYNAuj7nQRap3ZggkenhNfxOBMcWB09lES
c7+jRkVOUQwG7v+tier1V0ThEkcrtFmXBSeUFKtaAG3huGBJ3soD6DCFkUp00Rwr
2wzcuw51DUN+idMi1lne+81Y1d4cEAS0Ulft1AJL8jB5lOvt3sTaX5H0ooKIyqNs
SNQNdyfmqDEBygJQyir5tu5gNoteLIfL3qPityaUDHasaXKJ2aKboQyae6EOlxsZ
8DMw7cDGUJOs/6l+rh0FpjJbVIVhnWS+ODF7mOyipoDTtQwSDbrg/6yZk5NMzmm8
lkZo3rHjZOdOYN/0FkhqBX5uiOM63MAco2V5D50qcmXwYku8lETjGkKqN0EnnTe2
++69bj73NV8T5fldpOebcMBQ9z1FlzQz9dwRdueSLb4qVZHhSHuV/I+xsB/fRZm9
KU1uj7HJZbooAyPWtgjhv+G546kzFfam3sC2fOj/FYXKPww/YgPhGv0eBgZMNsTh
G70EolNj4YSQTOAnujwdkV+BOXOhnvdM2F4TyZrF8PJageTXl06QYjaLe1LaVzed
M2WJsfiasF2HG+BARTHRvs3RXssB1kLVi0SJ5b/dvy1j3/Jh4efudtz79BGIfT2g
l8a3Av+SbSc8ANu6bHbYGFZlya8hmPS3JprCaboAG1WsiHy3plMFqBXyKCODP8C3
IhbiBP6Sw2FDSCIGpkszI4zakMJcYryKDEl/h/xx+pKIzuU+AxUKBvAQn5+74Stz
XJNW40EANFGz2Qc9jvRLM43woh44RAC7Xtjy++XTU0qgDKhVmhIEbdcy6s5adfvX
znpH8ro0LLgxAvuloS8xBNTYp0D3FQ8qpVFi/h3TILM4l9+8tOi9HD5jYupNqCFg
IQ7/ij7MhYNi7NBhgpwJ7IsPOwzpsJjqlIcgpLlYapFhy+Ske16i308lA5MHWJLr
kJZMUd8BpW/0uAdCiuyg8nGWvWoSEPv4UqVI1sPCPjGiwKw/Dk9dAYoavcsdt09K
tAYmMXMEpt6GgikbwMAgEIHOgvLvGdBicGHBCKIB2Y4N+8ctPyTMG8qUm4ve3cKM
VSn8USzEIoHqHhC19ZDSJWvvFnIbHVlQfKpH11/rKi/NeVRYbq5ZabhFlGnJVdKD
QBzmwlrzY5b9oKV6Lwtj9CJ3PFDeRwqU7gBe06WoIHHbteV74GrKFp5YYHH1Rqd2
qMaN5F0S6clEp0Z20WgCiqrdSWqjl251UriC183nt+dXEahlmgsdCnqo8LMqlqER
qPnzMh650u5FAUVJv23YrvebixfXFKqmwqsgVYEApd4QA2PkUXt3X3Al30Ve90QP
cC+kDy32UTxVVd+5UeB6ISHk/pfuNPvA4BCIhX8M3FBr0OxqyLb1ZdGfSezE+K0M
b9DB6RmMpW2SJaqkvNRQyvHkPf8fSaT+RqwVxpsB8T44MD2ounjyFtDiTEx0shLj
vFC9QO9GrRcQM5qra20Zqz6o7BXMZWXW4N4GsZGPbjeO5qRn9jE8alhP2R6k7OK+
7ZeFU97mnPZrTK+nUnqAOl7T+W3Id47JL+oZiwrS4vHS/oRErrHHyxxV1pJM0dtv
PxX092QCPf4Ua7Xr/RszrEWWxiWIuHVhqn3fwSHK/GQ/UpAXlZEba3iik1oC4/OT
nyAqh8uYQGenB1t6TPjXoAgwNF4fuSpZARAZ/kZOqyiwj2Q43PGLQ6JnEqKdxp0k
tAVmzmph/u95RsbFIpXm2DSgWx2//3kczeNB7M2gjZhgeWl+KMIi6MyvDheA6I3r
Et6bS6wW6E9GTFr9858J/NIKrtEeZjWVMB3PQ/0W/ZrfTzomE95sfIunY6Q2FlDx
Ej2IozAaKfL5+5AFmimNtLVZEhz8YERr7INI/BGcgxL4hZduMtPjq3Q0TuWJbSkG
EzjgqPhHL8r/zOaqE5CimoGaM2PfOwiiC7oL56Ro4CXb8CYgVX7I0QU944GvOuf4
WXIzbrZTvIosZadkRV185/dU6hSUYDWTvWVS/ACKnCje3RtN5xHmhpKekFOM40Ym
zst/z0z+u67iy3ocC4uqahKDAi/6lbRAtQlPYESJvmyZA+rBQlU38/824J82jq0H
zCqNMpDQb3Ib7O2+mB0+9Il0RlDm8z2Ba+RBZkuhYldUzVawQI4LgETZcMukbe+b
MwpWfM55vMFP8lwwfK6IIu/iBK6BAkpvsnnL63XiOUFEJVZnLAcVfkQFtzDKY0zp
uyESjUAJMhaQgFQqe1DtiUAZkYkapnZ6oVlZEpeMdwwpkkz1DcwwNbZy0sjVMyoy
WpfPe9eFjiiySiR+rBipe1KV0x9XO2kD/2WNdspa3A8y/ruEp7mnjWXot5QF3MzN
1fdZskB9c+8NCjJWLflsZrJ8mFV+tBY18KsKOWrwOOMpCLAzHMnPAJj/ZP7pMShu
3l0BLe/r8d9oeJNXVQyCMpfzwrMAzvAIa2gxhjAlaVkxhWbAPST6Bn62muXQGozE
d8XckPlQdpuduqIy4+DD7McCf540AvUFVIyeDHRcpDc3CMZHLovv0qVkwaZ2U7Oa
jf6dsSnhYq4rlnM67OhAuFyz8BPdYjObi4PHNxDPpZQQVk/rRBi4AjHQ0N0JhtNY
wgLnTHozX/5JM7YTwol26TRVoukX4ghmiBeNlPz67JgW708eYIknS7WBfQJpDc5w
uLPE7Y8zBtWJNH4q/hPc38/M0Xs+JJ1l8f/9BIevrk7eLndAf3YUByhyOa6FAxUG
ZEhyodT9Wx6kicMXM+nyiYK6NeHF7FnYR/lwToCw6Rk8EgD8/3VlblSWm1E5sg/K
EpX9x9op6fwbPvn04WZp1i5R76ARcg+efI5bo1IRwVYWf/WPWHD6+kQZgFJ3/JJ/
8OoS43ODAFDvpvxb61CdH07wUmt9MkgHWF/zWFcB0+zKOzAKvJFdnbEQwWD9QDiT
BL4xCD8Ds3HwjTowdbZsCvThZBWpnG9GEYWqWNMNjbiECbXbVis/pwXOOITjjmUP
KddR3YKX3AuiFu8sN86/EHOW3Pmg9GDq4UCBddSzRyAYds81DfnRfBSsQYt7hP6T
1P0qc0Z3abKnQkfZ3flV0FdvMHd9NLHGO/jXYqaPZ0oQYPRospDsUzhqtsNEKYBs
gMQeCWpmiGkDoaWIJrtrJ6uHEjU/qRdwVh9h6rWUbaFhbFwfdZLLcM1XvwgJkbBI
plgT2uBuEeetwjwWhDqmVXLruTg6WLQ0llieqWd9ZIu4kZp1jmmaoYtrtu2nnd/K
Xgp8mRKQ/EPE/+zBp+UpPDuaRkcACXUUvm1PcUuWlsmDrB2Es0DL7Zl8FeoH5g74
Q8I9xMP8ZDttCD+DZBRYOzTzNzL6lAUvM8zm6dM6bpztVaQPLRuK/ATsNHVhP+Q5
xlLXpc7eewsdaxATSpxp1xvdtyfc6Uy1taWBllp2U87LDLb8U+i4EA+w2+QUWq2o
LRG+ZbAsK1KkIxac6jIafvcKVPT/lJx1fdCQKzyNdwoi3mZEPJ73RCzPwHheKSUm
B/bgK/iV3DBofbrwyxj0vtIGf5nGsSIGXIeXg9JiuSHg8n9VEsxtJ/Q5MsP/th8u
VbBMRsOE+asA4lwdqnqAJglXStXJpB9fMzlUQ31qV3q2uXGqkRXsza2JLk4SpQbb
ns3RJ/K/4Pd48foWJovBVFHAONAkwkcIyxn/orRnQWYtSpCcz7r6Lqnc/GzrQ4Qj
ja7QtpX1zskLtZwd+BsvlhxP7dl0i7PvY9Zuubgnut545Wj9JtCxObknmj/oeS0u
ZyBPNtI3EdTXjVj/HH2HFzRcltQBEHs4PT2d0pRm3o6z6zvMeeaZuy+QLIXK6i/w
Rn/P+GPf1b4BcbsRu9k/BcHfHPTCLKvDBNbGcP1PxwIjWFso7+i5x9topnimAi9G
eQA+MNldcwTPIgsBVltQrzshseSc18JKNrrxnVLUIbvHXYOljfYC3fxUxNNqyCvm
PE0zYcbdB1Bl9WX8aqUVQ0yPTEOuYjl3t91qgE0q0ECNCdFs3XsdeRPStEk//z1b
r2e508cX2RKOKSVK3ShbRqH+MV5B+3RwcNd6wTJH8UdK6K6ydd9/iDhIxZMi9J5Q
qZ8fVKSHr4WQP902YxAQWvXIyZFkBoASLInV7xmwomW3Cr5F0CXjAoaZ573MjVc+
e2bemFyDOzXHexVWyQ6h4OaV3FiBoutUzHwtUESwSqAB7EQ8yJQikTT4fYa+PBKO
G3O7J5PIngyPiDK5TigVbArnO0e6WhOH+KbOUEteJbrTSS1GnNp+oiF2rPIHYgK7
Ss3p6NvkDfGQbJJ5hRBkVzCbY2eIDUgVuQpY/ll1mDDeB4db9a0STxua0HxJPgXQ
TgwOCGrv+IBEFVC9hWlxBrtfU1CJZt6VEgBJ/GkMOIPX33CyJBpzvcFC6TcYFzZq
fjtlhzICtCsR82WZR728Tp1XUCVMWXCte+FupjJWfLklJLZxZHX1FnU97tWdKPwD
w7JrST0C9XT68hhJq9YkL5g7uhB49TEmr9eiV1sgPtaDbVlXu3mQg8G2snUmLNxo
gp4oIepQbUKHH0Xp8s/Ri3i0F7j9j19EoaJhi3yHWelNxaVrQHEMr6O09WQMNEJz
QZcuN49QXhLCX3YOsVtVrVa4rl3Zpr6bg2DuIdnWXHU9ZrR/HzlMXAoWXkoBQ165
ljhZOXDLgmSD24Tlw4LPS8U3wYpfB7z9ZDrA2FRM80g6OCz873WKxoosh9bZlpv5
kphHzIzVQtw5mRoOUvMHHZC1r10krPMb4Hg6hjVTxKt8namYq+IjteY+/HVE2OcA
AmmQPyoKe+QCjQunfCi9MLhfOV6/Wf7Rk6A048pXYIOkFzCEzD2taHK8t9olT19J
KWYwYrXiWKFkFQAQofUgTzRhOVOIHl+uLSUPUJmXUxGWLD3y5pVLEg7QgTlcx8q8
TPHEteX3x+5quRjv5ynC1O6ckvaHmG/QOvmwYDwzvELhHMYakSMyARiwB7oeoCly
1C45mhcAW8K13XD0fVITgrMDwUiBRmAfU5j4l71VebfSP1ynF54UKBTTX43QaGAn
k9Ur/G1vH0UB0z/GSbuhU/YfI8HcsZXj6V8M0/X8saxbs8h6AR/YC+35M4nHoyAs
aitI77HTY0lfypRXnQfscafIFET2Asdhirsks8HHsSK8zcbWL8eqPin+Iz9gWon3
nDV2UstVgT9SO3KoELb6YyauiIEl9gpca+NNoLpXGmEQYYlxe7HXxPvmY5S3v7CB
jK7n5F1ooi1HBsjbKrzdXd6Fx8W/j5QIZwBwCPgsNPExpfvDzzksT1lXwSIfen/K
d5Z63m6u8poGxnIrCcf4fMbqKOo1eIP25siHq9Uuv7Ml+cxQ0CcQLyCazHTnhGHo
/pBkBuoOq1xi1ruTv/0KrEhcf3YD+kb9wrL9R/VYxlO5AfRORmmhMqXOmSXAztGw
a8h6jqIhUE8x1W5PNeS4vbDsJhri1+jd1T9QSSkyXCY6rBGGzZjv5zn0wKD7CBwo
zEyaTxzqHjTxh3dzNpUumE0jUgA8/8rUUXKjKKpQk4jhjbzIUKzZmNRmRJ9TgC9B
6qi/PKpfSb3okUfdwm/RQkJ3LSyJP1BaC0FnbPoUIwfsGMVVXCnO8sCmd6+EGwwQ
0oFW5dJwjU2YoDWH3zm/iEyPagvi39FnmExuIygVTlZwhMwQ/LU/oCqTt37oJ1Ab
+ZpuDmLs9njfYYbODPqTNCNHogHnreTuJBR4R7qew/jN5OUaEBNOlqSJCDlS5IjO
hvXe9meVHd4WrT1eeK8AYQ==
`protect end_protected